

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
g7azmhtm6FcP7uNFjuXJjN8Z6yccOPk3SSjzvKB27peFKmnPmQmov5+YTGwYqqN9LpdyiUExk8K6
vPnJqontvQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MFrqn2K0Cr7TmQ5al162oDGiY83d+AkTWOgFyXPYrTNznygR/tx44RAp24ytphNK9p6shs2EFMg/
Qqz0l8DCWiVEoJ/T8vMpnAn7Y+poGVGS1qAR3qE2njrl81VcGBZJeFaWIudhfr/DLTuuf2T/dWDU
YpelM3KbfYNPPiPy8PU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FZca5XZouG+/BYoQ8qrJTmnJanku4IprIWRkO6VciHehE5WehR0wsZJhfKlqLEeY1oTPA4bXaxmY
NjYkrop4EOwW8t47/hj2kFLI1OKUAE/TAhCGg/aNSOViUbB3dUomG/y+TBuDt9L6g0Arj1vb/5Pt
IChc5ZdEfRr1lJMTpFfP+5qmEH6lePPdzgPZATPB4Zrj0P6EyiEsU1FKBuAKd9iYNGiLCxVomaz0
3/RwK2Nl+/l4mc7PJt5Hso+4s1qHb4s2wD+OgbIwdH26ZkEnKVFpaLiuWQKu9uhDLGnsBMPf7XDE
p29f+mrvP9Zi/3nonA2aBKrTwR7XuH+ZYoakxA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jP68OjlYJglq3zpmKrXOhq7Sex8XNW8fQKp4hUNmuw06OOoKhQASNTnjtyVjAIk/VXb64ViBu1ds
cNMJybDSWBhnChfJq4h9PNybShGJXxSm3NDOo5wUHKf10Eti3fSotB9rVks+tNdTEZo4O97kgfdD
G1FNOqlsYcQiShEGLLiEQ2yYtgJBxJ+jc8mFjIEfPhAYy1ElrvtFEpnhkNS2LfE7xdWOQdO/XoKK
ibeY08pgncTI3pvO6TMbXushf0AX2S7hgfk8ysZrT+0gktqFrJnyR6oljS6VVPLtRNW2vo/cC8XQ
Bzvwwt4cpSo5KLS4XxB6qClZipItck2AUEdIbQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o7jAZIoXlFbFtDYmtXhfRBlb07dhBb6Wp03mlT4T0FXtvccSHWhWZgc+VUNwt6TohLihOwvSipPP
XVXpGL4pUVYNdQBCVpFzhMkt6jhyUgsF5t10yI5Of6YEfQrDHigceoBukM3+/zJHPprrPQE6FUvC
wXSGhBCXnHJs1R+n4l0714w8/WftPQhlD9QGQp1qT2VARQXUKBRxcRjxe9TcLfs0P4xnN7uHu0R6
JTmV+MHmhGpetSZGx+B2Wa1MQofUPURqwE70IwBoUhdXH8+39DT5I6x2+wMY6RcVATnhNd2BCgPd
RzAhwfrcqRiU9aB+eNNdFR8ve9M2nGMmV2JxZg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Cl1Dz+fZIDYEIQuUd0pSg+5jknmtX/JERd+yOZ2SRaVra/4pU/eCTjEXMzhz4VFGYB6dgUxMsGBk
nL2WNdn/uaSPpi6mNF0UHQvZik4pUkYPrnRbFveVqW8i1t95SG0RW96uD19206lWrp5U1lqc4fH7
sfKHi8ZpU3MAg0DOO0E=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Qqp76m2aV9ue8Qai7QUavb+lhRYdu/txrnwYLzwTe0vS0S2OD1vxr8VeIT3bF/ZuXlTGm4S/UCSF
bgOPp7VqEOeGNfsSPK+VpQ+foQMENCQYccwKquBDSg/sLjpPK9uuoGLBLxjw2OwsRzplVFXiPcRN
LYK1/FmCP7RJBNgmhh/ti99a+WSl6i2YIIRGocNplQlG8FXq8ZTTHd/x2Gtdf/zGvJOy/fNsos6S
Oq9yJ0rMmbGeWbri5c04gZM08pUmXBsivgOHm2IVEZZFM4SBqrsi0xa52hs2kelc3iKJcWiTvU3X
0fJP9qNFuIjXBPPZvEYwhVtIh6DwiIC2viSscQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
aaSlSwNJkkb0vhahqqItym7j815+DDWdbjrFuW0kBHxxgCpB2qOcPQvpIaKa88h9gxc+xnhZhIJR
bFTasXM7wnGbhlQpyDc9zScLGhNlmmtp/SL3y6UgTCx6z4o8SkLPBxAGDlSl90NlRw/i78jkeVTU
qcE/0MwlNDSyfZfS1UBNxc1y0Fu47Brq0eRclrZvZ6XnWY84x68eBslZ8eZCazRxX8cnN1naH+PH
I/7HLehK5L6eKFbUimZQ/OSc96TGeMEqYI4Y7h/A+trtbTjMpLKrsTcMP2VpEfhbsMPdfDa84yDd
Gz9Jz//pCPDWDwiqVdxB4JgHQ+eCsiEiu/7OARemvHDobyYGzJYjr/a23lY7eC/VYISsfFWl5Lg3
HfMcElk6408ucjKFLGMRRsMaZODySrr72jWFJQSb2c0Q8idSez0/+Mk7awlsh0G9hzVn1l0F92tV
63ecFYAxe5ejSbi47kenA8p0iZBy52vmR71CIab//lVQ5HcLNXKSjF5SBSRrGD9XStur9nLzf2uq
/nH9QORkLeU9Jnb4rglfwkYgJpnhrFyNxwD0HYs4aypYgzQTfKjL+iIbvfUTfzVFlz6d7CkDF1H/
KcwTmlwzz1Mvu1+YmEcqE1BXfZ2EBFdS+AtNU2MluQLT3nR2qx5OpZ5Z025WN8Rqj0Dw5X+SHPnK
KJYvIN/TnbqV1GxFANLV70unGggph3obVUJG06a4XPTc0e5Vi4TEL3fKtDb14ZhXpIGhnfwJXZxq
g3slYoItu1RkY7Cq5Rr/aVWQh4W/MpOWgJL/iy8kqy9ycZZ/uTbIDJs+O0T8NOpAm0M3C/fPAkEg
KhRGXUW8GNG1K5svqPyQZ4h9lViVU27AzzMHC6NYO7In1x4akxAEQzhbQXifAnTRhrOX7WFxKkx7
oIYT7vqwPrB1KSPC5B3mHjzr0+9pIVR0FazqYC7IQqzFu7Ubw3wcIxz845N5MTKlelIR1cgFHoJM
b3Ri5zC3aq42nu5nbX20nd8BHSheiFFzYnNyzWgNdsg4xhr0jQCkd16c4o0KT+5ZtsScEbU6xeSa
D/RGIWHQI1eWzBvcS9f+8YV9aebxM+X7ZgJDQsWt4ye9Vz+GZd/QRzsxvOH8xRBDP9UpxH8Dpe/O
IqQoTOpnQm0ceyMY8vEPhBIsw5Enbz1b3yDnpFJtHI34PPvY9FZ+FKLBX1e3FkEKCq4uFPVLqZVf
942LDbBTWPZexvmacV++OKtVO18EoZN9UDMzijxTKNHMAKCm3KY5WjieFIraNfxNfTam4w4bIXo8
jCVOvjWtapVn188IlW9uFY/pD5y9XSQ2FKNl3WT/WyLIDjQ4ORaLuQd7ZAs5Yqhyh7xdZvjlGJGJ
zoidZlvSbOa9tcHhU2hudySY7S9PXJgcFRB/9iKGmqmt69VMeVoG/nmCEyTDfpnJBmAnmcmts7PP
b6EollMMHjLzbdmboV0AqsmTcZtuZ9BnKdmd0w6Htpxw6WiMs1w62Lj50+Jm2Uu51g+YzREvmflr
eQ5pU78HmabJc02Xrg08Vzc2Bhw03/kx3ecJp60qcikcpEx8Yc9ZQtx2PT9RlB2nQvUFWbOZp0Cb
tWuy0GCibkXHIdRn8URWu1F9ImvuAllwzxUVq/9tyhhNJpUVgAxqObkXBu3qaEZnDU/Xn/DZ+H6k
tMx1Yx9cbWL92FV0Qs3ArIZKJlWdJEd/7C+uAahdrd8j7qgX5yegxkuHoYkZM3t9+dHMrQ78i0oO
3+LzdfiUwiuMs2Q8k6VFcx5Ty27N+MDhimqsPQ6RaGLZ6v1PCsYStuI0tC5S1bKcTCLE7cHDb0aR
eP/IFn68ilqvosifl6e6NtTOsXKdIVII+k3WvBEwzVrHsyK2aUrGESIQqWtNVvbq9UCTVmbpdgGr
m0vIRKcA0WuRjhLQSOG8IuFJxwWNcg3i06MkAw+z/qh0bcQJFlkQZYCROoUOQzsY6UL3EK/hpYM/
JgLx67IYIhAPLdJq8keN5II0tpDWqhOsVMq7hq5YMQGno+coAXw/I/13K3wRKXhfzrBxZ2GdNemB
NWIbDSOE871z/kZLtx7vy0eHl+35h4K3dt3GiiH2p9UauQmujQo7r4F87Sd5lcDvjPDttjwEwF/h
pJJ8RigJNaiv2tvbXYPWbwAtHou0xACSJ8MwSRS8LTf5m+uWhyj8NH7WoxSqEF7moH3zEOaGOT38
pE2HMt19m//MZrzHVw/GSwb8YWY5w/O1V2r4f6oNcZFcFclBnXZ/a7PkuOscORLfvQnf70tkn0+o
6VfGvIqiSAzeWcWGALNlh596WBhVoCRd9uCjGJrAjBxwkgTqZd7VjvNtWv1rQ0WS0dda0BVapU1Q
fp4AT8Ufm3viNb4XI+2hEBOxmeIVOvv+Y2diEw13rGlKgYTA8AlK1oAqfdQja1a7VTmFyhox2Oym
jzzNfAw3dv2PUmdvI+f1T1OiVwyt0UCHPHIbZusF3c/Hvz3JlHN0KJgq/yXwz7Dqix2uu+HE7e8X
LcWzfBvBWmR+Ccqj8lp+MG10Eebejo+WsvksVmJaqc5LzlSMlVo8Yus76UGIEZPdDhPK1R/blOOO
3Azd1fAIRGfs+XAxfbsb6LIsRS2c2leNW6peB52ctEDviJgX7GyQq4wwZY/tpCnuvcVGNsnyw+t3
06GOWjpG9RvlU765DfUWUOcEsCC7ZVQqwdVpVumzWTRwZiS4z3eMoxPDBVcuZQZslXfRqFWENwxB
qdmtlpY/Je7/XJoc+qqp98FKRCGydBsO3tsC1E0ZmdlrOt/GtNCTMPyPKxhPpJBk6omvsuEYTSTe
JS1qxfqXzK5aysUvfsNTuvib4tscoWcbmFWaFsNfDn36sUV0/IBGQ5fIGpryCbpBeXEGOnUwPBWF
K8e62iGw3gT1DN2dY3dJabbo804WRtatRRIWzG8PLcWaiTNQTV6onp0Ta2w2QAtu7VSGHm0NnPm8
PZ1FXo6AwFRYMWCycUSgagevn04WJINbtgeKMWiVwUpRAFOWGaB4RX7z+fyxUUl93Mk0v7FIgNvZ
OKdll6cr4HqNuzSVWckmSAmJLFjEMf6KxJjAHuwklE7dSqaf0nT/+QOk4yk667wgK3SoGKpNced4
NpYim+6VgDDlF+4ZmhQPqM2NkbRSlDdTWE4a7BhBg6u5aFLf1wtgXD2wdF+uNr4X6O/iJl2jINnb
Q2b3xFDxKATNo29+uOXuT5ei10o/gp4w1M4fBt6OI1BDKCa9q4/tHndtCkXWVD8Qyz7PWKLDoZe3
Ts0/0JwBG9IMofs1+7BsjHnQ1XRjce2IZMEUQQf2B4f/nrvvsFhvhZTICyVe7zmzWOo/FgUkISa5
9OnukVpa7D3HgZKpjW2J/yo4JCmhtXKZhrvTLUNYSBG6Ei880VMkmgK5CTB+3hRU+jHxsOq2gBPC
HpsJRCyUaBKT43zGvJ0DSDbKRmZTldp3YeXewkTylQlhnKkuJbRydH0uuzb71ckzvlyN3Htwbn/g
fIosbhzieUkSsWMoSdyXoGoWfEunxNbkCPOcc/FWopEa6QHEcT+Bv+huH1nIt+LidijavG7+g4Kk
Lrp4HJiQl+hL30jizIPJe/Ra3rta6uxWBnc6+vWX6WVMNQgdhgZbTXf4w6tvFvvEGKr4Y2tBhhco
pQzdP6K+i7xq8sfta3BiTcaBuy8jDa+6lXKjsk91rPoWnwx/PRD2Sk5D4ET0ZxDjl3Y7U/0lxJVW
htMyK4Xli5M0/pv7Tsg/FkJ2qCbRabokYHtWXXp202At1iFxOxzHVy39J/inoj2bV7c6QKa6IZmb
iLj/U/mfy3Oe4BGypn10Zri0IeigQpnNfTf9hS8JBTXscmfY0oq/MrgCjd/Ghe6e34ZsKu34ZHT4
zAdn+i0zg0Y63d03rVu2IqHgO/CwDKn1toPqdpOjgoz79UB6iyv+3E05mmURfOBH/5vId2YOMRiK
nTKsmJl9oPRTN2aY+UqopaU9xgIxKkHBLRs2buPO33uMZHR93GeNkFplFHXX3fn767G5kG3IJD+u
k318f36dQ2nTAB9mOZsFsgOkzIlD8TSSxRJdkQ7aVUalYItVnPHbk2eurrcyDQlTS1bOsGjEDyUX
rWi6bGqRUDC85FNftVX3jjsDfb+HnzdqA6SQwevoNxPV73483GoQgw5mbyEEog08QN3Cl7vLjVL2
H6+m79MXTYvzo+2a4W88YDSoBi+aD71xknipVNE8mT28HLtou3dM9Wk16eeJQHpCprLOTlbeIka/
wZCULJ8hqHR+7V67Oj0CHzxlJdV7nT+YDZnJR8l2Q/Wv382DzJ+w3+UbWB+TRr9sJsIcg5YQTnxG
LNRP8EXsIh/DWQaTrRICAl1Ra5cQ6bIsTuAAu0OAhTnnmJ1E3nnArUoq0BBmwH/b+wcwjb0D5WGf
/e3ix1klFIuTEZsC2vC5RwEEnpOWWMV4h9WL9LOAqbFStj/lcsXdW9B6eMTbyMET6TcY+1aR/b/X
KwEgjcy5AoyILWoc8PXcEqA99cYgC9cKhoUKLCfbOuTVOVYq269a+IbiR8fInYrdPHHZT991unhX
FGaYdMxm1NtXzMps5+r2U51GR2J/ymOXJ6uOTJ8mdUXeHDNmaiE/ghoSZbShF7V0cWwrus+0TXSx
h3UR1I3OwY5/GQlcG/YEHOOWLObk6ksKAzDpf7L331yYxOSPaXj322B3S+5+GpIRh7GFqg/XFaxF
RfLO1BQVNDgrz8WAivTh55xR1ndOedLFPInoSbXIOLFNnUFqx+lGZ37tFwZA9EfW2OuS90Lbiey5
yEpdiXhE8diLSLUBR+JB1QAzaTFQDvQQXoJAW6LzTYb7lLRJ036lXxHPF/X22vF8EYQGt9GgwTB3
0/qKZlfdc9i3W/OLnRL0b6GR1lQBvuakhlEfqK/uiMFiYLHwMyZp6vhIRFLwqJJCaNxe9JlGO3or
JmS9p5zNauTfem3BAI7i4yb6A7Y02bNWveaJkDcHqecKEsMQsr0JUFa9pu2naApygNTGjEp8NhJp
ZxUBw7/6GfRMbz+AlKq3XtpYHjBfHEdWcdXtxwkZ61knX5A7+lNDNMoHmdsCoLekw4EkXNEaRstS
KO7ZoEoGnTkE+RzCVZnLqZu/Nxqlem7dMWeGDMeLyixD/zItPxFZ3JoZWWJWPKYpeT+U+k5kRnha
191N95QHrqkfjWrDsCJeAmeg/NS96RQuVeWXZJItA9hBLsWd304sSfWh/KLkxNxqLNkIUdg8blVi
UdR3K0ujAtD+X+tTCZdzZy/1SpOS/FjWb66dS6XHpNcfmvkZYw9/Dije3g016dWyDamrBD9sh85I
85gZ9TEFqOJ+saneyqDdZKY/Dm4ndn2lUspwkFHunyqSmFdmWByo/uYRgkC0/jenE+gZh/bvnbKv
oUGmQDnPDZa83rwN27e8ynpArw+qASHL/gz66eUVoaupQozI/XUaVne5r/sblKXEW8p7bNQCBt21
D72cqMMdfxlnaYzBsKt+AxuOy0r2Lhpn4FMq+GuMV0NoLygWpt2MoZEw2fBVYX2dU3AE8YajU60L
/flWBqfX9HNsYGkzlwMDlMcWKuqeJtjh+B59rNPwaUDBQ7NH9fq9XmQzjIDcc+ZKo4DSnwAlRATd
3ENJtcztLChbNzx/CaCJyL57i9MdV+FXmQYvWmU7FTBjB2i7KqPMsKh2nC02rqBf1p10x0M6bo9o
kxfwTWvkYBpMuKA36+b2npDbjIRoyCy/5QxezbH1yeismjulLWf9np7ZNlBZHzVzX8IotHP17hyq
taeEvj21dVlOCHCM4c5aHdfLYDKUOrrAGG7KB1qD02LM773ISMMvrT9nRQzatclKV+dBapaz+fOA
eLxTTjWQ+/7mMNqGmiZbG5M0d0byUaD8IJSFifsGemQneId0xhw4VMnRYmxLLB+yN8xYC6usTyGQ
c8KyiGXel8NF+xTiQrqxqlXHz58KHVIYqZOD62Gg+Sd5aCOeC3tNYrTVPogzZEpC48anmMiWpSMI
UiylBJh0OGV3bWM7hWr9xVnG2V6ouZkEnsXI+wcU1/me2/1RNBy6bUxVEMfkQggU1cdi+9YxhJz2
gniDnercu02hUO9FmDe6pGdVH+lYNsM+e2OdKEOvXKrobrFQQDEudvZ5XFEh+X34SFZb1LaIKaaG
V6vaPIw/KCuJY3c1gDG5DzMjn/lbgX4NRk0r7IW1xwr1SSGdO93kIdd/OUYgbqlNycvU76Wr6/a4
v08zEo528FM3g1EvU5iIOEYXqioZBotTEobg/JJ8B1RradLI31dqszvn7SBcX0TFE+9zvMSY96a6
/ro1836w349ZPQ0xDrgrumdtsCUSTZazxn5cJH0IkNJ1+ngub+KLffRqyeuKXOKRyLoVluh7tO36
1rgmFOJIg1vruAIgJBRIdROh6cAaD58GrEMk8HPyyGCAKT7wHnjNSZoGyLTXBgqdfBBcgCj9FL/X
Pfqq/9dLSIWQtX39Yz/AY6d1pQ/9RgcZWZdl1EFzGkseUU/0IqrN2vansB5VLVRfkpM/KuJy2/Fq
VTueCkdErUd0imywxgdciQNap6MsrdkSprjI6T3wLXAJPXcKCmqiOmC7KrJURQGBhtGI6ibKTyJ9
VYp6K95qdZFnEo4Upm+mbOXvfZtd6FG6v7KLpfb0YDcU0ueratY7QSxWpDiCVvfrndx64/A8AZmQ
1ISPXnWkl7GO1CjRo2eU7uf1cIWP4yjbNjcKK63yrAk6YAL2lYe1nEgK6Kg9w1ZDnl11BYN1QUjr
ILRcK8Al8BUpmgfqFyamBFg1zi9JDTapcahBuD0kPBM5BojDUNHCC6mM+c5r2HcPLkEIhP8GUE/q
TOng+/v3rgq5i54TF0OpZ6Gv4rKztON7fNh3aT0idR8jkeTtgtOpMEstwG0EkbteQXoAFXy+yI+D
Lb+Lm9tHZakuHxKqUfbaXalcBgr9qZzsn9h/zuYFmA2DihaX0DaDCmT23TTO/MAUZQJzzGNKzNwT
yTSg0TLf+jiKj+xa3KbRgAMYsLp00ny93ApE2JtoENj7pty9uB3/oD7JF18b6QhKrmcqFaynU0Z1
6vpfajqquy3djgaXNDbxo2O/5i8qqAA2fJpkZn8fqP7vpAE1XGyM8dBc5IdXrI8WifY96aB+t/Dr
51Zw6hw7XLfEWJij9URLi97BY70xFoI1K1PqVET7xTQTvaQ3HSWMUOmm4x0+1y54vQOfixIh9IRS
SngqhCYKRxNeBLa7meQ1/s/AhJwuGDL63jrKvi7kl1E9FZ1wAvRefUR8NiGn1sVtTORO5Tun3aaY
hyWvP8FkpQ0md9qbvGYm082gVzhlJ/5KOtYiv+eCwqsM5nvlsVWJBQ2vRVpPAfWSXNDQ2ai2Xkyf
OnFQbuAcmb0hT3PdtJmIxQD+AUKUTTfgA9oJTRHOFYRIl16bYSYxwLsh8jj+P3+4wMY2ASaC88jk
DRbe8HHELr2UDy3ixGWixAS7VWDGMUodk/hP9iyL+EhwWAUEQW/EjBob2yYMC2wgh+wTxt82PqLN
9HrM1avwvOyn1LcD/Sjhn4MTDwSHmhMzVO19YxEUoFBgAqBVi04vZQB5xtUihAOAIkDwfwr7lvQd
uQdMdU9ioWuHkHWIZC4/EMYNDQydnLWiCWbe/Ky8ciGLb8W+ypS6Tcmh4pD0Eh7CoOV0qA80QI45
EcRsz8emgqSPwcy9v5s5uVbzhRgoz3yG+fE5o7EPGYqdwsx03Db5J0RXYOXuZx75K7jIdumokYgL
Nm4iExJQQ2unCWt4+GcLNrfvE9LCg03ii6qynyPv70befvZWulU3FAMSU48IZ0Oh1xbT7vbm/Qx9
tV96LX3EyHlOryCAOkkHJqxbT3h8tl85aiTL8/9hY8yhJMIb0DKDiA7pDBYZh3rMPzI0e36cbgAh
dIFUvu1d7qlwk+m+oztkG9hQ5HjGv2x6JRPDtWYAwTvxJNDSkBEiLb8FXw8DdrvlZnJClGgQ0GNO
lGPRvAgSrtaxakuA1Pr4eFJxcmJA5QUkxCgME+lQPVfIM01beX7slhGl7rqQ+FsLSBevEPM7zAKf
HV8DvgVmbACJcqFm29hi5TExytvLlf+tD1JG0kUtpD0ShTYUzRPCwZxkYUgxynv36v5nSRy8YWwn
cGrwNV4obRfRbIFbJmyAbPjauFg9xOTmVyIzffAqb5lCa1vMyokZ8fDA6j67KjhWhDdE6F7drvGX
liZ+em876EX68WgemFvjwYOBUnYOR3dMQrJvatel+wgK0BRG2u+GuxM58alGJDfPky4TI9fwhWn7
p8sQAPu1UlS1EMcM0zaZXLq9OV6Iq9qEvZMVTlVRcecAwLFjEMw3znJRo86BSDisqWZdBmzFaxIK
ku9SD28UoQJy19kFbq2op/VKqELk1DvcYRKxlB6Tth7DaQIwgIPzdQbvqmw8NtErp3eTSMoYPg5C
es5GZ+VH3aHlaNjmK+rJmiGF3tn3ypdUglBFQkwptP5OiNWxAUlJOzWBuJ8tBNGZpndMsmINvqrh
Tpy1ZL0GeVGrq1BfdTj2DTTFvuVpK/0sXGg3rGRe1tBHMElifQjBtCQ89xZsO+x83We8WktPnFsv
oNDmOmd8QMf/U9ZjNYLSQ4yoxHjiEyEgYm5eEo8GFJbbD/JVrR9F93ORpdLuSE6kM2n31PabARvU
gp73LuaJIhLa6qtvhAC8ZJ9ePTl5L/4PDvccW9rW5/1cxpTONGHEYxp4v2pjjzt0rIW7h7w2xEoE
t4SxvUc+nwjty/mJctueJNvDh6tmiTLIqVyxe4UwxWaAk61E+hQouwTWMA/KuuoS2/WIrqfZ8OHr
lc1ABV0sMqNK9VCRsvaUCNUQKPHbG6SHTR8k4fA7THll+YuSyaFWS0HwKcBJITqceSxjRUuTMwIH
xXek6MPsc+tfLC76H1BTHMJAr33juZ7ZWVpgwJLWed+jl8kv8tpa9ev39QxnDNUx96KJ4QbmlJGY
Hn0VvoOJKQ860v9JXD1IIlct7KX3wrXwhxax761BwPdHk8/Qo7N1JnshbDXyhVyI62wcje211lgC
6yv2SYhoULu5YEqJbUX/jaaMZzE1FDJ3kMt+xsx6xUIGtpxuwIkdRdyzqxjHBG8qqmoBw36mPalW
Nb8upk44x2wIY5PX5PFmY6bRreZ+LXNp3ljejWrvm75GAcsDRdpqtNQ4kFlO/DFuOZ+I0GHCg/24
2NtJWHbKN5DG0/rEY60EwnIgaDUwnQ/ta0zTdqZ1c8RvYCL5cr2uTjiQVDEV6Rb3zmxsyLy5jf96
J+SVQexOdw5RgZhudP6rNlfIIqF3X6GNDhLRTuSqHDEQgJjMjWnQTn0DDvsiGWLmplj1SVMqaG8k
bGAz+l+8C2a+V8gQ9HVLzarCtfi2URKMRW4X8EwfO0daj1PCaTqk4/aUtSIt74t7QQFqOduZrwOI
Myvd9CLgRPss7+PhYDQ0pHaLf7j/Q0IP6/6LpTQuMyoEkhkfJ6AtQM+W2JvouptYFDKrn5gH/Y2g
x+qkThF0COlBYSt8iP4Kf+ldVXmabHE70t1sACvpKnOVUMsf1IXTrD1J6/BIkxn9ilFb/oZjG+49
MgHJZthOaobjRrAG72VwEcPf9Y4WYGBld1yryOZ9dXJcM7D8FccakoyLn7jQbRkhmYSoP7P1AW+Z
SAYpNJ2U50ryyaetU99TA7PG7BYuG2KH418Ez+tEJPj7V+64ZpDOQCpedWMi8NbAGaJx8JJmd0zS
UYnh/tX/5c4g731PH4I6WK5t4Tab00US8R5bRHg1k+mYiH//bwk832H9UfaaalHpJzINC27QlvKM
El77N6idLGc38FC3VxJ4XGIYSrtFMF4NrUMIDRx+9PqVdCQXUBGV701/ruC9GHJB5KfJ7wzNXLAo
FgnqxVCNncDU1aCK9ozvURLozw8BqKr0Zrp23kFfkA7hFVn6aqaFlqZFr656kgtsYdPJZIRxLrk5
EJBAijzLSbPVpCuGegvxQ9ID3Iw3MikapodhLQINeJhyIGOW+6WgAXWttDfZe3202U59bAH8eWgF
faLiMSKjz/LvRk46r14OBTvG4D1WAcrQmNUNg65RrS1Qny/sSD4ugR/gICrL364OIisbtylKu2Ux
P6MTuEYGSSw29QOsCVH33tlHeeRk1/KuwE7iwIL5Arw6Zw/C5sT7jaosgbNuLwCgPEnUWsMrwTwX
AKczr5pvloSsEpdd02oqO2YfUD4nY8Uc2xCSGb8F40sNRvCxlroTCDHJgeWketlh4qkvLAs9+eq9
i3IQbDHDUhUFo251uQG4h+EY+jGW7RXTgQsJVKgdg7K3YPRaH3Wwk4i7VMuPnF34tPoUp7wAbxqX
tMXopWvUZ+ic08nsJR4Jd/+Pmo2wGMmhRG/Ki+DWtWWE5RD/zWe67E5KwZnSsC+3V86N/WU4gANX
k1+kKT4vwAD0hPgcQEVmqzES2CujIUgBefeyHni7osJxfyDixbWVQHSeVvfu6HCsZ76cnxBofueW
TzkP0A4qqS83f6ixWhZWo2d1ZrhpKDgKA5WIFlS4ModP+hu488AetZwzjH9vj+9s5NGAnNW6Hwqq
VuvjIWxVhlbGnaXnV3vsGkzWRuDdQMAUE+hdPMZLNSzFjVlesnfcp+bcviK4M7XIw0uAb54dF7m7
D5BREe7w9uu/DIBEhhNfm6co0qpwWZytDItLHpWSYg2Dsx4sfe/x+PbgMDYQqD+fV3dXOoNoJLcF
xM9l/b5uCfmh2PiOZs6fhZMKa8kpG5x5ZsSS2u0ge0+9kmBwQUEXVmuCpTvqFUMS7w7XC5CdJn7Y
I9trMVG6xpLeEMjj/PecVjkgoXjJqNdj8F85V0CWcN5x5RHf9IxmWPTwgI+HmTYqF9pBFJSHQfwe
5EmsbNmUnhGRJh6VEVhwVO0rMnF4oUQfBTSwRRd7ZodJiqeKGoMOPieGPzVQnT0YgFnv9XqBj8jF
7auV6O3o95e8ialuTFxuIG0DtUcJ4aOp2ddRbztv7a0rCSe0wAEX0Ml/3QcS0j3Bq/YrWSjgfFtT
K4LoA4aOsxMw76mWoaeclaJErra8nHaO/sNTBryPA3qNJFP4x6rb1klsLrR8tDtTAzlV0ZQe/a07
nLv7v5MiLX6tp4btHO4ReJkUNM+p4a6b/q0OZdXJHvFXuGHyusZhgiXNFQI6xB42Aj1KG/QwN/6k
tS86e48owtkKgw6ZFfDiyVI/EM4JnOTHPT0bAHuvHaI9P7rHNixbBqHFfBUr2TzoN04cu54aE3rr
U4J1mohBkflc8o6KYEpe19m97vXFnH9FDvfirO93izH7dxXgeGzONHR2ahTJ0mkl5FkEZLYUxEsm
s9FCgXwwUpsIVWNDGzNYniWJnEQaV7hCq4t4gQr3FWIPij8RK8DpwneaCOeloJtJII7xLcXi6UyR
JkVNUchGkMnodwGKlJpYqvmWwo7N9QsxSnctrQes/Lz4PVJocLVfbQZuwi5VfhPOtRhkYVmeahXy
G1bh7bzAKNEsbTW+HmcfwMDk5fsd8GizcHtp020dKh/va4C13S903hG3ZSvC5LOSW5pnjYpgCJCJ
2+Y8uD1l8C8NnBXfyLw2Tokl8abJXoBByCnGJrt0Z8h+QaFno3rpR1yuDdgjo2CTVsEOMkeWDIdd
XXqtsF85OZwln+biH/uVaFDIT0oDLjUg3EWR6zgK2BSp/yffbCPeBUsktES3IGgdfXBFkZjiKDBG
Y+XJInSU9Wbkcu8+Djp647F25htBg73jWKttXdLBgt2pk04mvJwkDp6wceJaTzZotLyCaG/U/lDJ
a7SKSW5WzU5zHDWkbUKquDmQtWv1xfTtOzaICM5IjWvY9BT2WQ22a5Fb6LIkvfPkilHqvauR8/LJ
vburNoWz1+pIztzKhX8maxJS1GN/SIP33CeuEL/UvHFxGIlqxYmC/ByKS1dEqyPWS4MtFOvj3u+c
r4CH0BpU6YLe12xoD26DN/+iinFa+nD9DY0PVKgKtXCLZiVygEcpD5q1sdYIGHh/QG6fxVQ/5csK
tUyqhWAOjRnX1H5CfmS+Hki3h9F+QDDYCzlmaPFNym79rbuHvo7Bv7N5VUgWHDQyanwttYPcds/j
S9pSiY4/La9SJjXshsavrPvHzn0dOPJb0ijzGDeYv/0SQCy6nPvX6/WmGtOQd6pwOTkwI/OVDU/I
k4yEONGW6w/Q6L5N3Hl8hOgoHtx2B9nTHzxvysmKE7AKz43Eizk5g4ZRBnSR7keGtvAoe/nMddpY
ltWHtLcO9+6Mah568Q2cQ1FmqgJtZwKGNDAW8R8e+Sf03Z7MzrMNhMFWPzPCkZJFR8r8FgYWlJk9
MxVaVhRQlD22uhK8Cy8o/EYdlcM9nuVhZaR7AEJJQkgc6ULROYGJNx1UFn5hC4DtGQ0kh8utjErY
Z1mDJ2/ajqJIvwTswBqsphOgjbQLA7jPS0B4rckXn5WtLfXle8TF3ZgYgq4iPcPh6z+iMXtrIrUX
DIF3BFZSoblK+vQ5APskCtsFDPxLYmftWU3cOCg1+ODCELwvZAmmUXVyozRTvkCJYmauutOcmXQW
RMr7YEGnQ4S6j0kv+A/gSGjfRlDLj09WsN98gFJiZ+J92aty2/4zuTO3892hGFALwnsdG4kF5Nl7
NqAy/GKoflMzsR4SdKijBKFvk4HX4yB/Hyet+MhF31S+fr93WpdT+ANjt5wKNMWKOOxNXYORy+t2
NtX6v1dIKmev8V7Vq1gD2aIpWIapT85L2CJB70Punt3HnU6qysZlqL42gu5BFaZSO9SN6rBRsUxe
DiDGIw6veUnIsKUKFIZt8mlYLuRhhWBOM3kk2KMi76FthEEEfGfKJ0qKRDU+d5L6j59ClAfHxafi
9wz9XPEB6cK3Y73PGpkC1838w+0C8ivBi5aPebNKITVnaGQbY4/DULQWXMz2p1/fIsY0lefM5rE5
KStqFUaqR09KMQ+nMr2Ycp8D3SFnMvHH4FFWIverKgdf3Q+usmJT9gFUg8afLStLPCAgZ4x5txox
3WgzpzJf+9b/Wy+REjJcG1JDEFpbig6jyHoKo+kC6vKn9RCjupYY5jqeCUEbIWfL6gWLJnlIJNhC
tr5m6ffkbXnPb3tFdrxSRCH52In8vhicJqvLgJ9kx7c1CFK9KekpHas3vrpODyIXkxwFLnVtiK5J
q59tRHTklcfhuK1egqhabxIGbNuvcWhd1+N98gVFZ7LCNBw1AtwRjIfUOCDMlF900CUmUs4ViNRM
jc4EakdvgKMCJkqD3x7xepU/Cm+hdP3sFExGnQy804k2bPjFV1HhdNQa/HZhDWnNHjhUv0wipqM7
QOc9UAXyuVbtOxfYXMDqGCLbw4zLfM9IN1qAYee1L31R48+5MiZtj3bzLF8otJYMN5xlDdgZYKmR
aypiZIgldeKVXfKoFgGWNuOuSxnh9bkoOUqaZW9niRDv32Bka2QTq9PXl0BCxibf68y5fajCoqGI
e9n2qagCnUD9EtoHCDQT16VlgE0ARVpkDslPc2zjAYeFzhoqON+4PjRnvDzt24O8JZHVZmpdYuMA
H/sPhzJ1zSVzagRzKrIrVq152D1RjeWZOzElHIrhW+P1BAeh+W6Bz0deX8m2TELVHoD1AZNvkIJJ
HiHOVwSNwtEZBaGjko1Qt+WzsMYTOnEOz5WwYSO5Lv6J6atG6WmDdAqUvu+xZnoC1agbdiX2bS54
c7jk0kcGkuUIu9ChBmJG8Cn6gdyCg33rjWjfH5UnMx34cJpMG9c3AzmRKEs+5kLyNJDlh7iQOv0v
Vd/o5evAVXmHh6/ugSG/Z5UiJ73uYqWVo5T49uoS4q7J/sAjYj9RGn3HJYQsdCsHna925uEDMxSa
s6vVecL2/wTfCgHjrVno4d/wXM3U11U6dkvGTiOTPwBmFGsG0fNd0LfQeAOxNSDL0b/kPSEzQxbO
WADrWtwo9cYs36VZXQiDLenG1qDPAX1wZzno0qZ6/H5kX7y0HJEobFoz/EmNvZxRl2X2ZaaR4fEg
F1RoW+UQQ5dZzdoDqKvEtrdkUg6QIh/Oie5TtL5KZkz2H5dkeVrcGGJdGHAPjcO++Vdt5uBh2byS
5uq6K5kU5S8kQ6NbVG9PCtjVN1/k/6HQDTYKnxUkBkO2H+SQDXVXW+0Fc/pW/8lMPSMJ0gcC42Ee
R587X5BIvtvY/0ttfdlAkjshU+tTXvgtGHtjj6NVpUjhqqhyyTpt5yzzgkPOs+pqFC6M+Ayie0cv
6EFJ1RgY0UZkwh2aPFmIJvuvfIHZtRb/Ke+qxkJ0fhupIvu6L2RL9JycijVQ700Nxz0JeIDomVEy
63rBa0k5xGh2ZNOUZYv/tuMpwP71jOrbhPL/o8RK6Nj6qgiYuOZ92SZHE2tRG4J6dcZbTRVAsH16
vCg1W6kd34h1OKgoM9TvpLD1xkCr3QJX8G8Si7xnh6hUH2vpLrho5ONC9JE9IcHfcHA6H9S2RS0T
GAj2GyuGVJNA4LBIv4LVu1rXH5MafX8C2//SfTMvhdn5XdzVkCs8k1fr2+3QorVjCmZK0Jz7SO6A
YyqowXNFNi45VwuqiCgpLH/KJP8inR7puzQRAIm/bDwP1hAXD5dy9dBX5sfg/RfalPtIDgg32wuz
gCMoF2tWnoMptwNYOLcY3q7LZKZgQURRtvTGCviOctYtA5D8X+lGDhXQ91pBXYckus3ILWcBkH2R
jirZ3GSuth6ZRpXVyxvB/wyKYW7c8IG+QlAzD+2cLR0lOz5ex/Rwu7Xh7jK7bKrdSv5M9CzNSNxe
y4JBkSkVKQY6/w0L/83SheP+ZAf/xtiJLNgKNoIuKPVxRQpAGEBNN6WEDEq1/VrYpLLFzYO6uk/O
56vVRz2Ia+Q0ZSoE6D/QbMwpkaV+Bty7qxS2zHemLc9+UnbATJBXXzz7NIC6uh8J6rwR1UcS7R29
nITbbojTp0YoYy6gFH+BCT1qlWrmrCYllQLpXjhTrPBvXHQzgtuHvwCtFVBS34LBlUkK8s38iM4A
1rQxHTc7SqPsEvDXOISObhY1vIO8jBkRadCbPtOZZWLLS5IWSkqIIiYeeUih9ipemhupol0ddum1
7ZzieRjTzTH7lhN7Ub564m/FUePitAPXf3l135NTo5dldevOu4WNOfCl8V9hVdwf3SxUYoRb3YA/
3GiFyldv6CpiQmvDawy0EHgewRvnN6uMRe/CfCHCQBQwLV3njjixkJ+P2jBjcZexhll5akLRVSLt
eQVQiKjN64UvoDGFU3adPKIdjhlNmj1SFK3BLGgi0K1wYC5ZVM0d0j2VPRaTFZLMmbEv6ewKt3wP
Qe9git4FyI0aeZF8kc6awrSIww/nD7OzhiU9Cx4LfrRcc1YjGgSNRfUHzXGF/HNDLPixx6xt2CKo
Amp87nJ6oKhHGeLMK9bP0QNa1ylYbkKu83CpmpH3laubA8xUMzP92SAj4q3lPNUq+wfFySP/zliV
HcOduUa2dGZR1/e/zycO7gwmx64haQpCNLjlKff4OdiD/UlDYnAvly5VqBvH8CKaIZ/OztKPOo6N
XgwZU4DDuOfHyad3VAkwRC38FEeOBbVbNe53PrWICuecDENIbZL+hNGIo3JxEPS54Gy104GLgZV6
sWSKYQj+JrtvRIg4rrzf/A623IL+4gCAsN/MYyrqPIpZ4Xd7NWzyIAywfl9JBEhqodBo8uid0GIa
gPNwIKHqs4XoNzRTkTwc3QUl3z4r7Q6fK6tgzPbmtfuojpIqfPTJogta/NGe2xbWyRhEEe+p8PgN
XiaZUunuA32Q6XrkT3r/EskW5S7uYk8VUzKLBX8SjDaiY0vI65vpqlFH+Dl8beEBF4Jlx1Pfbdy7
lSYb4xU6AIuh9Yp3YpYUCXLAG7NRPS3xfqqH/tVzbRlzl247hkPqtegjcW2U3iOWMUSPhNdjj79t
BgrFkMAfxSpC9oQNph/zA+PR5bF7Y3qxnrGgvh6Nj2AkRD9N21VsvpzTY9qA3H79f5nsLuQmCVI9
dUEa5VyrJ3Mt5kv7olD88y0iIaeXfKqcS7qA4C1M7Kt5pHMgUkew34bkUo5EbS65KKAgETB5nnpJ
isc2gmy7oBwJ5FdL6npetKB6wQL3C0+WWqBCnRG01oMO4AmBirSLtBQL94ZV/BLXqWFWgHEIF5Cz
lIzV/d0GXZYj2jfFWbh59+rr5mTKUcIm+D/8Wbq0gahq2ROuiXQ3oBY/PuhKGqCWfp41kJxLVRBa
GBFQAN/WXDxq4VHgO690oC4x9m5kaHhwFwKIlICAThW+o9RzqfSx6NSDHGnimiU73VacjlShFK+9
pyTFDMxLdQD8SdSmgqSrprpfgX+cQ6i3PIpUfRYZDQIwJ9f9oyQ8qRbP7vzKAFsTFUa/CimOLTT1
Vglq1K5vHb8jNf+Y15Y1pE52HxfvF/A0/PrmkFld+Gvcbr6k/fYlqcL2i573qvLPtjnCur9LcwXe
b1uhDdtelR56sUPj+3gfSYaLYvFacp7PIZOXW1wpEeX7/BzdJBgixg6Bpq2h+Ux/VD8BXe1up3TC
AtBBKbWf2ajtkxhvFLyU+dYKLafjs3305cickMJBRuzXWlw3Kr1QbdD3WGUh1zOrq2nA5eNyislH
/Zuu/fRhrJygPKKeZv03JfNvibF15oRe1EUwV4qjNgB7UwW1wN3fcYHdeJFjPT5ZW1iqzTmUV//u
TKHK0ZfdBx2APICc1SuNr5Jiq50YpWej0hz0Q62SVe4ZjaLvzuCxCvoCzEatP2qa7tBdw8gYQ8Df
2JqgK2729bNuduJsq5Zw9UCvFOxzZQGhXnnVG49nL56y7Fcsv7OkcSWy2EJDA5fFurYOhljEwBru
pIkbtG249fYgNTERpZaaPsTHrVLTieM83ibn84xg9VZdJKD595a3lMMddg7ZcYln3BN6eK82rGsQ
qAyNPjQTZbZsMGWC5Fa/j/VNTEWte9rVvXknBpgY7MjEO7PskuOBtDiIlMvDe1UFlJUGjtv0Hx9p
WutzaYFeAeX0ro41Txp8JawHtiDEmwYZIkGd1p1sE134PDQ5SxS1NjrlZ7uknECmPMjzty8VOjpW
NxaW0gDKYZesogOlx2FOrL9K2ZW4e31/4DtEK7nChUm5yfArDXfWihJqP5p21auSufd8aC43QY6/
d/TMRZR9fWhcftXa2A1u1xD8fzgR9XoD7seg9U7cOwYMrvC845T+BfYOtro8zv+7NT+opnUL3Gnl
viX4WnRWwhL5jjSLADEghM2BsysnedQnT26WItkOTLkP+z2HmAxbTB9AlooJicVxpee/lLvSMqpL
gwNVDVqww/v8jP8bIbaHKrnKDZS3qetqgshpGze0aMmNVN+Mu6q6oC76pLoITxLzDHwcYrfOfDAj
BTDLli8BNPldD0olmaCFgFW8NIcB6T04o10ZVdwnoTlghjHOhNvspu4qXeCLiCkfCzos/lATp78B
2tI5NtnkjPxYy7znLKJFdG8Mo4t5WLDDk03DAqltpN2AbZ23uIyHyiGle6W3f+RZ9OLb1JQiQLPa
cWtUT1mqHTsRuHnJupWy3RgNAHtukpqzZjWcFXBIH3FQpiOuCGDFd3/zisDKST4zbuI1YTJmWrNW
RGQnM5g+bIVR9/HQc2y+ZMhNkjRIQBRqPS23UG7q79V087H1tvs+o3+MxcoHRWAt3hT4zb3RcWa2
1sQw9euN1y9EjZ/Xq43yhloQ+mrOrV1heUC2gpedVn5UnFrCs5+ka1oGIUXyaE+w3S0QO/2QG0x5
SOiJK0mZ8lOzGuaFzfFipCWM2jXvcwCuCKVahbwPUFC+M4wGmSTCXh6Mg4APIPQD5svWCSJYW2Ge
Fe4Np91/CZoRR2X2pPx1pfzoOS96Ka16JO+EbKryMdAnBwX0OgDkEU5YfWg4ZCEUqQ0TqSyHOAxT
67Hp09AU+fQwF2rpSZr+ouQRUkX9rHjwHzXiiLaOzOYsYNme0xEdTxTEtFKtYVK6TvID+E8oYQTw
t6Is7jlSu4bRGbTqjGiF4UbXxVjLYLMx0T+Pmn2e2ny17Ie94G62OWj0/7zRJGBVYZe7/aJ1tK/A
ts7c/Ft7baVi0Y2NHujcEo/Jwh1e/7XGDF9U0kxwurR7hWpQeiZbtqGaGkpmoFBPfFs+DmL0cnSJ
D3rvEDPcFvgFz9piGhm7UM+6nJSsheI6jFhdQes3AjO8MLScO2sKEIZWVdL08dH91Fpe3o9BER5A
x3BYcJfzFQ67tIlOZPG56Stqvx/aZhQNRZjdufTFmsLfwGRwxXi6uyfbi1X4MbRZFlLiEwfudbhg
Hzp1Y1dtmt51fNxggHWG+zV1bRaKHYSrQN6ZW0E6TjSnL9dPjeW6SpPSQhF6Kb3JQAQy2T0fhdKP
36Zqnmy1Tiv2qnbZOYY6jOIhza4NRMA4g3aVHu4J9gd6NLlyowkqfy7Gcjw2beCq8MOCcsFDpA/p
J7r8wfdEvJv2uJae0/sSYU0jR8MZiz2Acsr4EDxuJ2BpCg1M563xY5cq9KJFRB9mV898rvm+W9JA
mBt3UPl+a6io6jruedrjSt9u1C7ZvWQ4ecRYOZqt5V15QgTYWXJ8+aD0eDihT8qTNpv6cmAegOXi
J2PVmAwxl+UgepWlkY57Qn50naRI8GyKel8OKKxBIZoCDRKlH5K4w9uelZhmk4G7/KHy/c3zH1G8
TMVLDZRSWAEZenabpOPv2VVx2uM3xq7IOkig0/u+wSJ62rY4tDSLnhMG5vA3IcuNHv0NpemK+vPU
HDuEJHhPgGSBuuJ1NP3HLhS/1kNuO4T6LrWb+fG30zzDNTOkxprKQ4oe4Zmcb8H7DUSJF2Ni1u+k
8kzM53AhPjvNV4zBVC66IFOq3qu3a5lNj5ldfybiVGa7i/Kv4XQ7wpjMrPeiwV/Eez9s/+T3QLZT
w64FhO6n9pgeX3BvpgV+J9r7mnT+71ioH/VQLonXXSBvjCJzCVtoyxcfLjIHxRwZfVoSJYSW+aU8
skZdFPIwFPnS2Th4xUJmunrD74UiHXEkuVFUEeXa+MMoDFmE72uZLXj1FzHCMmSODDIlUz7lrUia
7Mer4XiSFjneKlcXBXHZLXCHOiLBSYKeZKgK86+P0WNWfF9jhZdfwy09DkfjWaUNS+G+qnV73qy4
i1/DQSW8I763KKNCSVXGfyLlQxqXuegGMU3WbXIPQ2sAkLZJwd5A42wktONsN7K7BNsl8HWGaUCb
+Jno/KMYPv4L6kQLUCuWQ6+Qbq38X0npXLuhByvJceIzJUbQf1wEKhbnSaPzhV+CUPiXYru2dJeQ
Dwxgq6zthbqjlJ3GJgNy2/H4j2BstB2Xg/c7BHDvJZsIvbgQyrOe55kA13ZPZPh9ByYIl9StkNtd
lb5iO7ANt5Yo5H3bsRTD+V/JY+RYXlDDKlF/MYbfP5ig5uZrN3koFSBvFg/DePJo7Ke6NOa2qVPS
fBAfWRGgnqJ6wJZpleLA++15JiYiFWT3b+LjuuLSfkRmIWBsAgO+S7kyntUvmFi39u70nLA/ozGR
fXJAWLJS1qreBEZqa0bIsEUKZNx1GJYPP95I8e/YLL2TVkkfAPK4oC6AopbUcm7CvZFv0cLuqSi0
83FP3zzV0C2w5x8nMNWXEN4+M3SuQK36uySNxpUWpyUCSucEnGXXGb8evbe6ootThchWIwiV+uPB
JdLLRDyR4WC53VaSOA9hZUfHF+t6EDn1uGJqrH15O5VZsqWfvCTWTYp52z8ooPGSjF7A4oNZY1Is
KDkxClB16AZgVnY0mSuE7ffcoKJ/Ym42rAghLX0PmvnqNsSu9bHTc6cwhz+G2g2FjIws9fB42dEx
P+eaOSIP7CEynhFFCt7r3mznw34m3QfwsR6rwnhZzJoTDXuPt4IeOv41N3r9sT+DhYPhQ+gqxwf5
ClMM0YyLOucVLIgvTfaCVBmK7LnPHwUOzrilviwMIdaIfrcXcCAsQsc4+J+Gn7X8wlEkDjggqDaP
GvtrKplkBi5xTtuslxoWBBnysG6mMf+iVVOM7y32psQby3gZe4UzaqJXH25+SdgKwGo2dxj40YW1
F4Y8K0B1MXhV1COY1FygFHKzOkz2HbK6iAzWBrQyVCzD6dJyR6Vm6Y5ruKtmaRS+UkMgHEtjIUZM
vdKfZ+ZDIpYxz691UNPsPXmzL1TZP60cxIPi1PI40VVJK11l6EYbmY9CtY7EUZbw15/KhvsW2C0k
6hqEikbSGQ9UGhRHepRwENX9QWSzSdEr+GUou1whm0Ud1JMuBivofydrkWpwpLE9Mcxips+gh65P
OXRv1GlX2kPqeyJlOklx4B8YXCxKXpPDrQLyEbJZt8t0lAMwBQy2cLqkmvumqjHCNaAaxxGd43Zj
JG2sSGCTyGo8JS64BkQSxikcboCzK54Fk6fbzzJOe9Vh5xU4JPctFGFp/PWzN+LmpM5Q9Hq0xT7o
a416WP4Jhk1zTSlAZfzH1fiYrmoWKYllPEJyBiMm6TXFuNm3tkWI1HoRSQJtT1W2lsokOhkbjl7E
CaGuj0nNcBlCMQ7tmaaWiczbKWcKkzVnL0MX/JzNFt1vXF6a4X6NJ70U2WbkgI9TItKPn6uX3DW2
mHqVnHgmoERy2ylqogkgbwAcLwphIipSMsXqv4jR6M/3E32ECp/vtkr751EMNLJasfzks2Mk/0Xy
FjTgJHwmtC74jQ9gbouj0CXtJFbbnYmHn5FVu7kv9zGGSCb+FgROfXHQE+ayXGqGyEOV3uOYawb6
NcJRokWc02VqQ5n7X/KJ2a5FzSuFdXBNQNjShRdAQ2pM5a1ltuDu88OHMk06SyYTffKrAGAM4pDK
wG90G5gYqqH4GHDZQgU1QCPIqZ/8unZ3azemGzzj/WOaoqReB0sTMd0S7CBJ8mZe+s+onNMd0hMk
pDd7M1xaqHc01pufKhi7gKVpmL2ALu6WEKbtbUdPiDurPJ2HOMC1fqAjJyid1dfRMytRC7xHfHsz
tUbT2F7FtS/wLVS5L9sqoh4zrVdk3uvKZNu5PLtHZkG9rqewXZt/w6/ulPQ6zbvlSYJkKD3DAY+b
KShtN7zNQNj7RiSysjSsp0wJR/SX3hOGH9zL1OHGB5/naxyFMa+rNS4xyttki58YS5K/nAL1+gco
p8DR5ed7BVqbD1ynwHdTW7ZBLLGtWG5nsK7jU+EZUf/inrGdZMJkQ8qa+qSZJDag20FqJDKe11kO
yTDolzeK1wfn2175KSzlFosfP4nqlbdieaLiEmuyy5Tap+lzSkv9qV9SsFUukRituWxIg3ymWOC/
vhpfMbfP4YPzDjLij3/s0ICt3N2aaBhfbDzFg10JTuOu8sd4Nxj+siDvFyDwBczXurWh6q0OIVBh
bR8LevjReXQTot3D3Z473JBay1Dn6kr+WF9llwMbxHObu0xwyuldc6kA3hrtZd34m3jOIvtMkEWM
Od4I2u7cXyRPW7nX+E9Lywn9I25M8WKMP5PXpdr5/UamgMDjhSJUD59HM7TRHU+WX0Prx2YiiCZ3
zJuxSDXrGl1pFRbZpWcOXYUUalmvZWJ7cVlLMuHFgOUVaSR/tnXxsw/PhLczF0wxB6lVDLrTEm38
874Ak0KUegoQIZXMWuFcpx4ssIOU+LXtqJID5K9N4X21Chbx2/oSHST+BxzaAE7KfTsPYZzG7x5r
58+BA64kaNCT2k+E6Dblj+UQHIdT3B7l0M7jGbk9o+ddteNEQdMkk+0JRNlvHaQ1eoiiPLiA3qSH
hrazu8wTg9fmmpMdT4IkCkWJsY6osjEP4P3R3Wzw33KIBN034AQIx7Lnk3TP0dLSvY9LkG83Cmun
nbg6IXhHu9KHEA/NItVbmYORGCFy0PcVaoD2UMj5/t17He8bPAoBd5Bs6Q8Bnk4tGuHNI4VTjj3y
/tBTbYXMhWEwJdzmV7J2ho9TX6mhUZuKGKoYAfXWlF7uEtvtgy8wk0AtdOWnxz8PKs6y14dCIdMr
iYSQ2eVscqDpKrBP/EVIrdPoEPHUraBlYyFN8Wl/C1gCDVc5WdQIH4h48S38zmBnQeaSB2pLGBTU
5VbGRTcN1nSh56EwJK4vuP7XW1oSNFIt19a4HulsN/+3Sg4g9U2AEuW8H4HSRiJEvf7SgBqcHjvb
elofICWjn9AzmuogvFdPZ5v7jaWe9UXkkCpvkDhH9wqPcl6Gg/AeKjRtD3OxFA8WM8ArpBEd5X6o
+HvezOBRdeb4QTh/cnDL24LitBLk1F2tw37a6p0blgURmtfbgAKm4HX0Ugl6GZH9CQlKGkY7szwt
MtzO7Pt+tkIZoLbmhOQeDbTBZMWxuQQN/r2PoYx4aNPyOjC1JXJCfO3J9xH++xM0Y2aSp39s3EFS
3ma7ENu67eS2KEjavpMDbYsi/MR2PrayWNOG2PBzVdtevvBV/og4chmf5BmYmlQlF/w3OTRU9AO5
iVtvANEaxflnvwwGKRNYuiFZHcgG6IfKxuMbfqEDuLfCGynVWNs2KRJgHoM/R8Olxvwm+YnZm160
EV/NiF28xlrC96aqcz4iaJ6Xrfu0XEzF+NLRlOOltFyrl/gNquzIo3lbIbztJWyZ/K3BRuC4JKwN
LF21gCieebE5q1VjowIWAEikSV5fs0Va03RNKZ+9oFn+iVMKng6A6ukq4Eut5MiYdDHufXcCDp4X
hWfLTtsBqhX36jVLdRsmfvDheJI/7HeyOlHuAjBu5UC3pcRjZKDO6jNAZ3FGFClYrGrA2yx0sNL9
b62k5jU7yFFQenV5H7ajOyGN1bVLapalAsbGGDc8MDxCX9On/x7WtPiHK3nIJzD1kSGRoX4v+aLV
aAsNFRJolJB9JlLa6viZujlRS/dVz7AB8ogdPGxG3yvf4vPGtEMtYYL6g/0p38R6tKiPqnnCWK8o
awLvBxLLXCF/J1g9n1WDSuVjOnYXA2t3I4xLNb9wgum2zNLnJdjgWb9Foena9WzfoNpJHbb/4uPR
wZbxuFZ6rCKye9zoYCVBrkho3QrOt88KhqBqxtNuvGPVhSIWxpeMmvchQNpbM//ZFPImbZcEpIlZ
YoVddJh3c5hK1COzHhmTBIn24y9XYMGgwZ8JpxZwrvfK0MgHK1RN2JXgoXAAl3EFHRLpjoIFElLI
Q78S70kHqkQnaVPEQgg/Y1wPhQjtya+5qrsE9g0eKkBHfTfp+aEu2fEtfVk2WN8gqMP/6ghORmmk
HokFEycKX7+pOOnLcx8vUmZC9aj523jS4Y9lgYqtuuP8z6pacp97X8guxn3yJhlklVLgnAURyvRf
GbAuP/VemPMSZdTMdy/gyqG5nyOK+TqoHchb9vd2+iNLstqqWVBhnHYgmyvMwKqb5UmBjv6TbYpG
2+5of7Vr+4ykiI1KCMKhUb1UwpTVAsUna0Ur9qvdTWwpGe+oHII9+5STfT3Cj5LOG8xYkcRvqcAK
j7axwxkkY9YnAp3EGXuCmMOY8zGkT4AucCvTK8o1MMeV8G/dbJKpTYAV/BoyjOF0CDV1DqbqvGJ5
5RcH85qk41o6/5NKM3X8mjZbhszXj51nw0Jih3swfbNKgV7QsdIQDgz7SkSTra9jMug8xsDv4MWb
vtBYDfzwgQNTyTNbDZl52KfvxuMBrOfc2Y3C+fuueKeeEjQjR3Fbd1GZMDCiraY26vUNELsmgDtQ
kFzDtYLrlbZtlP6H4Dk6ZqKVW6SQ4xqkELgj+SppPyiGx6rRXEVDrhlmOW1w70iduRsG/ha+TRwY
uZjqGFl8mZwAIPXQ5dslKCOto6At8xfjNkAuucmeSbq4myk3Wp7KisWSGC65amKgj8yiFshKGMCt
1y3Bc/N5/5NdvI8BbV4jEdGw0gbSSuW6YfvZgxw8LBnOzeWo+3Zs5+EvnS5yDb0eqqlFgKX61Ecp
oQ/TIOmk6ApR5PGkZZhuklAnB3s83qvh1idNld54PJRR6EjOyCpFe3Xy8++O2mH/ChWlmWMrzAz2
7YQsoNWWgymIcwluErhWXIpXDKvbHrYKu/ePie3U8HNH8UfId6p6IFSSLJXC0pe4NRRzFZoRhBCO
YMqYEAeiPIaQRhSB3+naAPiujGku+ygduo2auS8SFi8XCb0xlYF6hnQ0wj7wYiTu7bvQmXaHSgzS
pRX7WjQwtFik6gi+liPcZS+5YjacmyBP8ZAfAu4ZVgqFxdkg98LrTl5uissgPCoKDjH7skFjc9yw
JKHSYegFwKuhBzh0Lt1xByfuJBhDEWijdw52sLCS9cRTyevOdargCkpc4uIWeqs4rgHzN4BYr5+N
tsSuYlcDzAfWetiNiWsXFbSLLqig4l6ilwSDf7VfPcss+XfuFxuaR0XhLX/cKe4dskS53skhnYAQ
+8qyvjwKodE5mq11lFFbrQ99x9mzq+hne1r7Che3Wi6apm55ZlNmode8IC2bQvSEpw6YSkChNUgI
xo7OwJLLplAgDSE+J3PhB+0RIQFz9ZzuYtmPJg7/whAJnjhm/BpF+UOaiC4J01f0ym3+6uQ1is1Q
Adiirn4n8lHkIkDG/P1ZrSeq4gapa6Kn4VTUD80rXam2MR7gl9EbzeOa4kILyongleJjOLA2jgSv
1hSyv2TXNRK3YfOrwVsu7lsLzbm8MmBCRigORdA4JfwpAPaDWwHqVUW09XJLWzBtrun9CaezMONZ
vBg6WEVSU2t6QZXH8lLQ3xGw74F2pmAdU6R0Qbde4tkSdveccd7KlKOdX2Yo/Ql8LLUw2UaI+P9C
XAtVi2AVxFEH4zo0PEhGwM4tL74EZbn1Kt+atf0YB5t/X+7vzHu9nj+3vkX37Efp21pfkRb4ZS3P
KR2Up9NBYVARx9xDXvDLzucs+n8eHFHn4fesSPz3WP1V++O8Uuo+DJV+XoiAIf0AkMKvNsiiRYAE
EyB85uQEbduoAlbG+K8KC46qFqdj6KtjtejYFqYRmLpwN8uv/x0Da7SKMvk6YOO29EN/k6DUPdrN
jSzcG26bpGFNC3EVSmBSrEVce4/PEXy9jol5e0FDfD+ZL6xmOKT2EdX8RwsaB5I1CUUJtGgk3Z3L
x4PqODT0oBIvW1Z2bf/rlQARLESa/MSWNNme36RJVZHWxgT4dXw3wV+m1ZucXv+wsoElfTMMyzOH
bXzRO3puDuMY2X5zSjahoi9aZiCht7yqrZ1f1Vjh+S9Ydxc6WOXrhhFKerbkH89LsdhZDSjsTTY9
hy92/6Oz2WgHrR+TSfa6oD8QZD0eZYiuIV7xOE0NqNdV8i/nawwkk1Nbtr6+sz+FKW1FgXAXYjJK
GuDAjU2RjepGAewOLNQu8N7eXZPHWn/+6wv5ucqVRR1ukLATqps03LkntE08Zxa3dy5Vf8u0d9Q7
y5QddsYNHVV55tQlLaDny6q3jjw13BwuMt977n3izyf2AjA5ricQl1TIIMms6Z/GSeDWotZZU9XB
/CvpnfnORPGrxEKR26XthNsutig8BEl7ykaJ9Cx7N+HB1IrlngFXPhsR8SW+eMD5Bd1YEaCVdPL0
v9NRA6+n8TZ2xSKInLTHDDC1aHwLHDPUHzKCa4ydrh99xtxFXF0V5yE/DxpJrlkT0d7w+9X15jDf
Jf8dABLOszXL2UXb9T4trI1PJ1BevqE8zgqFJDwYFV8Y5+wJZ+WoN2eMFyjuXuC877QeH7GYexnO
rXx9p8INiljTkRS6aw/FLr3rWotPTWw8x6cSRqGWBAX520zsq0lsf3Kdwgx3AR7DPYtys0kS5985
Rg/vmlDrx7P+fjAcARO2Yw5EiASgu3xEBhgT/67z5SVARn7VgeiSszsPb4SZQpTKJaSldyjlGIoV
BDQZGKo6iR8v+DvPPkXjsK5lPCfzKxOaexuPs2oipPckU/2gWnhdswl24Jb95uouWulWUOBl/e3s
Adeum6RMdSezDlovIwBZYXHSSYALE0XEq4qYUItLFcj7qMoFQVq4Er34QA96ahfxHOTO5uUX0RU7
TRBOa+pFx/kaXJDVxdgk2XFDSTq53uMyUGJemE3Cura3zmiaDy6Qa/VBlmp9H/kH92xLU44ZaE2/
VuFgP1SpYnt82qX7HXil5ycCGgytwdiMoHNsGZG+5Ocml/salLcgK3+zsKyeZGv30N9BTDMWXjOe
B9mazXnpnt6PVfEH/DKZcN1SOCN35X25udQkak/c6UvOXnd7BrgBVlqn9CyHQ7uKCSA+d/KDYPh8
cahAWbIMfWEWso0xVJaG7JB4j8zgCezhphC9z8kwx1+rD9GM5KCuWk35u89DWOVejDdo61FtwuhR
V+RGuK+xokSgbcX4zynoKxhg6YqqioYWNplCPvAVzgLyQQ1kiwuPc+i9Ui/g9k7vq32tGqCsXqmR
UVQC2hbHuWpkToDoo/HPSURhaWutFG9jdla253xlr08vfvdGRCtuWWdlXgeqGGTKzQD6Dgzy1mKd
16xACRfhFa3MNx8qwfp8iIfl8k4X47J9mAUW5X6tYV4UdIKeH3MKWvPhBf3AP0KXOgNlcdzlpfKn
9LfcWV/+Q/LWIHHH8HbRdODB1KS4wvGE5yLNz+KX7UZPR2jssiQhL6wJiywAEIs2Jug0XuhTsbhe
82y3uVtLVEVRPuPqIyqcohoop2sQzXuN69rrd2fXp1Co17lbPz0jy/SZZrKNNB0aupZ0GN/0NFNd
kZbddMfQbcAlf42sbOXr/zQXdYivbYDu89oT/FMiqJesHoOz2WmZIcRf1Oir+tGlw19PokyPdG5P
5redN7WvXxBZF2jy+vc6qvQLCiqtkNJhxD5Tfr7IJiaLov3KhIhN/fC9zctqjWlE7pmPsrHzRHpw
rmaTTrRv8aA5d4REsn6ExC6HnzJ4MyjJ23SBWu06zHw5i6ma/jd9KqSdNUI89C9nCiNRs0VVmBS8
ms0sjg6LTSyg2Aylxg+b+CNJOJMZ61AY13GoAYbA5+j8q4GLv4VKtzqzSBEO0XbVvHaHiYTEKxwM
EZOOmWCAG3bZ8+aDaDWq1PEFdBGmNdPQawFqymR1M59v9qdgHdEKiIZmXR8x/zEqky4y6fzvM2Nx
WdWSA5DuuxfXurrDNc4ltrpizEtr3YYwrLTojSBgIsNd+8wvvd0n/mcroBOtZfIxumA3dOkwMWia
Eo6AZK+XnV2P6iq1UWhElYcsMiMV4GmL1baYlnaW44hY1LSOKp47uIJoWxwGi8lmNrVYVjJt4ixM
aCE8nEgyj0jz3dRtFqYjrowewCvctbJzFZN5aK6m9V3C4qMAy4N1NZXngrrSdU32LueI8Nyurdr+
J76vD47oJoFAYEvlZq1+qoGwwd+IQP1GFGkCKke6Mfhqp07I/yZ3djrKyFT1uQjvkhL3mW39Tuy7
Hd13EE0hGZ+vqZFBqkeL/N7Gl/RnTZL6ZODxtOtmZnMOtAHFwsrRM8I/5JPjQKNMbQPKDyKC2w3v
2wWEV6+w3P9skvy1UWE9TyKUszkYcZ6rYGdxie3HnfnP/IInM9XNDfW3P2//aqRD/Vz0TfPazJU4
FkDSN7kQ2USwT4r2XoTOmn5v+7Rm5FSXpTuCnK465sxgYc0YCUU0It+CGU4RhRJSbjde93mu9nQk
o6gaCpfdVFaAvxPDThzD+My4QXIavmrJMnm4zSeoFpeQfv9r5UJODkaK9mp402ySZobbDBrpe6kp
XZ8y/Y3a7+vR5VrcFjbS+c5C+MuPQcclKdFi+wrZThLuYjcsktWIN+RRPQY83WkMFmg4dQe5Dgj7
v7msBNa0hxQqMs46GVvk0qWFVcWMdqfeq3LcnZepsWMA+Soyv3eHtOQ80+TyhIEhGmA8cYcPCszC
8WsLxBggsyBsqm92BXJbFEZMP496EdRCZfbIN+IxFKHq2vHFWh+g3ChHqUntZ5xqTKn3cbMGZreS
IGZNwJWs/AXlH+NTUz/VvHUQbT0Sw3HpL+9uDNC6Yr0Rm6Ks+I1pSXXNYTMJJTdf1mSlaje1WpVi
t2h+4oH3cVxHw9Cyf30Oqqtzc76AuSWMUmw6fuvaEybeKK5d1QIlmqQtmGhkNEyM3hnJRa3YTSFh
iYRiT2AO0yqaWHqTIQ4omUaHs26gQbfa255tJWnJLGcrzJXdo8+k9nfVOeI2BjcUsO5p9aG5AZzH
TMNOG1Z8ZakkbjQ8hDLLgsWnDHw5LeLaiXf6XsiI7FRi5ju6RedxLQZEuwVCWsA08m7iI7X7uwwP
k+JqfG9tXc+90PYt+LsOwIzwJkz89bCOwLxwb4JbwYDkBelxBBwa3S6naXjU7k34mX26O3TKLX7o
NeQjmPumL8saRdt+XNIEOSWSOk4T8/ecW+J8fT6CTp6Tcr9xw3UPTCjaSk2zsdnmVLnO3IEc/OQX
xII+z5OBuCTKQ9lz2UNOcJVo+ZFDoNsiEL+9DNF4n7Ypxp1npj6/NAspf+TB/5JXXIJn02v2KCvr
2vMkD3Ny22Vtn/l71MkH43O45oZXAg0LHdHP8auxUH9KfJtv026785zgFYniK2RMmX4K7lz5AinT
fAPWRr/uzg7tPgSSEaAGWTHy4ryVkV9aiuZvEOm1g69RXCNAgn8fGehE29wNCAGNiip/Ukz8ljOL
AKuSO/5otuEWaQlg3ZU/23IJGfHmLbeX5p9/n8qBGchwxMu7BGWIMyqjkXvV5RbiLU6eIoXzLRdk
pgchD4Xg7Z23VRLjRnujrySkAZ2eWCKyJoqty8aIoR/f22tjltuhY1hLHueS+hTtmIIJQU9vvW3O
7RSE7gX+FF5mgk9VYAbXjE4/Kw1tkQ9YxPtNG7vL+UEFtglzlUovGJRmUhrvHqmkJKKD6WyHMXtM
Din9h0B9Vy4ykmhEkG3vKHipeBy1fziqcdmXCo997SDnPCD1VG2pD5tBa/wMfMFAgeKJEcm4Hh6P
i4xBqWppC06kBh2n2SwumLsFR8JLcqWRdNtWebXxDTEUqUcBmYq959jgQWe/CqgibUOQdTBgtxCF
XniNVI+infZsZ3k2e3KtPTD+r83ePY8iky8CH6rfZ7sXVGq8mV3T8NTg4CRN+9sdksNRV8PUR2eE
hQ1BJux6WjX2mXnVlq8WLtW0eT0XunPic4M/gXIF3IgOl7ASYa+PNEs2QwUrA5YJfFWkZJyBcVzT
REfr0GMZYfjF/JYtsRcZjv5SxSqakBEhTP5cMxfveNz2pJSRGQKb7Jvw3hgF/VtVuTMsmXSh5cpk
RTL3oFccZxPihfY2e8NaEWfzJKNA5M2M8pcCFSOfj45tEJ6zWpVvd+jGfR3qf4Ri4vfg64lJRWa/
pyvuVtqOR4aqE03HLCYzZqlKCUeEX7MsPwOvyB8Sgx6GtBQXGosePWdqThT/AKf+J/7Qo9ZA+oH+
tPN+Cz/qOFyVcPdFim+qLktoqPAuk3ypRvTKDojL5hF7DPY1nrYxEtvoHN3Pe6r+yfKQHF4G/v2h
YxOuy7uLuLiWoQPJ772rdx9HjBTtfzJIL3LGzF9pIxkR5Eq+Zwo9VHtZCKO/cM9OwQxL+gSZ9406
oNnsgVbMv4s7NAlL1LsRdE8tup2Ej32fqLrL5QJo7PfTSoRyfvR/UGFCd99y7lPCD/5fALyvLoDy
8o7kDdVHv7uRmjuKTJruTR9tcWgIOoNhSWa3rdK3nQCgoapHAsIv+PM6vjG2JXROikKJFgq5HVSj
GfTkTay733xEAwd0lefUKd+HU7R7pWiyEXlX1yERstOYBcfH/qGgeXFALaIjm0GI+0DLfjLfoeOl
GHi2Jyhof56+4YZ3FxzjQy891ABHNJtuSX30xR2NQDm7rMdElacA5OkRVhqlHQ4uvcLTpy74OB41
HW0eEMjPW2pDr8J1G3rT9MgUgs2Y3drMV55cd31K70IXbK/0QO0OoDXzqTz4/ooy8BJJ7wtzhhgm
4eM4v8tMQ+6HjtSxcBHMu1UDIz0inXqf7XvMYuFR4WwiDzD9c4UqX0IZiAfBLXh4dXpxkI1bpwx3
PpWGoDSzbp5Wn47k2isbuMjuG0cUS/IGK+aLmF8ZnFEA4UCnJTnxxXZLbaSU7u/IhAJiLr+s7Jsv
iyVoWzsJHtlZJGmdcaQccliZaslY1LeEcyOiThVE/NwzBTQttkkH20QNmedidm1TxGmvHgoMZcXb
LZuMjalV4c6vfV0lA7fn59CvQ/051d9fYkMx/NGYOCXBuF2lgiXR1/DpdaxqTm0GlXxxpytntlT6
GKBmSvqPyUnf8e7v5N7auVta8R6VRZ4EAsp6m8f4+HzeaKB8EGlXh2PDpegOm6b807D+WtaUv7so
64hs23Be51qA/gb9whpUFptJg/nOz2nolCtwlHy9AUf8TV6ZqGa11qMXSH8odMDU/E6+YoZoTSCM
YNNNcKSq8/bJu8JBqSaIaLlgdZj6OX0xPFNsnTYjAZ2VzBz4t+wclxC1t7MVpLe7xS5PqwehhSoQ
K/dklZZKIlVbVu1yp33iDpHmda6p/4F0TFSoyTd6Qk2hyYgUD13fbL27rDq4U+SGubx1FwtIR4g1
2WeKnBF1EDmOsnevsC4QU8atjqoQCNitFsbf47IoMyvT9pQ/KABc9+WizRBbGHW/WrLA1vpgsgCo
apYBW1vwWG8OAnbUaqoyL1MwcktuupSm1YvoaDJ6+wLpUHeRKkiz5xYSbTn9UHavLk+u8PiT2gPi
KEep2rkgMZVvII9c0ofN8x3O75nQD4Ge7Z9rMoSA/tesq2lY4a72BuvLuB8Cz7oYI7ea3Uv2liXV
JLm9SSQVW6MZf4iixO7MakeCz0Q2hI7d499E+dGEpt0yJMp/IvBlPmjP4qspUPS+56R9o1kJ5/ir
gLEXkhGQ6Y0TQ1X7Gh1/TONImlFEb0WxpZaJdyyYf12Zoizg8qf/Rl3xN1N08/qvrBHGAECJrIZI
NcpKfb1cbgLWgSMLUtP+8rNUv0QPcO9h1R5iV+4IYivwlsfFxTyB6Mp3WfK8t+3Hn2bXHVaKvzzh
8kODnxEDKghksmxJXmccIQgkkQlNMZbHcVI3f3TCBb9ymwHx62grlig0Y43AiofDXeLSNcqGpZtA
vkAUx73Uc/Z72RsO29DeoNSfGss1Yw3ugAo8kmghDSuy3h48MrJNSdD3mf9bTDiPc1SaIRs7Zg3+
SEObuhRZ9uIwgEE21LJpltlGZ1F7itOQU+Y5oQPdLiPR/0Km0DWMCTl3yq1muz86/8eG4ReKnhoX
bCcEkMImK7Ys9NS58qXqtxdcGU94yU+lmvqGyGx9GSTyTBuEC//hywyBLOlwLULOyXAZkE6XH0+5
r2GcGpilbcv74GL+VWetE8jbPZfszStyNm0sAwBD54BMeJlOBfzEDZX19etjqIo97yAS07sOgGeH
r1kADzbR/P8Kug1jJMQzOVa0zsfhiiU/WIm0ClzfHDnpv1B/Fk/D+X67ZPmFnnLHxtlXD0k9clin
DOovXHnLj8KesB56TCWDEe/YKRo3HOYCWEtK/dewv+hvpFtOjleZakOLl58zh0K4EhVBu1dt6x3a
1fAM4G6HbtyM1K3sULGwA9WTqdtGG70TbIqgucI6o3zLBYXKntPGYPJbARn+ervJVANI0UojDWkj
bpuL4GSUEjviknjN7Y+Y1Y7cXA1xVOntxiRgST3MkQaC+qxYODjuY2T+j27/O6Ag8n8MGrPfy15V
ZVpu/8VFRBrfIMrpE/LvwmPipgXXfPeJsIcdWb3rGLNx15qKY6zSSwAhc/STMUpikXFYeYSjGhxh
Wox7D/PNNiEjxc/aVBXp5kWn5vEXsmi9X6JJrycVQlgXjWoM5DBDxwW09N1e2NFwMNo5aes33+ue
RMnq7Dgk+WQJrwNKF/1km6yMqYRVUhHVNZSjmrMPPClhxqTuq2nyrGajQ7jaw/37wJtFhJnDtzlj
4FfJBJc8kZfzl2xtWLgN9Z8xEaVvlDg+hj+Ox0OYeXKM4QRl5U7O2edIs7Nblp/dwUmjNuJ0rJh2
UWoSAlG+5vfU6C5v/QFPOCzuxR3Q9Cx3RX/Ill7BfM41V7Y24+/xDpE7dIr0vQ5Ocw29kvGi+VbK
rXwbN2FfsJ/EJjH/h9G7fgbs2fjSfUfeDrmyH7SwgA4PQ1t9UbM2geaKuhQ9Fo2XtjpLly/+LUlw
Cevk0LucMuqrd0NoUAVcYGxI3CpU0BU4dZoMHYZQVS/4GzBZirnkBby0sGRe/LEEJv5CtLHE7QyJ
5VVcipAyZn5fAgUIkQFCMacwrlGnLzQ0PcRjVTskklCwYnnRgrZjfOPKHt52Q75PX2fD7oxyPYEZ
c7GQ1qn9HMQSKQVnhJTtH2oj+wTNWlYjr/jt1EK3Yw5C1HbG7wsoGGzsYHx3Ovx/VniQ0JgeXeCT
DFQqEfQjNZIzbTJrDOlWG1TCi4wpqV4xYYnN8dAPpHZj3OJXRSWkxd9lw+gILczkipgHKOwR+D8m
iNtBzxHDVaSgzFOWymZg14rbWqRRTE13FCiZ7mAN5mV47aPZO/mgkBSY0YmTuhsZl3VQ0gKRVju2
I8GnhkZGnJTZQNmEDJfsmW34t82WMxZ5RYrlONpTmDAe1pi0+cMCRsT92kKaTpdlQvqhAnVO9SQA
0JB35ToHtdJehfoFeBnexEYEDNCzyZFx5nv/WbgnIirYetDXuFh4zWsqXL72ObOk6JjXg0/8di7j
SXBevSGH7G2mZDdCjyNG4W20eZShNywjHl5CPTEGCZNNs3DB2joY/FoG+fN6aQyc3wK/IRdGUfda
+PjxBjp/BTOel8YmbfH+/qoEcOuMRM7moxchFp5IMqtlWnjmVhN8YZLYs0ly/g5/Kk27gDQ7+kXD
05MkVtcTdic0st9foAuiOtp42FlVdpDUSOz2hIsBjtgWe789ZydyzxLV96NvjLLjPpk09qA3xfGr
kbeCChCLB3TZKUdhaL86BwAwt9bxpIMMNa+LGOpeG5qEhFv99tzvIzcHP3YeAUQsV7dcGKSRAxYx
FHfWnOfN5ZYOs1TA1lSoAOkoAg9Kwgp4i+370zfHGr8gmszsPme/ulqnvm69ovpnj4qzp4/QpoXw
o0ygM0bti/wwK4qF6xgwB3TnlUI3o/5bUtSYYbyvWFWw7rFSGtZGQ1by2sx4z8cGv9DUXggPIy4T
MWaML1DyWYb2WoOHEEykJ0ThXXbwNXZS7TgxoATDgWZQZyHUybohT9K7oW81rYt+wkhgGSfQ7R+n
prvNCRMHK9zG7np9LIXiK8POHeaAQ0IQOSwKWlB8mquCdMkrFZ7zz+3boPiUtQuYBZZbXskg6FUP
jM/4qy68bz/LQxMDCoBKnnA+qNGcXvIOljR1h8duoDG8CEJMgn4UYoUopBBjL63EFQ3kJLk15S1X
Jp1KeCmHYv/o8Hu1Ud0f0Ol+f5ZpRg1glWdZxYfhki+7byykaq6hOxoj7WyrDjOTuWGl6ydu9PJL
ASXcHrqOml5rnwANCo7IMYFu5ZiWTT1fT1xkVOCsYC5rPcg4XCxV179BTcKxFdFoyuIUvubqSOCQ
Vi/4Kyf1yN0G+F6mSEKqlRJwCbRKStgHAob1ADM8ii+f628UJmc4ktwnzDFOBzenCVQ6MKaEDfFq
HkFMvjIAtpKgsWt4NquI84O4C7iuzXO9iRoMXtiFJtUv/Kl23uMHwSh0JuoJ8QIa4m7Qh848eQbP
vuP/z1r0DFzEnNXHFQjsHYm7pT2QEcTeAjpOhLcmIYvxteQbnoOpOvTFL5tyOqMYgG4jrdmeJVmg
fBsHn8nptBeXFSjBO9tSOPAUpwCQmcK8oeBK7S8kLhYxRPQgGt/of6whJu9Of0FheJcOHlGOvkkl
m9uhIG3QfvN3lwKvCp/vTBqvRnyyrfLhxEBDMSAho5A2JwiQxMVj4LP7ApNESlH5uBHUh7x+TScl
DWzL/Tx0qFhoRd9Hn2s1hMpUKctdnGoMPJPe9A7Uh0/PH69yJJLZi9MtP7FCYptJr694UWko1R5c
BUgpg163nt9BBUMpxFurCyweCFsB9CVwLviJQs+NK+wLyiQ3o11211FLnbK1VKJFPJkB8x2o6bD8
L6MJuSvkDrisUX/jZ7iuZMmyES0JHEdOT10jh47h0NYuO3ah3t92d4SDObQsCYv0GBs1/x9RT/td
G6l0mg5hBAHunaAEodfv/Ou1aNRTHM/puspj8WVN1yX94VIYcI8o3tQfK+Xwk0lfhSSKiZY6gGEt
m5aJ3zgSAdJeBy+2PtzIBUbMGD321IHkpAoxpYxuvm1eFv4WUd4cb7dYWWeqhyH+7U6fMEM4WVQu
dtZ/iGXzLN/9GcHDv0SuX0oMHuYhASjU7ENF1X51CYw28LmTBZI/1nStYjDQcvYT3chvd4+4qXzH
zeux+t4oKtT0Z3OrKcSOblqdiH+3GQ2gpSiOoB0FOC3OJ491LhPV9f2F1Fuf8JbqEUpx1BCqdMOe
YeEzXqWKYz16uGudC0zZsZkCfx1GXpvkuEpENx7Rvq5u08NhGVDTaqjsqORYpQLvtPQKDKaPyFmG
ITnldV9BovyYYLoM3ZugUzB7RIy+qqHJLUIfcUrYgwAnD5xnnVOMndhYpcXJP/KU+vtAqb5ivSBa
NhxNo0YMoDEaYixURE1vvjDFdyppOEmlkNpB+gXStizpE54iS/c6RdFuRSntTucigqywOEaiWWEL
ut7UZu2LembfmhknVev0ksMn9DAIAVSAzfcryWrtrglIWC7gjt2RgE+PTbD8k23QAEYPvS+8412W
g4Q6bI83/kKk2GrR3ZtPIGbS2mGhrVzTr6pTDyL013+lecDcJr/aujyYjDek5BDsIkvaaOb/f1E6
piNT/Vei5XEnFB8alDKPg6LI+DE9urnkRiuxWa5bDczubgLDc8cMXGnQS3wEF4nTHjAWaPprNvB2
nAE7bnPkXMtPd+wYeXYQyda5RK/MQ7mgh3pdgar5N81tsN/sDysyzd7zsT+s0PogS9+Vop1CMuzc
IPcBXwrX6b4UWmK1C+zl2LjxOXqbf1/1Y8o+j22vtEWZhe33sy/itI+jrZ4ckOEvRktkA4AyxcfW
ma30yTqm6O4K0HQqWy/CGfQ7hiqm2c+njHNNHueQ17SrkUMFISXi35KRMeg6jNEVf9hIGjNKzEhL
JM+lA3J8FCm2BqXSEhNCekBgc3WJBR48ZrJ9R+J4IPLMrjklz+0wYEaN/agHUnhAOGFhLk5zq16a
7upqwbgGv81lQnp+rDOVlK/TffO0YE0npV08MsQJyA6Ggp6zYNMghGjnU8kkw0me1hX3/x44+RC9
HxGuENNh4EAaET54QqBoUiaIoJV5/dhu0YyhdC1QUUZmdrbAl7UHYCjcUYEw5QcKuGJE7xNhqwCG
eafYcO/qtDm6VvY9LDa8TKkvtU8NsVmO8EFmrwhq2z0hA5NoL+l8m+ptsw7XV5u98dD4DJuPMwPZ
wfibhTyK8VUPiZmuMAdw7l2uNnkXQcEXTLNs+8ajmzoH/DV0/Qr5lB6TmEnX+Ua/js3+6kZm7CiT
JWMvffAoKfTh5BJoRqQzUiv17aG5FWo6W/aTaM23fC5/YCERGyz+/VDz9W+NiJVrFaS3lAJVafBS
0svlY3dSM2oG+2Ux8DqhoCWzzk9lzEhjacF6tFe1oKZVlv1/kotI5S57wSu11NYApWqe+rY6ndJz
GOHNbmltXO81fjT7wV+iDlYH0h5ojUMER2nMUK5ZOMmPFfnFk+o2a+gLWBjmdxzpFFP8+UNoNjWQ
EwDUNZ9FcDSzsOSA/0tjugAbnSJFyt8emYzfS5GzMfQ6RoFzpECyVA9j6sBhXfXELPwILre9+/8s
auWNm7XNyCDWEk5kPd1oyDholiE2WhuxzwiAjq8WJQnIVOOh34b4hi26h3Ro9M7y63bRqcBH2vZP
riITdUrwNXya6YrQjwCzjtktyTaMfEleurNaYqrBGID804Z5H2bGHZI0Mtu+/UWGzxrKjREA2eGV
1vZiDSiFsCYhdS1OcoQO6JzBf/Y+Gf2rymOTst0ZMjKtxQwEB30pUi/8z1x+sLxldbdOyRaYNh9P
Gk0ZaBQlwBTIWbbNaSAyiMDbZVwZQJCRcxYJ0enPkZtvvmNHX+2G1f/3L8nvmqXETZZ2Wt/2StEp
72iP++Cygj8xvLaepagOnJsBV59cIAbpwk2IFN9Nc/rOnz0M12QmmmY9sUQM7ATQgxXYgu1AqrWu
FgpQ48HLz0bjJRyUoE06zGcoygzl+Uc7g6w7mbMQuWVOxd8utKa8ZrZ64fX+uHS/hG8RqKBaQ3xE
oMTNdBTFx49o2Tg0QzysyjUGreCLvD9etR39eXbw6TrBftp/GpFVRMJ4MpxjTM+umZJwIEwPIwUU
PCvpjad19FKTlXxfIkIwYElYjzzU1AqiAEvz7U1JFQIVm8Tic2dZV8hCeoVrfPwJZhvE/qpibXbN
J2eiHKotMWCSWvOWphFV81k0Jrm2BWF/00LjpTTlOHzb0BJFQPM1J96j9UIvkt9NczDjKgw81SVG
hFF8TPRSe40J1VNIGgQBXEO1bLZrKQJ1rhpMu2r9MPrCoLAFvmWcXH0ZYIB42znekIbKn2dlvXud
20cqRtDKNWwH0uZchdBsU97lzWCbVQxfmVq9bJYPqH2STnJKFY43jP7nXVNZ/4w2/B8Qr9fVtPml
bZHJGR6rN7Wg9i68sN6v+ThEYaMImjx6yP2BnDZ2lFLnuAvHlc5ignbnPssgEN12wMcJXfs7Bsg9
WnLxgAvmLfDft6FW9W2sZJlsZV9jORCqS7mOznxOX4UnREHzSk+RSTSYFY3Ygu/nx6cBmBgHgIvP
f3Vic6dlEzyR2zeNru7DmiDKrjnUrud5v461rBmKekylnRexqObmXrASv848LtSX0hw0U37gVdHA
2Fd/HSvCSMGoNWiLGXNlWxwriYns+JVKeRdDg4R+uNA9Foq46wwRCynQvN50UXmVaZdyVYDy6gWP
zXBdfvZjxH1Oy2xubshlJ5+5B+21K+pSmR+jcAjpwLDBRBSl9FmdOl/tTJjTFkG7HCV4CY0KOVe6
TrRpsw/h1f5P0zSbC5HVDw5yn1GDLrFKZtKtdFdHjC1eAdxwTJdNFW+3L7Pr8Flvhn8JHNWjbsQ1
PcnKpP3gldJvBv2woQH2DZfOQnyiPLXFS53hRpbHOy8A2V3ILwhfZw+D+vaolGDEn0ki8kRfFMrp
S7EUciIdYif+XXisEhDZBO2yhOi+SYC+orSmDcitoAMWptk4J7MipzUPVvRixMT+GoCyYLNFhieE
TjKkW5ZzZWvy7YRoxUU0by9HFF+wifKKFaDAiBrfAzufkCsoHGtzi7hH32FkRH0DrumLZTDYLxuI
14aKcWgyzL696wgWuMb2tRLpe31g6j4DstqtRu7LV2jK6wMytgeoxE+bq4xdLX3XSUuC/+Gnt3Gp
lUAGTvuMzNq+f9fU9gOLOl2LSQEsMqhajjpXpSXVRBWWDadLd/D/fY68OiQWLGa0M851GjU3zQRg
6rBlNebM/uhkosBM6esAygq3uNkxyn9UZKoXRn4Os2bJk4nw8XrQWta0xj/s544Hz5zIN/yPofgL
f2/PySVNR6k1yrllSXq1ksUiNefwZlYdnfdZFfbN6lOv1JzhJ1r9vycO/AEbYnqe6lYSG1gsFLOb
aJKE7ojPV1l43+rB+1xM+LuxjgODD0l3KqgVtmO0o9xk1mNPEnCk8Pf8FyATYaXLZFOpgivRzNLq
1UhsT6YQGfxWMFYcBjYw6yhw4xadwkxulT7GLY5hzj9ZnBlqdXyG9aneroO23S1cc/iosZaGKVs4
p7W50bbErXSiFpr18XEFmO9DNgAJ9SnOh53zGiO62hcTbDUjuUT0vKs12Sllu66UVz5hjZdst6WJ
gzk1LnHDejLpu0E5sNpHi+X9LhrUr26eGdzWCDcwJpkCMi+lv+/ZxC4JnbNoXC/coCg+YOhKeehM
EzEe2TgmsKmlSN4v+vdezbTHc0c4akO/m3bwaph3pY/EM8prbNJczDpm2yYOGmgsM04dgvZaza6j
/f4sWwiqwKH/sS0zbJM5FQqlSjYFhCB1BUOyhE8oYhJuZ7eQjX/Xjtni9lfN/Zh3zyYJxbhnJ2HQ
DaKbBoFDA7NRe8V3Zf6ejGKXSia/djbU/JYwXH0hO19yUXokE+1gQ8VodjHkYCnHxjsyiRebrLo8
h+Ka3gSnoVsCmTsf0KW8taNRJVruE3GvvXJ8oTLokXl0Jh4QNVAxhRGpBeDoOUp/6DZZ3QUPlSb2
PexVzvHdmWVHerNdTMYM+C0dQqI/cehlxsDF9Y623VyBeT2wUZxVqWGJpfQ56Ix9x5iB8OyEduvR
qCCgM0wNk9GEnTFYx4ygYb6da731tzlKlWjoCvBYKm3WIRQGZTHPzJTnmGvP7WDRYf2f8a8ERr70
mOdnEQTGzJVPvxUetqtSXSKuGFYdbpRLQiWnT+rJjcl9sAsDdwtjr2GSzC3fbA2WlhQ7FVeToM9H
tsLmJSCzai8nU5tLSpKIqW+E5X0VwDcJzlp39NLkn93X2bDfFSOzoSUP3F10hL0XFxgfokmBxUz8
2kDIRdPhHGoPD4G5JSlGYbkJUHwx/GUigqDjzO+YYXa5uhe+yvPan2biSJW9yD7nNXQ0yNTPdEGq
chWw92k9s2lIkimbf57LqIYr9Z75ILEmt8ehfXoKGlQ07sEs4rAJzUTcTHmteB/IyIhZ1XoLmfe2
HrvPqQJHWi/hU4Eyr0j+56dJFLQ/QTbpDptM6xTl4VGx8b94C0ePEEUlT11f94phgDHovQDQCYjH
1IgAqwh2eGER+nkbi+0YwSs0i4+HxvL/WpbFBOwm37fHh/0utUHq6fL8v0XSBwcLstOb+ZJpg755
ht8LpGFVW+ZbkSs8KeeLA/sKBwzervLpFTnkP9Y6LYSE+AkuldvEIg2cPoteWR1QqBt4WpjS8w+O
g9rN+mk5ra1Jp9xjwxuNK8r3lMJ3tHXPUHXx5F/fJMgd57Lrs3rVWGfeouBTNKfv4CYhRnCpAaP0
dtFSVbS66PmNhYRRGIDACFrI+6JexVmKMCPYIwWHOvy9iz77pECRxcIdlZzwB9TkPJzPMYEmjhvJ
pLiBs5Y2a2JUbUZ0kzEz3/TPFVQOvxh0QIuuOKVQx+3AVaVapRpoWsR676uIze78NnaTZzC4cO3k
F1JtiDJub33OIaEpTMcSxp4gALzt/7gFsQaejq5U/w1FsSvtBFxfrvm3qBUn325kDqgTydCpjMAN
KDQwlYzPGA8dzg+Grp64fYtRi8XfcSa1MMc5lW8VmIDkANUazdh2kYzl7HtyLvI9+WB0JMu2UXbt
w11TcaGTTmmrDtVf9cx+RpaA3Hrcsn968jDS1Tn6b+ggpNDTjHv/fMkxnizLUM2WNWIOWeKWt/Jm
tL3j4kBerUH6rK71Du1swq0QH/crhp3Omoms/gYv44MaqchU6MIKojOclNEOmvDFn4AKKFBv9qka
tXQyEkbHJ/3GROlPp4BgG/gr5SEF38wcGVrcgwvkEQVKOKkIpkdqh4qYLorubGmbTZUSfwJLFiaQ
MBLthyOfuaQwI+Kv+jqn+l/UJjYSyShyxHDCFTCcmLaC/YGdpg2yCiOcS9pd/ut0zVY9C9TDn2Py
nTLxO62OI72zDXMj8XBL4ksp9awhteYMpfo7OzkL6+6nspVh3ngHHqjpOWcrP1OdQ9FlUga5pNZW
4dushT1kboO8/pp1faL2q24Z8hFgUAlOwT3oF8c40ma8/3pOPYDgRbq/eZc3YraeDlzedSvllWuJ
61XHAxFq0nwcvSut4SNFhQq2ZF0x3V/If3ERZ7gw27xVNhhHxxgP/KHOKbd7SsEKb38M+wuUx8tN
A7WQR0ZacRKdhQcgd3Lk0SOHA8GFU5IMzFbWd6JOoKC46BWgvvg0A5G050/vvATLjKG0l2G0+QET
3hf4uQWyru/Vsx8AGxjwgmdgOvK6Nla2/rYj+j79E7ds9faqgK3flTlWZn8J7Ro82N63zjdVxCQQ
PaMudi+ZkvfCwLu7TYVIaAPeA4t3gTY29eZEZbydr31+x5J6PE9UDmE28Watwgee2HGFKjvZzQHi
rbgb2gw2p0GMMEvWnsoQSzTmUJf+AhTUMmjXCrP2nZnKKY5f3TsYSyE2/Pa7czXsdATkmSQq7a2z
mKgc+eLXIkEqd8DK5VRZcGf7szI9o6QO84bJ2m4Rh2BjZ6vW0nFCm17QHN682Qsl+a1rE+RUjuIj
QakHVobliY8TvJhE+RJKG9sV2uSIkZQI1ATVc22gJqsp6UNTYZR6ik1t2z1bf+t6Y+Xgoiz5MnTm
f7WYXjV+aSOXT4yZxVxUDD7sXpTXajKJLcXeY1CTKGb1J/zpMGZpVcFM4MxvY58GWkU77F2UFOQn
reyWbbkjWJdsZ278/Zlfn2g5ytl1Pb6Mt/F9DNU6nMTavg7iqGuih6uvVatm/KeGwdspyhQT5oMR
1MK2zQTKIp+uEGmRUyjxoplJ8I26uMjkWzwXwCW36juD+a613hRxK7bAtEVBOKNFX/bJQqfnzSJJ
I3ZhrikGXm5nekCh1HOVkxZJlGW8TQ6RPf0wzdF0x2kXHvGKamWkRKbWojYgtd+sjX2f8VCh/cy7
LSne3fp77FpboJKJ4uELyqovZiuxMVsO66c20sHUD06eDVvSpFAaWKRRa3GbIBL6TILNaHt0wJAs
5ptuse6h6l7lzrI/gapYylqhnuOYY5k7QsQFxTyWhAJvCBcbmWkf81StfLl5gyuaUvaFpjGOI5N1
cWIsViadS14cL7wAD3BP0m5TPS8UNEQ5J1mBEzve9TBqGuD/NtkUp3O80k7JAuUFaL51Lzcz3Wnd
yIVkBbM2Xev9BrrH3+y3MAa2JRhiUojYgGhcBLid7Ic+wsCJkaX5rWKrPo3UZ0nmo8EAeE9OIqot
PAWrzhw4AlaECOrdGvFTi4JIYD+u6iDxEzo3aeH9jyidTHSJQcqdYolhSZ0XW61pruwd+5cZzbBA
wnKmo2l7ZswKM8gpqRjiuhNpExDDI9w538oAzSnFq6gjCbghFX+aO4phg5yMluAQenv+35ufXCgD
R53jp+rrLgKZqOk1FPqtbyAp1D1Fa/zvSCcAIgZk2DETiCcwTbEkt964fWUjVUiU4k8RRLFGESm3
GmNLTSmDzXhGAIzevh1mUJDI1bi59B62T5FQWg36MZcg6N92UJejWHnEqTT8H8i1u+Up5vomUflO
h9rt/2Z8Z9kRgnAgGMILSIiT2axL09tizUfpSUwaYjIKYBwM0QWXYjgg4EnXMnvEeujXNFP5YJig
pR6OaGz9PdzG5kjMzU5tTd68Wf4+qNyA8VtiKBGlM1cAoFV8M/YQDeGib3267HuU5fh5uGGQkR6G
zM2F/ZxItfALg5cFHo8ZEfFWenNLBmM4Diq9noqInQbvlc2IAQcNFxLvw5Vd/nvEoIYYeTs9yUzQ
XRk43ldWmvJLsUCHwlG68quGinolBL+8Gyb7Z1RLUdglnX5xs4kUR8Mk7GgiJmGRTqkprqM0dr+M
C9tXxA0DvH1ZhPk4zpN3yqaqG193Ftf8Y5h6/oXVQcJA4YkIWXpXpuZsXBPfZoaAu1PT588WBziS
7d3C5vOQA54HJUHRf1h12fmM+tTT2ArkiYr5JISq+Lagen84CRXY/x7VxHqSHbstUkGUmtA47JJZ
/ZB13VTqI2RVztbdER5jqWvRkC3dbdqpSmFTMMiQiRZ/KQwrYvTN9+n7GhcclnrHSHfgFOlgmIVC
1fnR1vr2oqggXjNgGhwEZ5MKZGwFk1mY8VL/O5k+Kp8sOA1uQaNyeZBrmnrtNeR2W1DVwQQV36W1
AhcG2mlnug8aft3lfemVEAICwbSh+sUT/aYPxJYLv8yOZA6zWVkYSdycgmnEdVtw8c5FnOxvhgSm
3LChm+oVnmlhmsdU9jBFzKLC8vyDN8UEoXq3WCRF6OK96EZ0lRf3a6d+PhNt+GeBmLFwoQei0KyU
MNhSUBJvx0OETa4ovb0tY/74puWHyyZcXyuxQZ8TpLCTR4gy1AbtZeAyq+pUakK02c+sq9QT5ICS
r9MT5acNq6h3CmKMwRxLYOD5j0s9Yhw/bC7su61yDjgrx7P4ClmkX6bb0iFMibwCCPU7boRXz52N
xG5QrffguNFS8fQ4nizVINCJ1sCu2mV2JUnwesGCQQM0oQdZzQBgauPMf1xauzCwbUW2FB4lxbxA
70vcD5PRVbKcfa2sb/2zOoC838f1VBuliumNqc60FBT44otk7/t1tzSx7RNSkvAjY/jVG8yOQ0Rq
SlJyI1wW1gMFTNIS6fIkshea1JuPDu/IXDgzy0BUyGHJnnAgvQ9C43jJ5tpt2uPIQf9JjXd6EdqZ
sX9UkCef8aI5k7AlOoBorn0hO8Ulxf2FVgTJv5h/KZ8JwYNx48DYAEXBwyeY6nth8BReMpTWQJLC
TqzfAwV1GavZWrsqPjPgPMIr8v3ofi4K2V8IYbsGIHc7+Oz9TBr5gMFbptsqUbRyzap0vOyPCoqs
hKFUSZ1SEKVE3xgN1kqTuINn7tgPZApeszFfwfOMHrw7k9h7CLEETOouCv7qQstUEigYl1aNSGGo
XOM7GnA7RoOAtckgnzYonkF4ytFYhx8nHfMyunjeAXuDjBvKuzWF5t2hcr9MXfpsbhROkSWXnek4
+apybOf5KbpwnE34uDYRC0XCRWM2FkVWncOohdeUnWkKwwwVptHC36ALfW733wc2Ip5GJxu3WAkY
ZNSHJGgj09Jd4Cdw4+HNtXjkbjDOCevWM4letfZ+2QVLiEkXOi5o8xNAMakFC8xVE5SHBZfVZEwc
jBYLq8CWMqtitVIjsFWuzVAS58DQyZ1W/1e+4C1Ljv0Z6qSQmwwcnHP8sZc/+5YFMdqcwgmWE7GO
Gyxe7YyIU9Tr5M2xzqBGkLrurEiixozm2nYqlQZ3cLZ5Zh4zxBHDtZLOQeoTg4QDNT3mFDrUSt4t
wCfsLO8RfXSIsjEOA3dRHhufFfho28QtTIJWf7SeB8rdTYwWKGf2qBgwabZ8HBL7l5Wdffsleiwe
5CtBcn9H6kuBgDq8ryBe4owPk1Fiw1s6ckPOzfqi6HKF+dCpZnJqDoJ4P0ZS9IXkEH0rxe9ulC+x
/hOxa/Ju8vTCVz3d9EA+rrZ5V1GkxguWxP++6ke3wYtA2bDCCpfv97m+woMECpdgler4VzAfTKyE
5pidNvz5WzZUwyBIl/+Jt06B1HcKNYoI4ffeWF8mYMlCH7KZSc5oNeXqaZZe6K+lzLGCYb+vRLrl
Kc++rNwHHSzdKSsl/b11JcOHS//yQgG34qBk8BRNVs3cMBaqHIzkzf3hQuLggJ4Ctdvwf1wKVkFX
K/Kdu9Ck5fcH8GfAsVnaU5EGoaRHCi/W2h50wijWW+mYJTBdN2lMe6wf3Px6zNlsSrWA3PK0XQCw
knmHlMVFGIkyMWCgXfMihf1hmzmBgO5i9F9WPqSWnWWD2NPZOfhneWiU/2hK1BCi7maokiItYoyL
9g5rlh68/VM7T+8bHWcmMjvywdfeV1f0ijX1FtK7WomdWChKnFfKtrQk+QuAw9NpE9/dh3KiH8Xt
YxYsosNnQuovwSwFHPmXqJ75MbIAZwwZxRS9mtJuraCOKyfGpM3rZ6D+5n8rMjj/XfeT9BkhThSH
266mH/7I7k+TQxYqxlMr8LgIqf4ZOHmHvRDu8v7BO8FLLj3Arl+ts3nmBbAoxR14Z6mUv2Tw2eeu
1lZoA1bEsQVw0h7yuS0QhzezBUkqp1oohLQ+A+IPhU9Ns4eda30brZVFle2FQAL8CyxWQuLblj+7
N6koYtunlugRCH2uV6fBaDcmQNpJrHz2WOy5w7TIMBqqNNjh0JoJ/0PCpNxJgRehYEJqIgCF9K1W
j1Wp0uTZHGdLuLlzbIEH+ShQTK9aScE4D0ZQdhgXgNAy/IUtqgSRX+U6mM6BFOu2wu3+z0eVeg2O
6hQ3qBp4czPIXQI8Udn2oUSVNCVvKPnmkXKDq3TOsk+CJvAksyr2/OGWcDJuuObqUgbq37HqdF8z
CFTIfYsLO7np4pWAuGPCqHgj6Df/vaugvJAssR6LLZTeWqvthVLTjvDJvk5jr/IcSAT0C8UK4pwz
e+9J8LHupl0CLmHivZgWi+Ky14Ym/yTmZO07ug35FlZfoJmGgO1s1DZqHFXcqPTB9e4CkM6Rhddx
xj9Lf3FYXppej4oeauJzEjayuSNYQolGbZtseGpU0dltqHqKvOttdd49rZgFCi7NPewHT6Z+S4Mg
N0mtPwt+UqWn2tVeGtj3ZAutEca6s1s3J9kroGD5EtfA7/E/I7RwSA9q3G9tegyR/lbExw4W8jNY
kimbndV2jeTJOAUYZfBO75lqIm0IrEquUaCafwB9baw7CpMCXmoEa2gzWuHFUCUZwPwOpfNOfHH1
9/T+eO99zweXD/eR23E8kr4VgkNqAOdNMF/RSA7moTuU4vbekKepFdwn8iwVgbGhsm1qNgWet1ck
jYQJ2jLYg0kOMk7k9MW/UKXWPlZjGV+f+5xK1uH42vitCkvzgjEAf1pvNAOUf35irr5VQZ7QxGAk
UhJT0ZLjkQMIIfgglYNoYQUtmgsulnrJvgtiv6w67vl0tHinoK0kO44L0VDGPLe0clqfe4PohGzB
W+WY8xvnx0C9bFAGGs5gbfAlNB+OF643IURsql+cJdq2cqCA+93MUihmBTC0CqW8udDPt9XmyzrV
I4CPv9Bklto0QRErNPghaKuQqKLrOjscR7KXma1q33He2p/lnWmMLkRmI+tft6DpfHrKUL2+abaZ
sDBPyPVIj/e1BCA7OFt+8tcLzZ0/zlrbC8saXfVh+2mdOB3HXe2FgEykbBFk0A5oPhQgFMZ4aEmN
kZjm1e5jFBU81xDWwQNA72gW8kKPV/JKTXbo39JptT8dcmx8IETjFgWPcWheO5ooWb5nkE65NGAj
TFbssOixqjWiWnJyUAyQdHxnGM967J6hQNfVFg60cgVcjx4FnudFdMWUchMChzpW3S4Oy+KqAeKr
mdjgUuex1Jh39OwYj1dAJQ0WYhU9Hwk2VJW+wPnlszqxHcHesoa4DOVRz3M9yLgG9P/62gWE0/m6
VV9BaE/67gHoLhD+7xlBp0LXeuY/Dnfg/3D/4oGsfBeuo9AdAOVMGHrizfFwNMTs+td3WVyiDr2l
ZrWi8lnJ6AYrmzzRTz5Ds2TCgWID0WeflYRFpF/OVu6lSGiamMRJuzvVhUV+b4j0YfEOTRGq1oMY
SGNIzu9jX5tArsxw4G+D6znGZw7CGdEr/VRqOvWBi/hBaxSMgZxMG7lAObuy080+/6DodgW/jYYU
mccGeASqA7YzAPVwMUxpOGKwqciWg5o15iMsfX6+HnA6L1h6mwv07L2579Vfs71lwyNgZS+8dYO5
yA+Ih1dizFJL08EIR33x/XtrL841iPBSc0vZ/2itB4CnsmUH6/7moEZ+r66KWPAT7qLKxYINziOL
gu8bP7fNlGHBPOdg0qPrhUFivgUrvM5HaV+0mcpkc9zvSXHoYOiHfHCZib0v++j0OG1DCKqmLJ60
JZjWRb+Ln4if6027TnlXpogBch7ljPlajcup54G57/KyI6TldlgFhofvFoXQ6Ssa/c9H+YFQeGiu
bZwI/dBNnWVfnaspDlPkFkTV7yCprDXmO+1oDhmn+y3Qla65lc6TyP85U79uK3WZlsOi9MXV93Oj
r/8VL9xzwagbgaAra+ULyfvUUbI1HxJs61PROrv7bcVcRITtbQaxE3ZBHt0A3Pcx0P+6dFC3Dl6B
u2QxJgKeDgLH/CregI6Ot5ZOh2HDuh1jOWNXKnBHhFdNHLlnN+5E0tAs93qR2W5lJperYcBtUid/
mojHs3l/iuYEexirSFuzUcgIhr68QVwel5sNZluIA7abqW7+zkhfH1s1zsUCrrfrlnkA5mbwvBNG
/aZLWweGTnfAklLcT1VNLfCGUx4DEtwSlXakT+Ja1ozMNcbXz42ryfho+9pLOB9piDzJBZxOxBcu
DwyOTnEML3AZduTsWYzBrHgRCObLo5JG9ydt9jAHdWmHzztEgYxppUHNaWNRGujaWxKseWdJwkww
/MnaBuUTlaX5JU09A0D9Qm3auC55/zkn40llXWcbYRrxM7c/lJKvvtOrANb9PLKOSdTLI4U6lukH
X16eFMulxb5uOrSaLhSA2GgtdyacszzfUvyqvw7KRsMpGLZIUEqlwSr96x6/nfFojPPk0DPcrXLP
7Y0fqqO04LArMTK+EaWySPFcruud2Upohq2Azs3HaFJoNIl2rU9h7nxtFqpos6QoungoFo5lZ4+3
r8qPutwCgBAf+10VGk+jpM/u6rsMQXguIX5XiNzeXK2lPvbvxmYoo4G3SXzjE3tkN8sn6E23DzDB
LTewaeeenNZIS46QGW+BG3CBkD1l1W2tjhtQcxvJR5ZiOtA2knBjWC89IdkB1VpGT/WaJLVAoKFQ
mpSeyBd9uiX5T5rx0fEvUECitvG3WTdp17086iJ/zXho/vfFgdGeWLh35oz01DIqm5dKNvtVVA96
Vccy+ylK2trwddZUQtGti8JOFOeNNoAAkA0katzYyGjacUbR+X+P2WQ9iuAIC2Udy/37JL8zFNEE
E0cb4rDO/U72EvhFVYsFQZgOV88+HBMZaF1kZ+fGJlT14Pnph8OWH/jZKp2A7FeK83PjSrcJt2TM
EcXLV7uZcPLBMddnEOwsZeX0AgqreLympsdEJUYt0S0DnKzICKuP17D1wq9/AvVUTSbcTg9cNnuH
sx06HOvlc4B2kuuxJ24AwUv4a8FD3Q6l6a1Lfu4ZXPdWMIx/+M76SAJ3yQp6oq9O01j2yT+6lB1t
Pxj9GTQNfDcR9/Ec7GWyLFbCl/NHAlB6IcK62pzAZgZyyEx5Rl6s9cOrnq6CznRIIGb5NRLx50t9
c7lxpmQaoFOSAa2oXsFmDK//hxudqqkmaXsO8mXMVkS9xX4rx7dh/COSLIb/cGStJr8+asVpFga2
vgJ11UblTp6fTRGGzCoD5jm1ROEf64AIF42jpMabfmn0joc7bDQM3hMm7facSQd2+OTAiWhotwTa
3UrPQLDtjANsqIra7ZDqXOPfT7ROH5/7KKY4Wyir7ICwV4C6bKyXjQkbK4XtgBEtbAA4Ai4wcC4u
E6ego1neXExRDZwuWUMPiorIuP5miSTE0Od2Bkuu4GU9aPfu6VlN3R6pmdOrGXbEfg/s2Sz3Q1ch
uFIbJ1Kded4w9YvieDaFwHBp412sGuX/SSYANTl8SIpYXcfTHuFbPHI2oiXP+4kFe+V8tYB/iCNe
bloBUroaSgkzawzCQPAl+IDpUxQR1/sReugzNuhk9eFEt9mXxseoMb6X+3KODXf0c6umGcoo3s9p
DyYhcB90MFoFk9+466k8kzfsCcGj7WvUo/bL5Vhg5+f2GHKFMG53x/n4VdooaEUUPZgRFNz48P3d
r3RICENdKFNRZxv+cxx7rbnMa633Dgzq54NzIOZhMIPWr8F/p7rLntTe2ISX3uwEKwueASd+ygjx
9ldDpW/0rtTmcuav5jSqwktofRdNiE6xs6zyLErBo07Oy7Tm8L6BROTGkNfZqBq0Jm4JUrmd404f
8SA0wNYeskhRWcuoAGp2tHc3/UkMTGbB6xnJPB2GVzcBDZeN9bh4BgaVzg8InS3JPbYcVdCzTqk2
U7BMLWr9XSZMiHpkG7ZP0spA14CqUlcXlTIhfhW2IkI9Jr5mhrykVTRk7jDSFWLzp836syf92iuO
8GUf3WE93Dc5FMCG1LLDLrPkMLT65JzjUJqja5rqw8M3BoJ6CE9ikiHoZ2HUvT19mTuVeEb2AJif
I/Za8ZTQPRk8q/Dm6Hb+QkdXUY2EhMrvLlw83PEPyRVMXGCyKu52CsAeU9pwAlXBD9E/gNRxwwJa
Ctz5iZNlY87b/7pe8VqZsblzIqO/8PCx+R3iHGm1kuo/iUsuEcEtYPJVkbDWuTdkFYBGn9Njxk03
QeA5y3RqUcGv4gHOxfsCa30ejYuGMkByOkS79kQrUOCfrUab2U88DS3K3pAD4BtpiR8yl8+Irb/n
WgNj2hDNWSIu5kRYBTb2uUr2Br9jJaLFsfr93Vm4L/AKV9zmcuD+xaUhyC9w6kv/v+v3HxaOrWV1
bceTCiBLjhJR8l+p+KbWF3nz8jXZUbFGnc1I/YJDumdJViGa40c1iapYSvw6ZNKMxPtHkU8KpLwQ
2WOz49qzyweyNmUT+ryDwKn7b8fp9/esSiTsj7x8mA3IQSyw7I5o62CF+NeV8+OzzLXtGaPkvc4Z
pyoAR20zzbYDLgxt4/M6I/SAWfaD6NF6D5w8n8eZA/fn/v1KnX+ZEJwzWwlR5WYAOmeX/aBYJg1+
f8SFh3s7MTQUtoDEiLi/lV9JM7GeEWFgjpGATtfw+Lb1Ubqs19kaGOtsyRB6UC/e3omIY4sFRfMB
tl0Q6bqBHTNi0AZA4pamhl1BdySf2S4X3r49zY8fOHmQb+CbIqjy1ZOuYuN+cwFcaJn4vjmH8jG/
/Lhjv8mKJKIADzKmJ+vA/JAAQym5nGb+JARgjqmJ6AxlrqyhyaahnM0q2g64VJXO6u3l/ckMfipq
+C3gulFzZgTEWBbYRv6jKwr4oVnvrvSkTx6ip2PQD6gDQUrQNTrCmxvKLMv8A39tzLwaxrgYnTWO
jhMVGGAzhT/UDo8yY7113SAnmiqCnLGT+5bVrhwa4g2eOJyuaUWfSXNeDSxsr8XPG7P3vx2yebiq
hwIGaJ/0RhHdLgcTH9kUO9qDYA/BKjEv02z5CmtrMhFS2ZvktNwZZJC9h/ajXQPKa1KAZdeVNmQp
hkj5UWRxlmhu9f1zsHmEKGCfFV2TYMklElp5VxCA2CIftEPfEFnkQp+ZoABckPGAROIRowzZK/yc
ulc1yjIkMnefK72h16NsKl7nxMDen1P36hAVKU/Ma7fcfZ4A7TFn/5Hvs/USLdYAriXQbWR48iW4
vmcahkZoNUcKmMl06RrC4LJzcj/5U7xSom46R8OQtCCrof89cT+r3RFb+KWnAQ5p9rLmwnzMMa7z
bMB4A2IaI36NFLHo+2WkMSKiYPhR755lzaRrGG2UqoA7t8xjl9/y72KueieKww2+cwA892Is/UG8
05xD424NX63JAgXMco9QBRl+diAnLd6di66hZU/A8rO5d9cRyB1kMaJCBuUUxDZ8YB8njOYX6YK1
ebZLi23kUCvXSMhdIQPbSM56yHOditCxrcuwtuIuifKMjTMQB9m5a3fDE8/yQeyQ9vaPUUTzQLfv
pTuz+cBcFU+iSDowVHcpJhmtFLtBDlvL8GDMcAs8pzVthd4R9N2vFSb6Z4gYFsjrotCNyyaqNBH6
Cj4Vy8TNFSYB4hxkrEEy4aUr3jgYfgwwnK0YmfoI7AUMzYg3CF71dtzAi8rl5yIdXKkl/Sg2HITf
nlmhIFqXjKtswP5kunoqy4Vc+3zJsnZgXqeHyI1vQ1XVWhaBBLeTxGnTq4Xrsp/Rw9Fys8rva8jy
CA+/thScAQkCRr3oPrUsyTOkOGRvx8aEzgm7q/tm4T2rgnFjtzp+wzcs9ymlDLc63oRm5Jq6ttgM
KNXTHe2HD4m1XYdk3hA5lWna+T1rrmk+aCk+Rd7mhYkG36VUQdms4rEh3srB5/DZt8SjgiD9DAOL
b2lz5cSxRVZQNtQgboDRwSc0U5kdMUXrftlcWtjxPI0yBaCZqtFfEAbgS6C+YXjHcLpyCXpRzSkX
paoXUtIua7E5FK5yoxupwouZSldMdNlaLXZcLg152jlrpj4FQ7THECdEJJoftkWBVwrRdyuRp+pH
P/cgAymsSVrK/n/Ch0U+E6REK60AWiOWGvWm/de6H/aDYKCsc2U3aghvBugGmO8Q+nMgq5PvoQpB
joa3dvCucxSmkUr9Y9zgTT71aw+0kiVsmH2R5/JKidoWod79/eUJ8Tbi0Bifrj1nvkM1dWcXhN3U
L/+uTmA6/UNbsuKfabja59RiuvT8kJgngYC7sZ/FnqhQksHxHX8msRULZXefU5R+PSf4PtTyHoB+
6Gz9YMUvcGpGbogvJX7tIKAcn7SyiKzA8Oq13A8D1PEgEWcvjETvCXEW+DZWdmifYt/NctdPJq/S
lzXU1AYCix3t1gDBVwKlxFpgnTLYEIPpgrkJ1bCfNy5jPjJnPYfsBsUFQkzxVVPE9GgfthmrI5QW
xRucqcTr2F094xvPjhNosfE0jgOOnj3tazxWDOyQ60xiz7OjGcCRGxy/4cuBnnmxmZP2PQvSN2s7
8GiEVc8uA+V8Q6CXA7/JvkX6MoOalXpKHrTZKGMWrr0tFDTPOuzGSk6EXz536cakkBdfooBahCTk
JBs3L/6hYTK2Zby/AuStI+XVXLNIMGHopXXVrfurjJ/qaGqcBVCGy5AVg+Rxfh+6qdrw28PYI41x
G6a2yv1/filPJfxUSRcS3M0NHSZxHju1wf1Lmi4+snMEmeLHko2FDtiHBx59np9h882cZ38uHuFL
PPCWs44XiN4uP+EmpeAC2xKODE+rr+CcKiiIDrjT9vufdPsxq7jcUsLDyhQP9WvdDLxZLfGzboR6
G3CZ4z/MRZX1BF5tei1Y6HEH2fVwGH2lY9/Ekdz8v/IksPnVx9JrkysBLyJ6/v5XYi4JWUE3ed8n
Muwwn17PZI7K+floN41uCXTr9JlmpDLVfCoOMeHsQJv7f6suThCSW+03nfblKE5eSoyR9hoJ1UKy
+dL/7q1ZHIz9aRRSa6gzCwAVTR2OQ3ftVU1RhmP4+phpqwLHTeBpbRtQDdS97zuvEDqYK0YVWzh8
344ROYQHTyQEVct6LqTywm6Qb6Xw3S/j2Vi/9W1vXraxeC+2TMh/tyotD+kqnzC1H5VLEZC7fF6H
2a5MhmVjCzINdu13y7JjChTMOdmgazAywr6k2N/fAU/Gm9VQRtdihuC6x+E5ToHhmPBANg26aU78
kX5sFoGek3iuu1osrdy5zKAASMx8DSy5gQVPcItewHUqQJyEXQLRWqvbZqy1FebgqFF3PeICXaNy
l0K8QrLxUbGq4qUr+FEvQIh3UmA0qsfdcwkVOIOLdvNez6QDNSLZc+Vq4IpIgT6CMfHy+MzE2R/4
8gO9JsVafCWMObGvWNTBUeERlITRgKF59MEw6I50C+xR36nwakVp2cCpXLti6qPr4iPkuUE1f7WB
Ht4Gj8fmwiOTGfNqiD8jQeyxlF/HRkStSSvBSoY7mKwC1FZWVJAxBWPykAQtW/1MH7xZBhtJ+9UG
HiM8Qb8hiPRIOtvh4x31L1/N7G6mgiOFHMpW6fYDDhPhv+9tWU3o3GrbgMbU5U55v3oYBz5it9yM
JEXWH+C1qLuYQQskCNVbd+iSBUczy18CweZMs1LpIbnlOeiK8Ar4fUsXhy91y2Mq0p1WEMicS6fq
J2KLrXL9nTBzet/FfLR3AL3ip7BEeuQjQh/l587E/O1MSlL57SJw93lemc0ClRuSC6SQ1cbuYQz8
GEMCR+3GmXppnxkFwU7Ep/TpcxXmmL747vPGRPQsSh9ehTn9SROU3ZcTiRQFXV8BqaP8AuZk7Ucz
l7Mg6OPoa9GmXTVzYKfDt4jrYoGTI08V8H4IqcpwN15I96Mb5CVrooXhm2pmEgnhRu0vqcGPUZVR
roS5TljARFYW0dqAM9umnVNfUpTimuG4bYU7x7hZiMQQq5GUjUuBV8hBnTkz2kO7BBIYz8FeO5RM
ix/2B7BSUxAGD1HT9bImojsgVlTpFQP5axjf4sluHbd0nx7RQOytRmvaeoD6XugKKZaKjCC+3cry
p8P7eDNGDps+82rk9iZ3zxcVMKYkDemdMA1iKmQ3hCGPWMzAmAcYfzijf9eI6kL1li6VbnsvAWw5
g0FxSASrpHX9MCaXAblr05CumG6v/sr5q3SHbr0aoNhmPQnpL1snS5Z5mbsjOUFIaYfwuB/fV1jD
tMihwWxjU7PeSirarCH3abcIEB+ZVaRac304lXi1asxuCmq6C1Dy+h439Blh3Pd+kYiUdR0I2M/i
ReKALxS3FKQKQhuhgs8YoQ2y9QIrMXPWZo9f6lnGGDzspEj4JL1eBOzB1Y7Fbi/UyAzdamcV3Zy3
De7eUwbxNSSEbUWkq7R8+SG+ZU8sts/VQJBDglsBkkctMVrsfQ4eBYiH/3yN1iY1aXx2/MPW0tn/
5w4bhL4XHS1eF7RXFv/dlFoz3i/zN1jwAG9aPAFAU6TMSEDF35a/VW1csxv1xCm3a5bJHWN3CtQt
XNCspYqSjqGCI4Lvq/WYow7CU6L5HzX9v3AillohRRf9ZJ0Tx/GLUQhZ8hSUEIJC7XtHD44YonPs
UfCgYfuCL8pdB9+ueBuwyJLnqdeCoDEck81WVuZY7ACvPewMtDzpte9Omw7TrcCUgQCWYblgXL8g
G+o3+84sjcFAzSL5mJHstHgQ8ke+RzUsI83dKdmzYV5SA2b1ZtunPvK3EyzoTVB13mqg38jnPzHI
OK+GRzbfJ/1udNZNr+DquxTvifyftN+jdG5W21lSCONVtLq7X6mpiEgoLZrqHSv0STPDKNV4dB77
V8pj7e05L/QkYo/oR3DDm7EBsMJYAP8FBoJ8U/x18ufrA0dE+UayY2hWEhlFBgaka1caN1qY4yom
hSm0NKWfZrbMDR0k00vbN1A/FOj9AGZlRZbijIAYsVlyxKW/+3phDB0jpkHkS+sP3oCHGvjPSx5a
6WRqHSo7oRepNPnKNcNdCouNme7AVE+cH6bkM4fUSfTX1okpdcPrnU5ua8zJ7B36kZFuJ8ySw+Nn
M/j2qmY7V09euig2CYpLelk7/45yqSXnCsW6wf4kVr4oBpL/66WO+BlJRLf8FhoM9NkOdsq2Fcky
/rifyPX7I5zIWFe89ISuzY9m6yQHtaYVeNNk6lv8noi7y5Irx5ePXJUXllRX5RGE0fPIpBevlYhA
eJG2ZyAY3OWLV47V6ijJTxTXelPzq+JgEaretNDFhZ4yufxsWSWmCAKnsWvX0dp63KGF4LynexGD
We4d47vCrdOs6XhltnyuP/ll7hJZz5hT5NA+gbyiKltpO26ukb2cldLYxQ/lp+uZ/913BiocOsxq
EeBP5HxyeHLl9NnjeiWvQ2cyzxdp/mCQPtfYtyAS9uVhIkXqe6fFw7Prrh1CPT1FwEHDLWYbC3CY
NLIRG+YqBtR5YRScQNOw1HmTorLEelPholrDKchZdaRq/LbsKUGsGeRFN+N4r2GTTBpD4nIZ3Kua
uMm3cIZjNhfiH9WuOiRBQc4sq7mb6mpLI/lbDOxPiaprbspaOiZ735ZISTyTzPgYD1fDkKLO8RaL
a0rGHaCQTlmOn9htxAoVko+YZB9d7EH/3i2aEFycZYUrLjjrCCq6gs6Jd7ByTSCq/RfOCvtogQEZ
y1RPlzY9c7jh/3rrT/ow4hPBVBYdGWHZ7Ukw6zVdVbdiP/YTcZ1b+PEO4cy5ZsWZ4EYij3+M1lHf
7jq/AaceEfREruUwZdSn9Wm1K+D1/JzmJ4UrZeZyvTyLVOpn0p3DVhMa9xdHjaIAA3dbgOyZyRgd
yq8Fz1XYBv/IspuMcKbuXeocEztF5TCQY/NgoiUHCw1eaNCJXygqO81622WtxH5NZ2j5bsrsGvpU
Nn1lzv1DyX2hK/csCAF/Y/6WXrvw0PVrRzHso6Shofz4uQ0KFtvP9DQf9mv5X+Jz1zWff2KE7WuO
7yaGgJl3nHj1Q5jUKbXpyEm17buoymQkEWs5DXjBw4haUTDB1zSkuWCga0bnoC0pwuX9q64Dsn2o
dK2zJzO6V4vKnvmUo9fWtz+6rWUyi1jNw2tm/+2S7PEaZeYog77Aw1rpFDrvVb7EksLDD7q3T/+3
47tm0/i1WCpSPFzckyWAfP8F4JeUu+SP0kZ6E+nz5ko0QOtaYAGbZtqXbrKYV6/5s+Iay5qmimdV
pgB5M5Tn3RWxt7ERegRoEG64+QC+4+kp0PNad06FrsTi0Vgr/K7s2mTara6Pn/Gel57qzYt5oBnq
FPu0iXyjTRk2jIHCoizSqrlJxXfI9o8ID6ZEBAHamffdfLvDdwwYRJPZNKPiK9Uqd54TJv98ig4T
9Snkfh3TZ8G7q7ziE0MkGEMfTsKrCMxofgQYQjNorIDtk4TYTAo/esvNCQyKiICjpAJ06cKNvKiY
SlRrPtUzQKkteSYLrU4Qf9loaUuEdcXoXJnU78q3u26GhA+aZsbTxVYpviyLHqJvrStJcBRc9KQf
pGOIoHePElLXgXmwEtGkDsivEBhBybGg9RUekjv+5uUpmklv7bfj/Icxqof/DiUe1Dh5r/av+Ex3
tTbPKQeWt7R2DIB+aEge+smE9/FnPhdSPCsJpjwzjaqOSi+W2MyJr8b/a03UHk5olZUmQT4c/tSo
5PyBqgc2lDYjvCZ6sHGJeg97tNZkZyKxwguay1Y0FmKp/kxT78aZCEYItixmXuP26z6TNWrF9kKc
bU9QlQDKXU2tBOU2HYTm/er59xsXnefgPyHPDIYrL46sQj/53MzYSrVR2/xwXrg8nijBXEYaWWBG
4pIBgt7sBY8pOu3g5gzG9ya9r4F4xlrBLpgdddZ9QKTuIvnejotWo4uzly5wViyu2ii14Pp+th/n
YEQXghxI3VMGwMA3MDRKV56mh3RtN8qvfsr/NVKaRh1Nn7DRgnxxeeo2zh07oNVUIDIbnIp8SonE
Zrf6XCr52gejJlpvGS6Y/T4JB1YTks8XXoLDCO00q6rUlYOQOlGW+ofJFjb8359tSsRyXYcUoV2a
Yi40xZPSipebRm0K/HXXP6EK376QuHxjrUUkpZNV5p4n0KcVPqmyztTjs1l4dZeqEKGlqgYXvsD1
u0Fe5KrzpDq5nVbEC8RYe2s8UjQ9ArdfYAIjtoMcz7qnkDnMY7i6KhPUHYjO/UWkgFqKFdqy06NL
Yg7GMSVHVVNTJgn+CQ4ucNJsZruVCkAn44V+bCvTnygV/9x3zm9025gL6PptXTk9uEbmJEmqsvKR
84YnA2fDCFDI8Xn824JJ0NQjDjzohwg2eu+6do7Z2tpjNzJOeb/NeE1McxHjZv94O/1CUDgkO+XA
z7x4aF3U56RSBykCET++aTW0+fJdcfXmp0DJAgkV8kAW7JyHAmwlJMVDteu6fQcXVzTwo2ncUa9c
taD0n5w+OhCh7fFSZQMh9wcbjvkk1GWogY2/HJKKN90vJ5F1InHp6vaTf01/SYLEVTrDsUDvzlR3
9peNWVNaiyxfOIROtxkyNlShfY30nu0KW/8UYXH0h1u79i8uYtkjFieiPpVQzfYqV4bnzcJ7LoQj
YT7SUHcF5x9YEcsW/rKVSSxUypoNaPDmXd0rBoVGAQiUEa6AAg+iTeH91EVvbnRykrBM0SRFYDeF
dAJVfRzSgJyMa4aJoWKBB5HcQTSNTs29fJckLLmAW5BmmGRqCkQ/i+ULI69+kUi/raKnT9xy3Ont
aYiJ1bY1nFpOUCb/5XV27836YOA1T0pbwx6sYt3ZTfEHQIUjSPNOLP8dIGXDqaFgaI1J5mxHKGpQ
UhdA0gLYLLBwl/jeVMZ9TJ24MqnPQ0bh9j49+CLKeuSVNBT3br6u06FJcsOzFoi023KhCf5FIgzq
F9G7Kjaqk/D9HDxbYgahS09VjVPIofYmM05XlsHrwyzD+zc4s6af863gn/5G6SInPpNdXxwARANS
QuSGDRmyxT7NGle8CgjLL1qqc5fu60JtdFSAk6sZlbpTltNmS3ZeFCa0f9DBVoVINDOecBbbyyg6
q4gGLJOTBx64k4ARC8WG6H8nLDUdOnIlivVc2TuFkEW1VqfWfdoxIZLBXV0tKiUAcMuIkwqwyeYK
+/ZoEyTRkaHfbnCbHmrvpBHDcM4i+jJhGIJOv5HEUeSoyrD8GBmnvMuk2DcCHsNOcFE/Z7KQmQSe
mUZ26mxOSL/Ed2mDw8PcA7iLSixfIsrtXSfarjtsoCth3JKFs8LyIlfp/8oHQM4yllch7Br2GQxs
ps/u8koY8yLCzmoyjCGB4sZQ6yv1qQg9Q6CSLMr1HoqJZmpkElSVRgVutssgf6YrgkCq9PAxx+3y
oiZOKtKbd74zFn0bTZNJUTdGXe4XOD5HwtT5qi6v0Nevicz/zJGSIJ5NtbBBm3U6vcNRG4AtuNh4
Hj6irMvi/Asx/b/TrCNBZzH4BJSG3IaPGFMxL3weeLSekXDbs3SOpk0XSBtHljiRd1Uq4cKEtjdW
5UmHvx7P2woc2mOPGCW3hr6DxPQD2QiYt5Tc3MKfk3cBWo5NObCRil34wT0eUaboiAM5ko9khTTs
SeGFvAOrT/SJT+jeZVtzbOfxXjiOQEAqI+LRVgb6GVe64eZp7SmaCwzpuqHp2YkQRB70GigOiX3t
KUehCvdlC8cu1nuyG5V7qoZWpA4oR3wJ6a7KhTqvdm/3pkl0R+uZ93IJY319byGQqHtftzkGCxXn
7OIBV7rx0QPVC15MVgejZ6tBL6WGI3yfcQDsux1mQ3PGMNGyGqov1Sh4nlPZt8R39W4VXCzPkIes
QGY08Lr58k4wfl0Gcg8WjydowyzYo+ccIWujYdrMZJvFwP9xA3O4z7F2vuf/IA67JB2tiXeXD8xq
Kk1cVD2jUIOAC0Ol8pIANGx+PJL6A2kVSh4e4sV6nxsF49XOgdvHTzKVUBwMtEc2lfjqvCbzKXV7
cEQYLsH6KV5vT5DkLsJdePmo7JqWpKBQCDAjMSlYx3EMx0+dU1zWNQpqm1PhrI8lNDjoZUIfn97V
+rp4HlfACF4ojU2ZUQ19KTx92NnMpJcRy8NLpRR0Ebr+LvAe2lPTCVbOr9dgcsbN4hGa7l1PpVV6
D/Hl/+P2wqwOI2j9X4Dzd34OLTUV4nTaK09MeamBEvwbAMNYB9ZSRmC8duga/kpoxGSfIkDKXQ7N
kV4kbSsUO6LZRRP1CKeZr8NeJdRf7PI+XsC9cezEL26+JWZSnXFqkSkM7i0IFgU8tHz1EVC0+Ii3
khLprozyrUWuFppp1RAmldukYO6vGSiPTDYJtdCa52t5ydSrgP66856sUmZSBlHP1xJboZNNaVnu
jV88CfzVAeaqSa1lMEiQFIJhDvTeBbC9xSWJYrZee/DJBBJGtO7DFP63wL7LBS7vWKIRHeB/TGCN
DceNKi0dApJYqj9CX6chP3Lxh1u+nEVxntZ7aM8h3S2nVxGSVcLFey0AK2x3aGskEo/6Wh3zbIsS
Ro5TbPO9cNEWao+qH3udB+ABNH1MqSmgnG5RuYcjdpA1APYtl1bzXrUWIf3gqxY5VkOw3hmyVwC/
T0df7LqcWoRhzTPqHZpeJEmo9l1rM8nCbrwOXxyd9Pmuh3DsPNa/yJQMkpe9nHRfkdz0EL/qDGjm
W0/r8fphPKXffV13PWCiI/gM6djjUlhK7xdfO+XBZgUoCQcLW51XgkAt52l1lpGVQtJH9EIQp3/+
PryZC1T9veKmk6Osc2UZqDDeQB2qvPxm5Og2+9Y9CcVh1EtVAjoLPINPz2N/UC0kvvQdeFmOSU47
mgnzkh3wnLGS5skEgGvpQPzjZYCr0O6FmZ1BDmVXi/IgjKDx+fLzAWTZKyuHRewBgC9YGukcx76N
FVKo+4Mz9EaJiBrET0DzOkymbrfEV1J+5xtsR35aCyh5YrEUwrk+3h+qlirKEtyERKjTr+7ar89S
qhtxlU78Nw75JhxiX5nnL+0xdYfslYJLLhjnfXx4qxqzBUEE6MXjtRoiETve1QVHQQwDqST6EMh5
+j2R3/cdtRsjm6Fo4xrgxavyyj0yD2mae/SaC8uQ4TugpRUeXqPGT+ikmD3GU1VL4lvhaqORkweN
Qiqs/MlqaWkl3XElbVLWQ9B7F1VpoFmoW6jPn2/XMQgQmEEy0KZeTGpO/oHanQrmTOaapqS4p8QA
L2wZ0RnmGK+hbjhktRcKYGEZGfEUfMk1OYOggytaYqYd3VemF9J51vV+DGEKB/XEYV9X2mIzB1FI
XDnlR4CbO+uF9dZgZYM1O66b4YLHC0PsmuXwr7SIDM8TTonR2E45FkvTRNqiNs/BujNyW+YOC6lc
4uM4bDTFWIHce3FzprZbECpvKdJCbJ7Rv3rZoujwxaFMu5D4mr4fM0RifB7MF8sHiv/U9P+qGOEX
EJfLTzDHg/BAvYRusROr8m4dxZbLc9ALXrlpmW60dz/Pr6yL4qYi7CbkEbB63NHkMXphKJNYQTcP
7KqPAcWnhJMfWzn75yyJuZvaI4yEXHd5nUzoy3hji4A2s5hD5N8TADU9LK++QmTtNQJltwxlIfUq
TRVEZOc6VDCvZi4cxOmA0q5XRgzDAaDBuhuPm2uMXxNL2N3Tu7JpcCv4PaBG6xL1SjyfrbMn0ZaH
GjcvGNEhwkJMirpHeRTigbhmRWhLJh05EiXy9rlkyAcUCWw4a3k8veX1ad6PmKX6q7TtbZKA7yQ8
Yne5y/keKYLHkdpqcvpavdf/G49ItviG1imOE+GE9Ey5B5rVqKZMIc2CFB5Q60h0nkom7NUNbjWD
Apwe0iX5THibr9kqlyD5bBHMnFExAuDTZjr+ZnxNI+8hqbwoYWCyg3qssciBGY0ABVu4LAX2YcN2
FrONN9ORCwzAusCxZxoRewNFndtxhGsyj0PVj0faXjIpCVft5W2mTxKXBC2jsKcFsmiwXUBZOJpe
y48xGnXuu8YjZ7J6lbqoSEOfTFSsLX++ipIogDxzxBSAG8SqrSy07AG4BmCZn3IZB/TDWb1hWNcW
JFSmGrJyx6iD+4yexO28UD5PsbMQcl9asUSWFBrqEEDYAKcr66PJ36WWq2S0KqwCEAkDY/mUyQkO
JGJLJTMuv+nYItoKzUS2eH6UQSj9k3Zl3Hodl5NqrbyTc0MBGebb8anuhxDFVF3p38qjlznJpKJl
VVnzuVfs8ujvtebJ+bLb3Xq1YKCPScjbnu81ndT+frktX2vhu+/M3S4nwF9EdcUnQOqC3DeWCFZZ
rKpZqJ/O8y6c2yxTIfCadJylvwUA8bkWCN/NoxG/bzbm8pyqk6mjVrggdUE9OqU3Qo6WuHjQpkqN
m82U6L0pCy9wROrwXaqxA+OpHRH/FWpfziq2qR9Kje8ApnjacYYKuWI2sYoa239KwvQZk93eG/KV
d9y+HUf64CDOg9aOwrnnaDswzSKuEt5Ld2jYtJ1i4BX2qV8GejA/p6AF8i4MFBklD/GPKWqOopJ1
ZtNZSliPlOU9mOYNEuM0VOK2iZm8MwchGxUv69iNPc/BghkeNAsy7N2FCpg5JWs6Q25FnM8anDwy
KZXNZ+mdNR5ox6KUDBLdcJ5QI2ULcJ7m9MTuZ49iA9HGqkH1QWRJNBfW5N65rmNGgdSIgmVs81dK
+McMkb6ZsL2X5dN+Wu2AvHfLs8BRyaisHLvrtlygiB0lzpSu3TjaCQXV6MFu5lde4TVgeP99qNfo
HexVY6LO59GninwXS+9NmfkXNsKsQydO3S2Ua8hkHy2t1dWoFZua024/zsACxl3OxcTcynVj9kFG
cQjIC3gNVmf2f4orTXQ7MoPm+9b5go9yY9lCylXZB8bQYL+CzgIor98DN1XRlvCDVunHuk4ftahY
A+QB+naAjJZFoldTsaZBbkfjUchoi1PMBjOujgKj4NTGBcTsKquEiBXQdVuzpElalC0ys0oY8bOd
BztwLTIGuzSmbpINvz3LcuL6wjOWAnF6kpQci2l4dNMcC9rTB0qwvjzslpyjUJg/XrSNLMu/ZIwE
aF7H2hZE++G8pGgaFD8u14l82uEdR3fxjT7ynyVeJUS88NhGToJnKvfXcWkcs7CtWJRhfRSEteoi
Bshtrw2g9evHW4gCHtYaVXFsQKVWXpiWnzuxsanKPlxsuXxhZHBfROp3VmtLPCueDpB7z8tOpp/F
rg1BoyUayjppEBjZdsH2jbVzCK3efLe4bkelFrw21W+9STB0Nk8Kol5SmazbFncbx5/AnZou+tv2
SypohqnzAstADb3a/bVpuL4RmPeI4B/RFCld1+wcZom3EC+TVW7ru7qrWZ3VMZQR86MDA0KZLvgu
60PaOUzrvr0PTf06wE289yy0imWiDi5QoEhuPKbxJcdDHQENqhDuft+DyI6YBpii1We/hwjzrsBJ
0NYw9tNsBgsxVu0vVR03+bOxY9yiwsBz7UegZR5aq3d7G27AK/pTPT9cN+Q4Nz3bywRpTRINBRZi
Ou1/oSaofwLM407+3yDAsOmo2paIoCtn3X1njBHJwofFCa90RGhF5wZVLll+xsovCzAulwRkcn60
5mTJuhOu05MefELJTKBoZ8WrPxGDTz5BrWbYJNzB8kyCh9XxPSqlF0R5r0QDiAEZVOS/+IP34aSU
NVAInCMsgaLFmNnOelo9o0lWvJ6dtWlu3EGgrnWk2K0hA1CRiVxbM75JRF/bThiUn6SW/psSqJv2
NLbPeB+mJKkBNb9otsWxo+th10O81ecAzogiZfeuQ0uG4Y4qjtwvlFX11DpL2XAL2Z6ux84ggQto
JWiK1SISJzNSSAA1vBz9LCQEETdbKaxcfWvqxaWsvYVfPqgoHRBfBtDFMNzEnkRPq73TfSIwf9cj
7lLgVmswzJVxsVoh16bv3R1xEf3HeeGC/azEsztJ7pf+RVwphqqMn8JVa43gS38WLQ4Kmi3is1gG
uhFci0sWg/FCd4QCQbphG5W3nJntBptmQDlfnefti/LCKY7TKUW6o4Hx7VnFqN6KaFmCSSRDg8UN
tUMOTYD1wrBBqGADBxz/UnVTSgujGj67twyRJW5Gt2SC2Rz5+lXhSnUCv2Eh+K1cLpz/Q9imlHAf
pSJhevFbMaxzzlUHbtogOWOWU0kBdNUl7CT5/WDLDXJQb0F72c4ZZ4tdQxZvFAmXrPTYJo36OeL4
Exp1LN3IcScHjOWltZnAaU7eMxJSAdKvveCgqeBBmBt3RPOBp5CZm3ctZNs9dsyKIHzMwSuQfDUz
40OlMmhkKrm3WoRo+DwoGeLqKzsjm42k7nSvRywa8Hb6sh86CPqelF5ayG4Dr51NqiMcIJ2ta7eC
nYgeG5YZ0X920aAGANvxvC+AIv1NZbOqz0Rd14ZdItzhINlfQHLyF+VsWzgV/wWq4BDNVp0ci+QP
RiDvQnm3/VZ5jxyTkvJSIkp+I6bQml3OnkuMfG3BF/DuPu2zJMGoFSOIybWmL9onLwG/BreoSLB3
f7VoAxg7tfybLHw71x1y0vDmZZAh6o7gSFE3Vi+txCpPVdF8PDdhC8osbOy6KclB2gk81ASSfxQt
8kMOYFW0Y6xWG0o9SiENHJXeCWCyd3oOjO/ByhtWoubA4FnNo8CK9iGVbBN7+kGcZR4JhkdXmvsY
oKka8t3qpgBgkuJhUE/S+T2APKu89VsnBf/durcS5v0a3pApYyQOnSsRibYxksvZMD8zQ53NYZnp
ltBpSN0D7VHdLAC2h6NGklEx/55hwhwYtsHP0PfnXm/FJS8Da9a+LgRx/ziIEAY3axh8ksCATwFh
4gkpNb+BLPPFYvdnlj4IzfoO7nszs/LTk/kgU1Fqb+cCWYd0uNy+nJCAOGKl9JQbh8/wvg8JJ2CA
AG9JEmzm0GHf7VEyCgj3T8fuML7LAp55MO4FYSus13suXq1fNCoEWPUI1IVcm7TDCAHgC+tAHPLo
gH9Z7CuwHNmoEVGDQiWQBTJbm1ekzFV0RG6N+yOknAjrAuhqMRkVXc73Kwz+RSZ6tLJOVXf0ho0O
pdX8kg0WaJI3qo6blhfB2gwQD67QGlCUY3oDuaC6HsKixRjhebdWPGl8xvRnxZGkUR6JUkmoa2yu
z552fOw6+LoCae/hEDSPRI9vstyEnam9LmQJqEBIznkqRqNW4wmj93/D4TZvvcHKjaMYTsvRnu+y
zggHrt8RzymnvR86cit1dKhE0uM60wFkz3JG8JSP8mWCETEZmrxoc2c1D5kCIKcaamHIeYN34XUn
Dsk64hnLxcRF4VOYf0mIkMxhv8dGMggbqHPJTwzjflAIfYtr4O2fG7vV4PsxdRseDu5GmEB//eua
zKP9tZO5v4WHyzCg9r6YmRctvMq2KDHhr2f+CcUWgqT51GhGD9DN8ly+jN7JMVYWAuAl/hd57tnd
PZhJRVNAgccV7fjFrt1i+CEqzGSP5xJSc9yiwC1s9KWOR8X/SAKxvuhwsBfhj3ukG+HB+uGq7r3W
tABdxCCpsupmYujl+FoKQ9GazsXJzFX9TjC2jvJJSQou8XXI1JTptuiYqHffw0nYmboZWSGNtPJp
2/35t5hYOTKWUavBcC94uOE+gNyVUgGjC4CwumiMY+6a/Fg2u+NRD1chf/nUJv+msw/yfeijt+KI
VHOBdClhryu0vsLSRT0LhCpbmCKXEomvWVCyCQWcespTwC0FxkwRf29bKDDM1d04BxsUR/aXfAw5
kYeIGdn+b/nBJPbDJc4fHiPUE4YQZpLHnW/2qC3uHQ4ioqgP5dDXGwKLuJ722qn3tH2uSRr5SKZx
ZwjZ1vlZXgJBi3h+asWWq3ipJ9z/z3+Y0IvdigfxWDu1xpBnw99gbbgT4I/d9TAvVHbbPeyiaSTq
8wjTQCOsx4PfnZWGq+ks5iC4iqG+SkYuwcpU8Y1l4fbqUJBN9Aat6S8ZiR9+OnIEi2HLJaPz3eXd
gv7ufK7p8/kaj/0B9jojBgPh3hZ+IDQyLRbZjECwVkQH9q1TBDge73+s8HjhM6Ef9i2gxT3KVRMn
YKlSE5MSp92WicsX+9V3BytO1iVKIvkbudoWM2SAh01/IDWNtNJdkDtdUKVTnNct6ZZpEY9paCMc
wcMzlxSLiucuUbRTEmlgtVxpjzuwMkAoV8XfC0UmL0QIQXVQmEWugO4IfLnOynUfWyKVvkbaOCFT
5QLiCvdkI0+oMuvavzKnrvljEOPdsbtfke8tVjADvsNndYo+O1Cntr6tlNxkE6nf47vvYkQ7xOpv
sOeGm7zBHfzGNxyFFfJw9BlWlNA3aXEbeH7mrexS00nWPsmh6Sh78/V6E/Djh87IV48IBQkmU5Lu
usCVZqmABGh1VsfPrGC+HBAPGx7eioWiunh+mp6ghirT1XvMGmOrIL8A5JLSWzKfv3MpfXN0hj84
1v+JYoo8YIA+34idhn3h0+9S/K0Ips4sYVDG/XLWPbFyAD3YsR9DGX6+Xl6COI4nFzvdkedv+NVl
YqsdgCLaHbSfI5ISx5ruoJ4oMK/cEVFQ1fkjuT+Zf/5AtFwBh0Yx5GFnIse3i/KMb6IapkVZbGLA
Lyf9apatiRLauXM038+SrbATzrC9EzsJUhlSqpc6pae2YROfU7rE/9uEhZh5mXuIsDS2OgAp9IFL
Ifs5FWWdCTj0nHav7lLXuZe4kSi/OfVS5MKQobLpxywkMMKlIvmvKP2o9jwPLxVTKoUWYWXUrueS
poCLVRD0WUWy/2W33PAZG7nvMlmRrjuwY5rT+5GWNYhWjSIRZduUfc7ttpW3BIT31AGSv64awj2j
T4ou1dTMg/QcLSDHcwmM8NogcVXx0Q+BA1LOd5sVUQp26HQB/QPR98KgZN/wfIiN0OPs4ewyIJNe
pi8hGrYkhxBIeFB/SpRnqewIUvJsbR1V0axj3gSWa7siOn/hILzBokwKgUdnFTRJt9pi1LjfDtRx
pc5UE8O7GNZf5L6DNKwWSRj0hvVfiTcOISQ00nrHTJAi5FkrRhlvse+RUVWk9h+xqf96Y2h5k+J2
5hkXpx8EKb0Bi1ZJ6jx3eipEnhXbWAWeKBFOFFxdYEoagDjWADaFnFTVSm8/s/MNwmTrWRj7yf6t
3dQ1BX1o6lRKymjZcH2EBrvAtgL4CqH5fklw7Gz5+bmXMe8n7UpmaekXCfiy7xdpRTB4Fl104pzb
zeDO0eHfQZuJeUlWyigJ/Ugr/qqU/8YUV2a1WkidTNojTIm7FxdUHtTweVQAksfAYA0bkF53/1Z5
HElabIRc5Rq6IB+L8WCDE6/So9V3cOZITfhWwpCzdUnxFaZM78keegtvY5k80nyYHbkit/OdSeMQ
XcXXUDpfcb3rf0o8ylkRe8B2XNCrd62cawhs74mvvA1uTX++Ski41Tq3BqRgyDxDtKbl6v/qJq+a
6qyh+6crUwoEr1OTz+Ukz38YkQ/UsSwmlmt3LYYuWbbukoqa6A/NPX5mv8ZHkUfmRTkji5TZ9RW5
Yp7NZLWIA7l7+7uiBl4oaXtGHR4Ro9jD5fcduRnRmlVsXBfip9AjHoeNEFGi3JXLKdgWZ10zUBKs
xa4aEaCAOtPsHT9NB0gnKAuKSOxzQAznWxNHdv86riWD2ooFPDxKeiPQW/TQsJzl8Xus1rGcbW7H
kiepd6sBij5gJrEqBR03Sq9SQM1H4nWW8d4sBtH5goIU/K78Hjsn0CYLWR/jEoZeK9HuwX/30qHC
JYvvtpPdSuuTJvXPRjVOBq0lSaWhivWUfC5oOYzVK+jgU+rVDkTPh4poTSmO4o/q6zG8Sy0m5/dz
M8J/wvx27EecV5ZtJe5zlIWic6+lGNi+oVzMeN0c9tHmT9EltqTIpAPt4WrLYgcsdmrRI8OukXhV
jmnkPq+NG5pMihCFZX7RMnPHwMilFAYDClqzxD3kWtUNoC1t/jXMNKbdGSg0t8HZtuFvE0E9uAko
LtiM+lsrRBqMwx8zBqm4FdvHNkxXaJz9oAn2ilqoEpMB+X/0AYD5YAwhjfanz+6G3EL+sKFxcQW+
YJihwt6noknjdWLqvJ8Q9k4eVgCmPebi/VoeezAhkVJnfkv44Ae+pj5wec/eUOKNw2OfDGFajm7Z
2xM/cXFQpUs18yzdxhNNwttTR0YrIZ7YquIXvzPdtBy770OxPQzmVj0KStlL1eJhfOfYoqhPV6sH
M2UNBBMlI+vpRmX0+fiqGeV/uQqbKahQiPtT0BMdYaRvy4LNg0srn/RA0woF8XDTT/ABrV0wksg6
TWgm8K6mzaDNeNfLlUfcpsYmKqk5SIvQR2FDipyqdQLlf2et8obtFwEc7lfn9n/8T+eCc6ZiSOBU
z5svC02TtZTdBA96qHOPd/K+3XNagUXG4dMtX38K5/YTPMHhYS/KHGK0H7/P1Uaui3cXxIx8mS0j
8A9DWA6XEzwRFgDaE/E5vW/X7wFvlZuegHng3M/OyUQc045a7f7pzXRhOxDg/975LAAie0tAXQPi
PzGDJvsXXQFNcq+7cE/3jBKLag7j5/wDvApEBSKdMuqyRQKHx75M3JzKavVWkKmnrEfBVqSzj6Zr
mrtYLgvKvQni1PNvxyzqEyRb+vE1RVjLgn8oCscWimwtJrZUdPHx/X7YQ0X9udk6px5Ic+TO3+3K
Sq/gNVA5xnwBFUrVMUvfRwkSmTEvEQ88WD2ONsYEJDQ+p6W1M9DawXHVGU9f79I3Kdg2lCPAF2uX
6si9453q+/rk/T1tdePZ9rog6QtrZ+ghQR8ofeav3inSLwITxE6mqB7dkq7lpCL2986Q04hmqo0J
Tjlu56F+bEgkc3zFKxKSsfi1JiVU+3Pj+t67EAHUk2bfu5kqnl81rtEkIq1MrLT9IL5tiVYJYBum
fSlj6rApOxbc5OsVGavksCzCuaLQPaHiOztTSNgkotUimCs/T7KRw7ARRC8jiWYudMBE0E1mk6BW
zgCgWRY8dPdBidAfVKVpS+t5CZrFbp6WPAlpbqmP4FdaCpWcP9X6qOTi3S+Qxm1Ng9AWgIY32rv2
kdKNvkFYpGwiqDXWuO0lOboOt0kPcbMNEkA2NZ5bXODYX0RlXzoxrwDt14aGUraMmIHZNwS7IjDT
FlELelgGXhOX0SMm8xVQ+7rPhjswQSRps0QW1g5x8DHv1wwflAQDWxPpRKycThqYINZFX+lhjsTM
dWP7lsEYGlmhuzN9U4Q9EbQ5+IAmqUKJQAc3uCNfzoEtL9pGeyS9guEQ1Mn5H+oAz+L1SxVrL1Xz
+WeMkCICErboKrHHAv5vsa3NKYLaHs/S9osUWAfLGBQ+jP66YLPkOIUY6SvEfeUXPcBPyZzm2Bzs
prQsiPSHIUYqdwDnez3kcwTWREbLLjfHmr4+gLpG5BcIvIq96RNBtOOLti5jj7DS+fakZAnKOG5Y
WvXUlW5bRxrRwrb3j+sjvVEFIGNwu6peZorzNcETS2CsjyTujuYPZPv7LKxxKqkZh5TdyMaXIH10
37f6f7aWu1gYGz4xGQQD6ebaSOr0wDGMj04P0dPcNlaaPoPUex5CCCnDKfa6ta0wLULnX7czTKg4
nZSpyqsx5+e64d+fNzRSgiiYLiQ4d1zvFzNOnVsCSUtkbUVSIXFScUO6Zav7cu4mLPZd/0eD3igx
J+A8NoRqNLmrPHvSHN/ZaHeTHMGIIiMPY6YpEobYw8QLlwqsnr5fkrk10gWA/k7F7CNhONsR9Eri
8xSLHQJcSQ9OmaqUUH+DOQT+jnMyqYBiYMq/Ok0PkliziqmMPeUoRQU/MZfTpG1XIewcL4vTd4vS
iNNruQ+3KcgqUX/mUDkuJngar1r4IspfgIpoa2Z9cSS6MnPm+s1mMD2D3/wtqn/AgvZ0W6yo8bTC
Fih1qP4/gZQ6Erk6UNqQJrcrULjyRnmV7jZlFLTy1P4t2OkN47RehILwuPt2ypMKG49sBlfW6TtJ
qNrtp0lG3qUHwd0tHfdOvsnYNun0VN3uxByqwPOb/kWkzKseshSQKuNkjqouyh9lNE4zlZ1X4nIN
VenYdoZ43hH3USSyC2Zv9ljRsvRK+K4Dfm4igAvpjdS/I3p9L8IS5KGdC8lwDPcrjdH9c9sbpUB+
ub0q7607SyDzrmL2n5JlFci42/L8u/BEDQx/vCP3tpWx8gBmc+LJZSxnXn18Um0KAyBUQItmWvqb
U0C1abDph6Im/M0m/n47EC7dJiz4Rf3DrBq0V7N/84LnTErHsNfJdoOZ0VIFMbgtFCN5sqRXeATz
tZjzjJdbchCxc/e/5i7KWHoqt4orxdvLd3P7J2Oo1rmOECd3EvHCaW1FJS4tk3XJdtupTFMHp6a2
22m4VEToG+wHVq+ZAwd1w+zWj7gk7Bf3OOO3bbyi/BFLXtjJQ/jYbYmcGJ1oQ96Y+GmImtwWw6Q+
8AyjPAQEgzIlHOVKihhLl9l2GdVd+LD/k8f5sQAyWolnRT7VP4W+s9CpYIau/zzEhLgCG/gLuze8
ra1nUj1zmMewlSTfBFLZNWob1qDF70G++LF2WaU3d/4qLjTR2pBLr4krWgvE+FwiINv2A91BQi97
2tyccCrRY4pA2qoBaDakVHb7cgZmUb1GduBBRulUTf0PrFEEKmJiWnQ2VyxYVsDCw5qDw0vewPf3
A79RCwLB/gWgceua6aXw3LhltTpi5zlfLmvZv7ir43VeISoGDjiVhbxggFSPvM8cJCQBC+d24uSX
c4WRgJLsxKSR+F16eT5as0UwO9vD/oouvx836UbiKSd6AKGecnEmM+RLN601m300teXFFDflBsyM
6bub6UzTTdl+gMIpUtk9ZFwJhWtksxRZMR4sugQOrngto3Om65J+2XNT7CuH/cJODBUULqaJEbAE
EkptYhZwRLO2XSx+J9w16oaB+3RfMVR8IWiE1AmVGuEP2svCqIm+Jyhi2cvsL4JN2wDHFlpdr4Xt
AwwQRo0/TCTxVIuRHprBUhsrWNQF1a+6rx9vOaHKB9jjaVXejtDrgWAt5o3G+jVMTjg0BOFx4y9I
hxvXzo1yuIi39i7Z6nt/bNl3Qxnhp+F8479jPAZJ0gEnakYiI2a6xJ/zc2br71kYb4A/pu9Vv15M
4aT7JfCrohkhgHgoBPRL1oSc74p0uuT4tSkTXodRzmGZtZ8+rs6zDkkL2n5Jgtkx0JFwjrzpUF9T
W2BEiMbDRin4O/iYJrK838UnqAupqkAJfNkCy25a9MOqaavFiztG9n/vr8y381acN3VDphewZNYd
SGL0m+B3wNoX0MPOkZM84sk5mQd9r8wH+yXW/diBt/sYwH1asKH8Bez3HUjLcU2t5zzHmZDUaQrg
4dTbaZcMY4qNJkYp/xX8/PESQSq86G/8bQSHDbuey8SG6z1ReyYeM0eSWCwzfgBmxsPoszX6nxzF
wmOUI0fAakCwtqHAIM16evpaaPivN91ykh0Y364rgkbRZIkGoV06W/QPwsBJr1oouPsYI1AsIx53
npR4UTivSvA1H1ndRcHcSCqxOmdk17n4M2BFQFwctSiYkDzTmgN5lDGd4Y2S8sUV/lxYE+cQdEdH
S6oAOagk8xCUCvSW186UDIzZTW2D1EeYkPRqebuqg9UBVxlTFtJK7eCeBzKclBBcRFjB0Tqz/25I
JzHAQvnLc/V44K7G1DlvNTkAE/sWD5ie4VaoDxSgoJyAfw3/boQ75TdhTL7t/ef+V+TOS5x+J1uL
+2Inld6KT3RQYlIm7KKrTru2jcStMq4WYGotMid54y/5Yb5yLrWf3r0CSk81U6wIMeR95xqthbZd
EW6yPyQJOzvmiVlzsb2jCpsCW6HPxN/vATKbQSu2DdhG+GQmn7QgZ21HH8RRfrdMQH5hZJISJElt
vagXukiICYTNOYqD2KmQBbCk1pqbEaxC/7F5Bb1Eyt0hS5O/MXedTuH3yqZbWlWkc/JCaCzIkmBk
6w0aJJlBqPKUUIASK+wgB2Ly1iHpVe9+Nm19P/GnF6i1kA3FhclsF4Y6y0gEOT14Z4Ma/s8gi7Ww
V+SdY/k/ImAmouUeGyD7YpJCWYtwZQg/rD7SJwMlgoaSsEdfMlvX6zmoMgLVcdOiD6ivNCnarJHE
msIs+1Sms79TktdnoxvdpLbMkbrQe/emc4Ga32cqZy27BN8l0GNwJhfJfCYsExathasPZlA0pTaw
KVMYm16R6LngFT9pwQ/M7rG/JgLuJ91DXIgMC6dGzhiXKCzLf/p1bB4KLQxml6fNUCEhrN89CvNz
BqshxyKY9d2iLgz1YpNfa7gWO36UKJauHImohraWubDfOP6YNeHhOTozmIZkkauT3v5qJJUFYl+T
lg3/K6rn7yNMYWY/YHXFmSoyjLIbIrIrQUnL6UpLo8mIUJf3jygbcuVcCZ25BeLvxAyyjdJqEcPY
rx9f5mm282+3xp/O8yX8DdmnDBla3TuUJlQYrZNiHzCtFkPaTyiJ9CCVv1G6NRp+tIEed6l5VvED
mAzH0CaBziG/4rqsJ/hNBB+T1T8TCdEFMouRlpKuDBqj5vqmv2VwSmdHOk3qziuP7uf/WEQUHmcI
+LY8scmjcyDt5lrz8AWnrmXzBDNIc001ba1aOXKntdzpbjzpxWy+18DHCZ8pmR0Oy2GTuW8zv92k
yu6+q3ZCKpPr52T3Hx4UyPdsk1RLIwJahn2TaWUKc3r8aISj3zwPBnHcU9k4B7yITABFrroLxkKt
EKVGvVlmZnlrm8c8fhX+EYM41hLVXF9Da7/QuVBOCk6BgQg+ypfQJFHcfuxh1bINxGJdweobv6s0
2EdM693i4IqX/pdhz32iCWHQ45BBTcPd6JQZhOSHPZ6ctCAhlGPa2fvdQdyi6+cFZyqMkt1anP99
zLkjapy0DkzPseOrmh9fy/N4aPIrzdcMSNuCaRx6Lwa3U1TTth+otTcOy9rrJmyk4wz9z84vjF1s
bobN5ca5YxRiAFDKWzuFjrXpX3dt4PzuZFah0tIvC6pvf6HpIx4zp6tBbRM398H/UZUBUweSxavr
XoCYn/p+ZsctcpESDPSSGapgi/JgxcmNVZ7mdr4YkZJNV28Il6q47GqjgP9Cr05yoyLPoUzf8twk
n8kW2s3IJlbsUEP1SpQgL/7HPFE4cBHA0WZOjH/Qvdbr7clCOEEJf+cfoaHRUe0PMK0BtgDI1PPO
yHFxjrcZnc8Qac8LgBr+LZTPeGakOkFCMZkHx5KMf5iqSx3EMehcDL08Qh2l3HimXO65JphoY4Os
EOO52aRVy0LHRm72+MSzplAEGzsLbejP/p9wkEbkNuBCwYZKEeRv21CQxG1DIk1nPr29ZMqnpg8f
bPGnrFuVQS90KEWRjkQDA1Kg+qcdAqCC85Ep04tH5PhkqvDczUZePlykeWD+ikPNQ+GbeUYJ964m
QLFVYZvr9eCy9Ms8vuLpbvNBetxbeOyc5D91byeFdlvJEwpSAR06QblcD0k87z4vvufLjpbdnwDw
GLDvbqvDYdIx0fPeFNOgCAwYI5QbKC9mvV37MzY7O59qb9CZ9Pk01pGOd7I/Z4wYJ4TwLrc9fqf+
LY91v1Aoa3VtBVeVpZ7LQ7l8JJKIN5whFOirer+Fwhdav/auPaSshQa69g+UUE9krbE8Rfmjjrca
3aBhQXCKrwhGDzaq9DiRMBKP/A1YTZuSVHASTs1qnc9P947kMUnaISlnJ6KQ/gNlsVl8UII9T+Pg
kaoUzZgYnzw8Q1w6vFvk/O6Agtp18Pld7nnqonPpSMJYgZ/RYJOfXRB5RMbdxMDgQ4XRzQiiLnlj
rVq8N9YLbOTLMuEw6mGNfuhauptPB15865EO+6lx0R+Clb9t/mvZ2aoHJbkL5T1u8DyAxL4/hZEB
O8JGmWym8gbWZjhBWmnuOics9y4/JPTwvd0lo0EUluGinbt/ZcJfJjN1OO42zsfLWhfRTCFezZ6H
d5AaufoD5NIYiK3VGRzABFSz4AjqZLrOjh2yUwQzYOZbURrUofAs7XC0o2FHKjvs9qk5wSl2Ksqi
dP/mOVWupMlH+PoO5z5EYyyHFDdAtGlwmIdcXPLwfiKuxHQkOWlEWKM9FdRNiWNWuCtFjwAq2VzJ
xms9L2LbH1P5U6jMZxaBniROM7p1Fdvg71mJkdK+lKPrztZ7dX/5CIjKyboPaJ9RVmzpeWBJQePr
XM0qoHyXxv1oMIME06nkaj7Jk4zoQYuLcmxa4G6XsAWO/vAYeLUT43y9N2xCKhCFZiTwVDJrTRWJ
2wVtW6sw5RwUWBYvZ13cm64Qgl/S+enBKhdqHGzuLYASmacDP0+eqzl/L54N/In1G3W7Boj1fFWQ
jZW+eGyygJ7spIECdw4PePI0mzUiJoWVI4tElBnaN7R8ivqSpDqhL7WT+vGPCl7+NTBXdG7nMSOd
YEiO3kJjmSGw38UByrYt3wjL2zj/Ud4VPXr3XrhRsFyr3dLimsgyjDNFbT9E3SRaln51He+e2xag
zSQSbR+coWosR0IiBZF2uU8fRUIaPSA1gX1CoNP42cuFsCGx2pmSBPONiryKLgv2re405wdDocIN
kEQ9MG8jR0+bVCmR8DGIaG9b8Nhg4Uzdjhqlplrz8LRU8IhId4sNM1MCwKqX6b5/sn9NeoLlQ6eC
znHo41uhw3li0th9zPKAHWWr41x3iBlUjRV7Tq08Ow+gnZGeUVLBAOXsdYKOE5YpZt5/8i35MXbY
mhnVQHuC5KlYgFwMvF5iu1zzv+PUnacNIw6Fnc25zi494rfrDIFyxocTLiAHIyImms5QuM+l99Kh
MV1eqZFHMokl7ZFzL683MIAD3qDx4o6i5Vr5XKB0VfylSjJChQ4jdDRqmqfthYACm+4gceKSlMz7
EwNemOQKh39O9K72cU2mmevVZ/hyG2Go9EwYi+NW5d2/u0d5DCVbL6ij744NZcdlgP6qcQCd+ZQJ
9jGbOGyB9az2Dt/c83VAczs5I3wE5bsFKSovGw9Sv0ZwFh8hMKk0cZ2Ph0gD/VyvGLxtJ3SeZm5V
uMkNGc6nnCSSQwsGilTM4dz+y7F6XCTTEbZCEZ+TRPQzlLOG1PVNstEMDongm2k5wh26dVLWmAfh
6Asmpy5vbc306XXaJ8phfq0t580qh/dJdEm7ixBALzrpTvO+G90tyUMOU0TRF7rzjfrBI5BnrxDD
VRqlmlBdDj9BMXpiYNPlpt7oJNKsbwVgc40CQuTDjYWqAEG8wlaJ+eD9tn0KnHY1oMLWYQ7DACWJ
waO0Ep//Y1ax32dBN9pOopnEurinidbcGElK5H/rKTbLKg17gqBulxsWMm2cQnnTurFsilV3KthT
LRe4+D/qXiBlUsGlaeqZXKJzVHtT1GKYa+oUZzchanL3ScriPuoPIlqcbqm5rjNWUQ85xIgvZ6y3
JYnHdgOCsdCVOGEwIMILaAjE6pmkEKoYGboba3T4hdkYFAFYtn1rN6MJi13GUkDVUlosOFg2Euf5
69jTeKbbEGsfQxuBR/IXpnY82ddAhcCeGxQ8wu6lAcoHjr26kJFG6Lxo0Ddai3qa9prJIJNCPhYB
Mt0bBGfws6WQ219L6cKkShmsgiPm3PkuOIMNb+earP+Iv6srZ90blheVXN5Pslf9rAHnwAwPWqDf
ZrDihK8V4vnP3CT9egnWmeda8f2gb5/vZhkKOen7dYI4FnAxvYwlSTVuHtXyXcU7M8rmyGLwjbaI
avf9vPmoR5ZccqZj7W+2GtLu4MoxZipzgdt8D4CSj3mYa4R8eGaUEcPaU1AyXcnmoMNxHeOJq1Q0
YgpTuT6FWyBvzRUIwA1Hba7e3IgbKMTB2QqV9A8k1/jAdYAiAilL8+dq29UslZFOx8CPifHriVqu
uj93KTzUB2qE3ZnwluffOM9h8lu02x0P6EB+cufZBmPKyr3Vjomj0MNyT1sTvm6vqOFfAWptswIU
vPaE/Kkw5beZq3E9UdsxWkrIS+c2WTzI6VgF12IR/5JKwfUjM/C1fmLI033TDLgL5VrR5t1raDu+
MhDA+ytJRnbC0gtSg9camVsA+atgPXhQyQC7DJKdnMTHhhCbkqaOZ+MOO29+/AHLw3sjHhH492Z5
WFMfEd/DEKA2b53pekeae9de4MwAJmHZlMog/xjzClm5SJ9vTH7PagwhZKjEnp7NdfVsj29EHSRV
FA2U0TAArixIze7q20eaI0pqo27NS5IrGunScK9Da5MR1339CiFOlYXJBzRHDMxHnDpNiNrz0oEs
uRPNXRXZ2+rOEQGnTnU99ggirMCobUa7kxAtrpYP+t2zxPvSvAy8xt+hXlc8a9VxH1WLX4uhay8W
7hx9kfRjs/nsFnB5zigOpUIv8/EbSqt9i2S7mzgEo5aKT63aDXrWOxArcxs6vxjRRvYs0L/BL+tO
BZrf8UP783IFy8axwI6iOY0j5jtDO3PB4lRS+Ui8AOz+aGan0ZwWpAalHDTfnqkyCv98bD7CxsFn
ZeafEwAGcNK40UXkguWPlhlgwHAgMoIHGpTjSklB+GVSYInfC1UPgKIcRJMj8PNFq894IwA3eENp
tMoI+Zrtxtjz/qOPVoQZ5l0sYl024PWHFcsIeIyre/RgeD4kFdfRJeOZTQMlmjiC4JooLuSslQAX
NND7VpswG3nNzjGqHz5LjDo9pjARpvHUZgtLviZF3Kiie3wRjmA5oM38RMJwFR58trJqLvgY3cK+
nmryDZ+FNnGGcmEpI3OQE2hfCJYAIv5Tm7PnpPAfaf8gPetVUWGMDZioZkFP4MI+rM97LQB7o+UZ
J4Y1GxIYfpkxCemYtGqibM79LNaqDkFIsT11JiOb7QWsuR4Ia5Of7tzJBtjicGlxakQbf7hbgm7E
hKs+Y0ofAmblQeLNaOX8pAkxGU/SJIhHw1DQABdq1xbMQyic/u3phvYKzpULpBKrR9g7vyQTeZA/
C5EgEmXoSYw0CuRpCxyXwvwVGFvVszLO46l4TLHbbCiC0HMoviKIwilf34IFyH8RRbys1OiR4Hqq
s9cB5wpC/n4TPlZ1bmrvmoOKnU+U6rM+i5B4EsvGYFYnW3P86VTypXlJVQHCDudG5gOIrnmtlZ0I
2Xqwj3ocjhTVmEdbCRuW95B6MeGirt8ISfsV1sj/ig7V+rNLgD2wz5z08p3Y6AZkmFGwNViMtbTl
4D1pLRENM3BnBlxGW9iewUWCyARIXqCzkLyaK62VK+U075kTAXUUbO1x/vzzhlvULz2X2gxmCBhU
zkARx3YuP98fj+bt6zcG0tE8750BGaoEMXfzBJdjpjlMCJMUJw1NLJlNKYNrHydGW8HKr3ndc/7g
t3VYgVgj5jvLP1/TVKyZdl6320yn/hJ8V5EHtnnZD1RAQlYrIC58piKJiLmGTqR3nQubXxJiUfqG
KNBaDQCVA/EN298DpLhqFN0TT06Xfk48eq32/CxN2+aaSGrdcoqiUTWthjnvQr0KmeyfFoFqa2Hq
v4d+rhuzTNFw96TteMMR42J+W7DXqJgAI4ZUBGgd706lzaIPfFUDrMX1SWCarqK+eplBcSInbrvV
kXIK7fKgk+9b85NO9eZ6om5FGJ6w98q2VOJ6O4BZANCIpmk8UGSmZ6z72nc03JrfbADkCFoykztq
9F+oM/AtU82z/6GEyEM6SQ+DMq01DT9UBb9OgtINrIfvBZpdA7kJA/MvJW+S9Ob4N8j+rr6hAkKW
hEwx/alnkliUwWl/bJYmBnL960QF3GnkespYz5hAe0vDQR8dflV0+B3OQyW80itZ5KxLGiVSRU8s
gSNrouu0QLHrdt5FpX+ASynrYSp0kUbR3X8FZ9yRqXKLVlYSSGcT1TxsCnDH73uHfrj28AOAFfKn
IBqULyHBZPfNjclXa63jVdavBcZcAmbNZ1k5d2McBHpKsIeaKeIh1imk9GnD3z0oyHulCO1o4f2F
X8OoIWCrg1qbPiD8WnxUCnkLKE3dCCfT8XE8RBz8NGNQrj6PN0893agYbaRMpjeBOGlrl8vSION6
VpaBpumtGnlfIcR2yjpsHcbMvMzHhWUjZ1nusKvnTz6AtxLghmDYlQoBdI3Z2QLhe06Gv8qVaYRT
+ekagjWW1gmGNq8bKwGI7mSlXvpp7/iA2ILgQOMV4sjG6ecNfTltzqaQwkYh0fODuq5a73wfusOc
iX0UMiFqOk8mu+eOfP8ek/kdr8Wt6BvApYRp/jOCthGUOdU9aJBXhDhnvoLxoylu8Ghb6nBMH3qZ
AdJBQQMhh6fWp6rgoqkQcDWkRBcPPm8kbgfPBa7vCzv499JR+LMgUKTW0sfA4dJRRNV1wCH+Sfsu
WQjafRiG79JiBUAaeYoNj6Ej2sp4jYMeancYCAD3c1dQWLUWZ0AwsVbhg3ViBElcQcWw7RrIXwI1
J7ZUCIkxuGV+G16yX4yE1sCjjsIPQLrQTbv7fwKGUzn0IU0AkrlTpX+yyjxtrp9ihhbfDsu7Mcwx
yure6nm0g3MJFvSmYDJnO9a6CUTszQFxw3YaX3Y4Z+T9YtUes8kQcuKwh/8F5q9PVNuAjqzRgQ+N
jAaI8onAzFnb/tQSNXXWaweX1DABPOYQw5hQNXW2kgmZoCIqVC+lzonzh/ZrPQ6ytljLaQLye5sd
UyHqyj1scFZyIFdcexzo8BJjjX73nNFrTIXG9gs9HjjaC+7GRWbS7wEa2MNo6HJbvT8BYVQdvP5P
sLYamPMl5Iv8Fux5uBySOCGIiSEyNa1gTjS0sFQLBxu3maU3FexBYwNwn44xqHOCH5gKbRoGpRnS
10/MrNp3XME/IoYlBWksJH0CGRI3wcdLSANOfd3fHrwM9qDVcQa/M31rAnQ5PoYFel5FiyvL5tR8
5cbVGbCwN1CTZIx1nmieEzGvBLldXsSSY3Xj9UWApwrqELoCf6L7oIuWnHm2iclGf1kCAIZ+Gb64
b0+dF6QcOvQGml3qcluFFOyoV0kPsfpAzxoQ5hPbeZ//sP1S8NjlAUcRjzMYAepyF17lVZqQ3cHP
rBCSKYNVdFxbvupjWpPCR4ydCoe+cEhsRhipx1IsJED7ZEYsKaDmuWQXlZPYPe4v6F6UYIV5K+ME
lhMn22nWszQZlBMwIki+fUMDge/tMUF3IymeYtzVjFHmPmpgwAGRKH6+Qi1pES/Jo2tZdZtGkBCA
KUYXDSViswip25jP133H4449SxHlHCUn28qS4X1qPC1fyLSjAH7gyTn10w21t6W50CpdX2Q/AT26
DNBHID93LlmGvQZFkQ5fc7dLCVgYNDExwCwZzdV4/1aFAZxFHlRL+OQtr2NyXLNtsuUp0/X5HyNY
2ciW4lagOlSjP/SwjjdSLqpEHAqXDhbbgGKlGfpo2Glr1nKQ3ErtBrDO6MgX+leJoyAmBqOAXkbG
1uz2DipuZ9UPsHyyr0x3x1+6wiunWowBYPh1D1esZ7g2TRu5X8eJbm2xPlArI1ApKs5sMj5Xwqry
azuStfG0dF2vYPqZzd0pfY388hfm4L0nthYXyiFJ+VBlYLI836OjYHzCWEjpJOHDatGs57s7m2Fq
Pdd/UAF54Mw0FF97h2l+h8BvMqnkplwc1jQyCSopNKDFvSC7PAEPnoD7Gr5SzKzbrQxelBbt5Hbc
3xxTRELb05mCtXonc7zaH2Ldje0BY2zaASPGG7oyKHtPjh7plswya1cLKaFjjK8AN1s9EQY2OLRD
88qw13bOhEH5s9SHp8xf7nnTNBzcj3F9zCaOjy9EEoqydrlyyCI+NVyXpbEqRD73yq7Bd/dDsVj9
ecbA0L2eNeqt6GOBpWkjBDlzL3M8vkSLz3gmhzlsG3gUDq1qA9iXTca+3CD9fVg0FJK+3+GA4T5O
batoIKAfvu5HKb6MQuEdCx7/vJdO7cOmt3mLptDcmrOdFJveBpSt4lfWAaSzswldv8IZm+bVdsDG
3kEqc/NYm7IAvj8KisYPJHJ08dS95v2QB3SWGOSAHrd+c+Di014M8P/TPCeVSb5xojqAHn9YoO8z
ccwmGnOkfZFI3ciduEwqgc53qBaEL0/FsUFi3CkNNTqXmq950gRFOtHXoRy6ShkuT0uQfNj6RW/E
Nkt9sJu60kDntdKgiaVcjumSkhpj5BDjh0YMhq1wK5l/5fg+3RQH4LJK9rMIgTVQ7itp/HbySqYd
6OMeCdmP7zYiIKdQS1Sy2jwqa0pQv3kmYwup3/82oUcvZnuJvptpwxdA5O6IC/1h+4ALvrh3oG2d
9Y16NETbbFziEY//ieSmSDp21D5T/bS/ZwDo+0J0bWJ/zU4gG2Muxn0S4SXj5YOaKlFyKBQM4hZx
jtOVqwlvCWin1Xq6kptOoruRSNz0P3nY3hD31OEjCbxFxGcjrZXCndlbhzPNTCpw/Ps7mpMLY+NK
x3QYkDk5qj1is3u8fZ5DYiTlEVs0SQNJCrPCvHNMv7B+CqFu8oC3JomJCEj32/Bnjl7A8Oa2VEz/
f0sre48b8gugfeT7U5E/tp9lkqjssOD7fKyCdjyn8l/KQY/8NHSuxjNWm87NSt5EC9HSZwPPqohO
A1u2i5bIALHeOAy9AsARmSFo9ZfPzCgOJjrRyKJ984oQuq3GyJEErbIKVA1UbrqHERdd+OrewYzn
ABYv7CxlIZEtP9E++6wjbxZTB77j734QsV3+H1dNPCUhXHW4wPoKVD/SjJzUmpRwR75Vv3ywzsNP
MMjqCLHChrBm5bHyp9rK7bt+g0SjOdcfUBG947ZkJJnjWxeqN4xzFgEo3OAMnW6ZPkWMZNsum8+l
fI3v2VxhcQTlApzXCvTHMZTdMsoDscluhO719+X2TKLiPfNxMY8wao9YKuzE/ShMJsaknlcHGn3j
yvI1g0MxZxfnHVapPaEWh5JQrbHWZvpNmJEzrc5+1tEZ6MirgYcS3jjqUCWKgFDemGiy9xeL4bAJ
EBYK7I9tK9v11MGndlrfqDdvJAKVz8FVi+IT1AjVzYFc9gb/bnJN/GF8w8Q9iVkC1jHlH5PQo2Gd
M9LUU4sgmxR7BF8l4ixvRr9FKO6GzE3vZeS7azPgxLed51SQmKjzwkObRyl16HnG90L/F8u06vRP
pY4qHMv4XDRaK2jGQPSns/t13EthbKSpPcsD/kVRRxPAVCyLmrIiS0CxmNeZEkblmCpWLGTY+SDo
kVTbWl2fRAYt8w5Y0x8fWJgohvZe91bW8SeOspBreqZ36/YfmUCSV7ifsK+j2w2WOSyv6U6ElfxY
eFIhnkvL/+XJz+s+h1N1ILAEwv3t2mGMqn1gTBErzZ+fW8130LmqtDFISagzd70+pFNMTIPwvB8N
yU3umrrmZFj35M/RaolfQgU3nip8zmzpLrf9Duauh5c6biutDvebSpeRS6Q6Q/R17kgWnBD67e1E
j3OK60NrulNqTP14PRyAWEL217P8HnbgNIn+Dit3JcAOM+6GB5QUR1GLOTRno7YNohbqnQNp07D8
uFfd8bgALCg9bh1DeZwxJ1jgPVPYm5CTZwXgsR9XxvBr9TIrtLNk6YJLu/8P9slv/4KMAziU6r7i
BaJTpv2Wgh+qiMhlRdCvw4qONJ8J2CiAasK1twPfqQxcHQcmNxLBtIn//wrRlBTaB0bPNNlTLRmn
jVyevqi/02ftN45XXfSfqfZ4mRyUL288KqYJMqwaNdO2VR16aeZOciywoB63xZnbVEsgpVpKEUON
af9UXMekCx1duEYkT6/pRKVxmgzttSNihcj7SD/Cbj1fHApD16PWjYIMcY/QCQ4esi/Vzyz2GUos
sRY2z000UULz2GuSIBCC6xdegGnHVLN4jPJ9alOH84FBzNZokXtxCsSo7ceS9OXQySjs8E8S4FwH
qXClMmGPhNuYKbZp1k1q56y/a0nhjDildo+fT2RWWPmjKkQfsF4BzG85AG7pI1Fq67iPxM1Kh7PN
GiblqQg8pdxe9uViG4s+/wMs1aFLi7kaDf+p7+UZPYX/WLbmUv11ggO9hM9tCr+rsj55ExN5+H3K
Jqo00u+iit6eZsSSTn+kw86po0q2NaTWY17/c7IDYi6s85GGoaNbYnJTnSWPG17EUStEkZ7Xxss0
chf0G6MBR3z418HWq+N2UuDqcBKOo7F1fjjcxrrWcMt3PI+1NJSupgFCJUTb/Sy0t8r5mPcNizPm
iT5oCEah2KgQCenNIbDhfqenDrLj8XB41k2BXShF8L4RuYMiglIEJjRdk1/5/DpFTrVzunHIhJdK
8O+nsCQTubvSv1Y43ZwGr9vEqZ7VhCDnBHPOR7p0rWg9dkhYWbeM8gKUWE8wzVGeXAVdWlmfeiXZ
w0FdwcfwMlEonhoXBvugr5lw/InPztjG16eKVrI/UHpelElJyKPSxlTnqklx/Aqx8HHAvsjZ0pyX
pfrpPXWNM3vNqpNANgmMb0dFN93grLxlMhmgH3NI0RtiwAC9SDbHT2WCNrDjDmONW2yVUXiP76Pj
iTroUDcRzYxB8LB17jZV0zAhNC/oX/Hmo356GY9vfJvstNqvgDw7fVGafNBNIj1m0QV9H3KwBFMX
Aq0hunVE6Y3JF9zw01lcIhCXlCBvafSru/wEc0/Vj7/XMYV+h7CBK4J/zs9kdd4CGdNvgSVR2VMv
lBrZDnBEXXdxqsiMr92chNagyjB3W7ddW6JYvrChOTFhZhFVOkHW4G1CpLHHhSSmfwLx2wSqRgwL
xAGQXkbYwz94oYxgDTEMUXmwvic6lAsPSQ/F3tLqMHr3JRU00l5sCExruWCSyAOfNuS7Ssoy0RVP
FjM84d8Q1hkbOFYSgGdSW81QXVF0iRDWt23jmYGbVhbZhR0VltBkaft3Ct5c3khxLGp5PotbIHJq
Ozsw8KZQLibYU2OwcnCp/xgO4YvkXT7CUF7FdP4KjgVWSbAvxXAciXG7zZJy6VH3arnHhfu8SlUm
0lUYG4AcY7MXKe4tcVu6ODReyGR31fW8/FOiInJOBcGyvW5Q6MIsFb7jUz3JP33Yz4hmk5o7KDnt
1C2joqQbLccil4gStW5eWNY3OinKMk4mEsJjQbPaEq7a9fYKgUDtfuoEQVwHFOMgSnsyYAKAFRJ6
PdVeJ7ER3K7ctjV3/BpZ0My3P/W/MG2jaGtkqHSgZLykdP58tLdtbOxJNtua8fU8ZM6fErJ8W+ok
nNy8ig5qmhe0Cx21mU8EvB3UaEgmUJrAx7XmXXLChqX5/dJUKxRojIfzbF5lrxUBKt7x+MMX+/Fg
RpZgutWtuJpTbCPz04LF7CreAv8Lt4+0vRIcphrwUAsZ6xiM2KT7Jpg1q6HY2C4efTBjFeCMQRxs
ru/X3oL5pNdh77AjLEqfdnIyfaDt3WZJnsqjKfvN9PRqRQ1ZRKQCeCu05CG38QXGBrqjIlpornlC
jKD3VDW5VEPYvqWA2bU/3dGZZ0tM2blMrJ9prJ9cdXamkKJQVYL4wLhgEyTOv6YdxRFL/hYQ50Fe
vJwlkjc076o3rBi1VddS8qe9kGWobdDaML190f3ssSNqrAoO92ydsLS5yYzZP7vRMuptWLp/AIzw
nKVqhSQlSDJ8oGXLYvughTVAPu8gJESX9WtYZBZBservMv9eq6tZotvXODiCbyzIijgjHiOzKAQi
KfSyz0Yu2a7wmjuY3XG7QKHohs435k8DHNLG9wcaU5KA/VrUW4MYw13t44EGU1i1BPtqjP+v0cnS
mkuMjT8W4IytQPkFCR/oYaVCDsJ8GLHo6NQaf/owMS+mvfXuhDRHc4MmUITul2g/G7ryCYzSWl6N
T/cNQVDSrwdFnv6k4ZDOvDd5ZYFEqdl022CFsElbxIR6qRXcPV4Uc/8pfr9DKsOvMhvZRkobUXdC
iVEE8vBA1fxboLyCuzT3b6uNZYP1ELI+ODY2i3W3CfuwxYyvhkYw1D5PT7PgTgDqtLXcRlop4vZG
lg74deD14Vs61TTn0SSzML3zv0BhC5QdCSyrUuQZ0iWLvuLimHUI9kCyC+yris/lbGhMZKeiekeJ
vgxL+HrGhBRaoraDxOedu2SeiGbGqi8wp2DfkQ9KKrFI/3rpIBdcr7HkIjWJdeAiRE/BnMKYJmpn
YZWUwM4sgqBclws9lFxN3Zt2Mu2PGFbqQegfOksGm12Z0628yqPdyKnnhu4+I2dWBH7+4aaTndgR
rmZF8KD+fLoqOkxazk54wyjMVvnDc1W1zOuMdH8bvHq1lxlmvRLHKZGkh1ItUoYqvsW9kjfo4tBc
nIB79pc1E6SURxbzfRwZlHx1JP49ZfKdfOoxEKN4Gn173ZNgtvlnO4F7SNGqyBES+J58qJR1gVJg
olgbskg4pFdAK8BBgdC5OIqUyUWOMpMdx+0mT5TNgpVlnIV+mh074yzVj6tU6TYd9O+kE70SOGEw
FgY5uYBeCNrKXJbn7U2LUs/WwKDLbJZTSj+d4SXnvAkghk90D3mtM38Mvqz8kdbEPh+x8+FEbhWz
vQ2RXWIcNMrTdWELlrti4Y2u/3WkX1H9gVZN0GGmeOq9NoUp8dRHhURdTr3ISHy4/PPCCWnTjVk7
/cIEQ0J3K6mxt+9/mVjoV5PPza6ykRVagSFpOpncQwAU9bAzNi0NsGpL6I3pNcIG5xJWPzrQhvn7
drFTSJYGuGLzTRWE+7Mn/EWljWf+5/PtpCMkZeOSnagZ98KWiiLgWb7AsHv4My5ZtidTppzf//Ww
gP3KUkXLaj/QPU0yQIA4iw/K5cYzEG1r1L88g20xjw570zTfTFo8F5WNm9HXIPwTWUAdpjgKsqXj
nhA3nSNdnyh+7hkcO51idIJAv2CFhChHTjuFnNshJHBTOdUe8ze9fmkWpCfEIwBU7rZzo0mBzQqi
pRBA+kc+jC6Yq4KtVgvDsYYBvyVNs4Qg6NB3JWO/u8vMFbbI/K/jRk+fRZr2FQtJMrbR90IKHa7V
2S+GXTBxf6omdwsLR0gkZpYLss4FXhgvh7NS/KoHQRQ5PCbTT2ixf8NQ+bJ0X2Y5gzxqKdMvBGY8
/eanfk1RvCzboEWW/FXTfp0459WmLJ3gnbE7V7EZzosNAT50s3Ng7VFKqlx2Hb/dEGBXA+cZVRWy
YsM7ShWoSEJ5YW9zn+RK4zKHKB6DNI99gi8ATO/KFDMNuV5J56w9frdp0ZG5LRYLm50u5RdDXoXs
liyBHUbWreL/6x0wbRhnfW+6E4Uq5FIc1PiTIlSOaXk0EbfTYP+PLNZr+cCrCnet5xModHInI0YF
ZBgVZuErOtqnGBlu943j8Ql4WWd/ZFLj2rX464hHonUIuKypT+8AKmj03IqMBDXM72k+n4J8cPsd
B9VFj2tnFM2jye0asJr+3UwExv2RJ3ox6Oxg3PNWA7Lmjp4QoFCoylphamRUplLAIU+q/JX/XZK9
grRLqjEeAbiTPKJEeqxkMNe1ajwmNjQPuEjnqAWl9sJM9P904gUg3oP8Huclziap569erMUAr8DA
ewnnbhdnBWZo31FPHM3+Cfu/rBc+4no32Z7zfFDazwMl4UMPl5e9dezT82O8Kw7ueV2rMVuU+inR
GiTfsn5Ce3v01T1lfQENMIfZaalZtIuJvOV9i3DOa8jvlIQaZqxhS1wDcLTd+QLW8yU3j8jMSizi
YMzSdFzP4MBFrjS0zHenklvDUWX1qWNGI/Oo6uhgLjM94a+dEmFX1cY56ED+ylDNUEUR9nQmjyDC
X1380n4E9ATs4aBCp4OHIhbS6CJKCGUaNxsi6faOf3MXJSYahLtSZagSvycUb8Sm9pd1yVukFeiX
SgDR3y3L5d2eEbuJf2O0lwiy+MitoEhIJA+buzdiYu5/oSIar+QVjbxYbD39MlFKyBJHwOXep6LY
cHTX5vDukMHjfH38SNNJFtbusOUAF+H9mPXRrvtBA7UMg4kS8n/qcggFydgyAr7vnuzN6U9IDdM1
vbGxB2t5ZbjXNkT3FiamJ0SYBh+cAfwjQfcDCsuLOZcwtJXMQjXiC8KxySfKGB5OT6SyxoAYhSxw
lX2HEyOobh/75q+Y4DwigkdxZMGdp7D1lksSIUCWmSBC81i8Dyr8nUObKRrUIvbODbftvTxuKiip
0ceznS4IY6wLGnJra6ZaOwitOR8P77X9ARvd66wI2h4QEV4hirl1ldqntjmcyMLah69ac/uyMjBy
WMb5Edx8NcbTIKuajuibCSzjs6KAhdcVQQ9GHhwGQvvYJRc1/moYBnX2kSp5YDkKDzSFCLwhCSfh
TwNQ1ikUeaJ9PVKplc1OCCvfa34+Y3388+O6VXgiAhR6WU3+fAc5WrW8MTDMgN/atvQ2vgot7bK5
UyKEiDvYoKV1aYPwttGBzkaOGruj6rberOafrdYEfrqdybLAr9UaAyouvbuTIJFhyP5RU+Yi9g8A
mKqtFwckQqMH9pYVZApN7sujK9oZQTbjsNGP1DZWwQqJGHbeaaG3VgP6bqw/ol5EdgoHO+An6HJX
t1F0ozCFJmGKrgaMFHa3w/PUxbFlqwSTMgJQGq19FHhYOyvd9v3KSUBMSSvsboxkBKEwv+1IsALu
QUED2kk4r4+lMaT9HAxpmWiAy9IGHADMOTxdka1ht4dCsSxTTfWpUVZMsrUkIEClbjJ9zPUAgz57
F670jsboKjmP3AMHpCOD196zcx9KdnTibVStrSfa3BjXAabJHWg421qzgpIxZGZ52NlhZqocm0bS
Dw5lFFTh79GE1NyCanIskhZP4O7WBj+sc0dT7DW43XUsJztPKg1CAy9Fo5bRo5eZH8xWV/YtBp25
MDA10xzW5URKK19c6eNPDl+hl6jrcbcF0V9MUHKHMUCbPKOXKPfzjwWRYyHNQswc7itT9/2/JfOM
62RoktiHGKrShpGdz/8JtV9Zn/E+RdzjvXGF/6tKQF5m+rcPLCTn6TasraH45KU9QLuoFcBa6Qn4
/Ep6xfv08XbUMmYhDTMxHDeW5bEZvGnye1x7zVWwHZlcU/RK/uR5lYe/uJs0aTddrKcuDgLGtlDg
5sZe/UiLU+DfeYIg2YUKFzkaVI32T+Vto5uyus6Yp3RJStyfTkC7XSX1qJGPu1OOA/Qo3VYnfVxD
36LzzsYUG+07jX8T2XZgYY1F3R77Ad2ZRk5idChjWqmNqJqBS4UC6AWJsBomU7dAjBPV6t4fK00J
b/UTm0StzqmYM/kKWLJY2idoEYNKlvXLOG/e+2tN04rTW35zCJ9QWUYT9QFVBfrE5AQCQBldvhSi
AKkcZJH+94o5izeqTMIY8eVS+TrYmVbzVab7hsAXRG9XtFmyJ23F0Uw4HwdNV2ED6I0xVRSKQp7J
3QgapSmEDBoy2c+1fzeu1ut+AdGZkjQsu9cSfrUjNvu8qK6YSHhrabc+BImvaTupP1EvrguOrikN
HkU96J4Ujjr0N+ZHMQkMUbjZA3FvzbR+3Gh+Y9mJ7HRlCY/SESMNcGAEaPToj4g4KpL+gUGWeHYq
SgoeDz7MZEwQLxKHNnJHLufBRusFBe/u8oqAEbLu6RKCCnql1xWVlneAPOWzkZVf6dZHsx4swa2E
v0qmq4aHXRhd/HDGgEZebDYASnlxCh4ufI2JMqFZKbcg38AmzZMbpkWNfNWrO4M2IGCCyuc2LnAP
0JMPeqi8KandjmXeuPz7xsp5l/rwuO+1JKyQzQJNWF+kOGvLgObpADPMqUbrvT5+/egFyfnYtJ6a
7mWtNzXgr1Xia/uB6s7eVHrPjFo2C8R5Rjft0yV6xnI7dIoXrRdp9mMMrFcfu7kuot/BU27hYJ/j
6rd3VoBwlkXObl6+gz5oYgfD1O4YMsWyWFh5vwmMpzb0GpD550n8ZG8tYvWOfn3fcjdZ4ClXXuck
cxwGjTBiUK6CJ+U3U0HoJVhyl4gwyQTM3Hz3djNBS1vFJwAUr/YXmivWlYG1iwYfggWW6awh7p8E
1biIiq/FeR6SZ4Ug1L6Wyfh6vNVpETM1sRRJa48M0XZqoiBfxqoDLym/c3JdArA7L9Xg66P//njj
byADXANO7XIvastTV8rqr/s1QKDzalbVs28sffIGLwdnKRDzvhvJ5FvboUcpj+Gnt9xp6EDY9sqK
RiAVuZFG5xr7WVy9/moCYdwzsVsgTpWA7mWDCqmlAqtow/HTmt6+uP825/RySbRKZAnMSMslaoZT
Crx3EBQQoIQB2VnnjCI9QtfWSdkkw59lHroEatRl7aoebBFzWS+AU5Y8WcX+8qt8YqtWMD9L8nla
C5FU+TmB9kg2ieqkdq5QWJ0jnn0/wzt/0kaRieoGmOSsa1iUK5mm35+XuXvmfgufX/76JrjkvDNS
ZuwJIm6VieXOw7w9Sk2GNyGWM2arfqLdXInsqFefmZ6CBZplowLWqv94JCpDCbqJ7yfoApsuYRra
we5OEsLslICmb23BLoRWiuE8zRlsVad3UkLgtKOi2/picF5SktQlfU31lJmwgI8clvNtbO6Ssn9q
OQ4KGFo6J7JLEGHU/JSM/r3jgubp+tJCE5WLABycTLnrp1DEgyjRaPdZc+zPjZXdZSnJ81DZEe6M
iNClqYAJx7YKKHAc0Gz8YVPpEz6R+pOorUIr34/3u7mI2wD7gpnfvm7Hz7Ed0a7kC/WbtpvRYqa9
BH2f7loWlOZLrMTVClVATNelYNPUHWkDl7HU7VLx1/vA3vFj3f+phUsbjWP1hx2W1SGKfXoXg/q8
AI6R/+DAeHlkXNl637ppL13xK2owZaKYik2GsOEqVd0CJE4cW84L453pr1fjULCVdDEh+QREHPdl
wH+dK5SidMuPPMXaTE2WFvqT2NBvExRVGO7XuVi8EWL3NIOhZiZOXAm9MPHoi7wU2hUZh0BpDeWo
v2xi5yjeMSNO8kjrNbA3e9AUoC5gQb8vU3Eb9tO0WVgqbpz/xZG3hYh7tklB6pmv/1AQGeOWxhNW
IEovlsgad5QEE8NLjQjmKhCgpj1tvNSSkKUm4MjLDItLBetFsIUAbif0keJSf5HAb0RFuu7V6ZLS
2WXs8ESCAGFDajLoG1vmhuT3+Qkhtx0NdekkdMpFXCTNbq3O1PhcXzvSGVIw0vezKOGHW7Dcc6Mx
kkS+1FpQBVUjoddT4FiV2ufGrE7XpyQ2ipIPofI5WfIpFXJFJBS1AuqCdJyGXFsT7qyLH02HxRpx
Z1fUIBiwAq1ucCVk/9z4A4pYAAZG8HEJJIzT/ge9eS2Mtoad1h2ZKk18D4S/+oQXsjD4meng61hI
E5ZJ7IuVihz1FEdXlruJS6mhoQ8YF0JrvS0GaMbTBaXY0w0EJU04PJ78nQb/hpeZm8D3QZIzni2M
pA2twZ3kgFoWXm0pIAppFQfiLQnknUGngBVmqK1vMmkqO0RW5RXZCtj2RzPRpq88WRKtvRKSBO6q
owy6vU9QMQoNKosOC4DQO0jCa9VXRst3wCKdGxiiPE5QDyyAuSbHNy2Btsc7xm6BFDJe1E6LDpwg
QsqadQ1ZjLqI+N+fPs0JPcfYDHpjLrVmpWUreLjn8ojBLPbwwdsEsBM2crS6BGj5FtUKMXYA5WfT
QtCpp6bMQbU2V+6pGwoJEULleHVwg2aEDPmeBiiVHR61OkQmHcLfWXtGyk/rzeL1cDM8sAiRop/0
S6JRwSc36cRZib3DyQtOUWkFkewAC9wVNqWwTciULwVcFyi17nsmGM4Aux7pWsDCcsl2MJ/5Tx95
gIey4WT43CQGN8a33zUSsFR56UKCV+lc5kZDs/WuUFeeaps1kPb5WeHC2WbffXR69Tx1bJGh/nab
FMXqsxI6jOniHOU8JlfhRLa96GI+hfNLS25KRASPcGr38i3iaNXPJLTVh5mTtsHV9t48PoQbdi1L
dtc92egkDDWcE7FczioTp4BzBs4Jz/tgOJ7KqSNrtunb2L5VDGFkgtLG2V7CW3oPEhE+Xa0mfW16
Wnhrbkzz5xtiJgcg2dhXP7LHTEjJK0nTbIKnqvNp6rfhPTFf/jNe/nOyjJwQ2caJg53tOoQ+ZNlk
DYnqVD0dq+VvlnLS3Uf8EeKk/oeYIaMy1c4AvCi2c8kJ1lD3/1lC6BzlNo1MgiGiAYXYLAwkKlUU
PKCDqr7NuIUtZYTPoWtkINFexRbiuhwbRGUbmJ49fa5hQXLbBS/hQzvIU/4CS9pTw5fi+rBwxGky
/GYaVW7CP5z5Lmoh6zZI0WOiGKZgAzm/ATON/qWhV+iczqkUt0r44TFQVmTx3rhI4bYs8fRgRGak
V04nGLQ1BWGHdL89sVjBxLP8oxbsm8ASq2yDjBOM7EOvowE4Aw+BnkIWLH6owvT8crCsz+jRL64K
+7mPELERrIrrznfwKJLWIi9KYdbHJ6y7LUGJdtoytuPnfRaMHIFUelhlyNDZ9qXWg82g99i/7l0T
4sdlPjxOep+cYirFCZ0DeMauFPO7OmSxtPzoiONEm/orWuCDB7eErpys/nqK19jiU5CBHmvUf7KR
Us7JPlWuKUPfabQ9UrOBnLPxWkUrOGVMYUOcU+7JcGRunJyimj5ALksl3YoNv+yHwVsFIQaMNVK9
WyIKlwT7XtBp8q/HmFLBtQdTlrkno0mjplEFJYrcNRAtCq4ThjyVwxZVDOUYI5gDg7pejYokRxVz
iezLOljK0Tl7aq1TP2DhBxbkMrFNU7jh3+xKiQG1i2IaI6ezLvtSC9kWYo45DQ6ZKnTA9EHvcedv
HuBS3g5O6t09HpweQ+Nv9Vy7GDfXnMg6KWXFtyBuUn/3jIhNYrqlSPJVJ9bihtcqxZHPF/TeJVgW
dTwvQWaIUZfxgviBKuByS9eVFP8dqQFHXVQnrMDxyq2s2Ro5Fvemhe/NJ3+yfd5Q/JoZpAcSzOLW
q01K5sueepCFhZAOBK2hmzOyJwoTe5+pcca4LN3E9Tkgo+2idJ260LKf+oQY8P7a8gotYvR0haKd
n8a52H5KcwVctZ+AiSyeoKjUK264E1gLKU6uMhYNERdLd4p8O/Hi4dyvaJuh4CAP0nSgH48XlU2t
2x7423nmXx7t972muvtQFeI6V8x0jOniQbuuhFh61JfmvCCyZKCtIv7oQftJG6gDFd/TwBfNeNrV
LI0nRuQFR+Hq05R/Yu6Ql9J/YOODisZfvEW3xFk5pJ3cjjdWRoZAg6I8KgBTICuAm3Bx0snm7vuO
MlCdWGJBZ+PE/CW07hWqnqvHh7p2dB92Os7rakD1Mm7f0BEQD0QJkEm0T/YUwSktdB4JbOpoq2sO
9sQKrax6zOuKmQmZtY5PkHJj4ohnc91jX65l9yaFWiOuQYbIoG4o+0Oldbt6fNuuQ68EjhbLuQif
k5Lmwx7ZOm2yhD5Pkt+Qga30BIRMdlLwVN+TCE9qESSWKb135Tgr6OcBOo3WDO6pAmkJjs1G9Ks8
hCpkSdu6ijClO0FUZqzlW3r/kR+z73uFdwUL+MySi3iwbrtS8v2iw3km4dAtpe2LmzsA3cMYOu3L
94uVxR1EssNjI/jryN3T/PABl70dNacKKTiFSHp/ZbEJ41lX2KN/Y6ZuaGHYmvjFPuyriVSYWMwM
22GMoAVMDCzxlb9dAKIon92kjYNM4ZNfAKwjPcCHbnJE3zlJRJ4lOllTl6iI/tbhTDqhtilAwvJW
x3uIfcYNaj5szsq1iJtfTVD6aovPnvCC5mn4BKWMxoD3bm3OhBI7DZ+hC4YoF6vRXuL0GLaY2IQS
p92vOQhKndwbVtuAhBTvQZQpEITL/KBzyMWXBhAkJFMpR2sq7TCrwYCzMQRUWJlNV7SmlY8mf1Wl
VBJhwNQdC6AMN9Oi5iDBxDXNU3htzs3G6nHY7SORGEqvqmQn9tnMh+CGJSJzI+RCt0V7pPfzbOG0
YqbFRjx4m233LkRZQwHz7LjCBqo85p0AJLsSc1/XA1lsD9xKrruluPJav5BIh9R/fLQ7afDIEkWs
oEV2Lv7F9yigLShaTNnNu4S5Ew1GMrETkgKABMUMUlC4NLb9TB+dcwtTZ5s/dwIIaXxjlNKULRcT
K1l6nu/384LZPSjaoauUmDriErnaFYEwBthZS2/k5UABDa3hqilEAOtTfrAj+SVpBHGoxftKY6hA
kt5lnLvX/K18my0WoTemg40bhgaWNnLLWWU7/1dxLHTqgkPzYVusqQJtkUip+8ALW37lu0bTbI0q
2fn7Oz+oY7Ju56qczrjSEuDGfkroU693lSyP5osrldEhHdjTJO38mD64jhucms0HUQxkjlVT/kG9
pD+Ra9b6P5MP/r8EnV7Lyb1Y44S0k42KufQpNCpmmnrC5is4jWUnIR9HV3llg16dLDXax+cZLHvz
kQS0Y4YC+bvhCwRXai9N/u4YSKVlWHZxarjiTDxpUdkYhmaG+NnBkOY5PFIJbIv3qEtDOw7IfBQd
5PNvXf6tptk+TKyiFMPflRUjqnqQ4D8CuYiBf1FECmOQDxtNtWDcFPzF1TDzKSRjVlcAJcXONitl
Kf/8berbYMJXNu3Yxl/57jwb3h3DYcbMkZu8J6v1r+JE8phQHWE7LmXenKr4sAL76cuQVH3gs+ON
HaLlhQLKf5vi0DskbGOSmkHCBGAJMpSDA9sfVGpVyQZiI1F37Ku9Bl72c0/BlJ8QZtt700a5RL/c
VMmrgJVdkQ6MqmatRPBEVbJ+xNwDCenUobKkgw0o0nxR/5vT4jHfKMOrcNMKUVdjSgO4emwZ4PCF
0lh11vGLV6b1BQjjLzkMqBvavxwI3c5SIJVlD2OCUphsVJKYFeRjotSXVlU5IWrpjYmjq6O/89H4
7WGG8t7rdYFWAA/xyvC3/bDIlYrdH60ijuaXoe2qadewFxMk5HYWo8MlamceW8qUmDRbAYwxHIAc
mn/+RmZJ4s1mMl4I3b73Ots5cYP+mgipfAj17Qhf0RAj0Uwrul412DF10sGcMecJeseWe7MJW2kC
pZctNrkbIv0Em8GV+t1v/cC37J9lkkv05nHSxU3Lt89S3soVtUlDmv0qQDR7+IN1Iy8ot/weSBU0
SsJurddAAFRcxuLqo9BrXsDaIjczn7zqJqeQgyx9/AcaARgGUDaWJyTTWho+g3T89b25zzbWqgmS
QhY4bZhnyiKMb4ZVLSgCzkd+P5SWJTA5GX9/9c6R3bRjG1ngtK0Xs1kMBkfPKAkb+GA942j9pcUm
vGRcu68X8Ash9OXsvWcssJgojd4eKDnnC03AGuvn52imkl+K69yCJATDt2XUDfHHD5xA21hhX85P
liEvDMx2uyupIilWjvKuhcy7XYLvA89TcKLi3JTsGA+Crdao7gRQ9a/Sw1K54LfROPtQDOzMeUw7
q3dM39R++6EpP2CZT9YrKOheo4mBwqjYLboQti5m+ZMeKbA2PMsmoydF9Dgtrj707YbRfhdHsMn5
PMtL8lEbo4BRCkKaPqf9jkMMY0QfIP65YR/ctjO9ie2UdlgYDOTIFYlHDw4k3J2WPvvm7So3lwlz
7JR6oLtRTPLPv4Mpz1pmej3N5TXmxcVkd6ynzCEhy6hcipSQOniAsGC2mRrZyn/Obwjw2eB+DYd4
3TVCimPYxNlqfXHhgSRqUJcNIW8V0EW9MEx8KMXue87Cu/BfunW3IOKLdE98k+eP/83b/+oFMxYQ
WWXCwvroxZRdIHZYJ2LJXHd9r9+hfilcSTxEk0q673V6JzQPkyIOQ3SiSG2tEfNld2B6cKdNyp3a
5MWXSjGOj2e89TKSAfR8oWfFbwI+94rJIL0XEVbSQLUMbl1aBgbiK8N8bZ8TTJuVXgumxPGDfU9N
ad/ggrMiFGghrcOQqlvsSB2wm3oLFZ3uGlfdQLRHxg/zwEP5VnDLIXhYjSYIlteq4s7qKS7w8odZ
QyR9sNIBRjitipeRynIDpxchu5zoRkuGFCiP1R9oteafzAU5LX9yr09r1ByhYzWamVOfGJLKNSdV
A1JnpFEyWhyWetO57lUQAKlnWCU/M3XuSFX0wx03LG8USSM5/ZCDcsb3TYNCdFWPKuenFwiO7MEH
iXZaFqn18kSJ1+IuiO1JmNdArtRfidju8l9GiWYawd/E/VUkmKa166HJBtkWTnAAEvJLFwmsZd4s
/UFma8M3TLh+2+1gzuR6dqbCFwgohAcVY3OhqploixX54V/ogp4EEKRaWetfluVu1SCVu5pvKRLh
IZHlER/5VFEVyyLWdtzW4G8Pv+m59SjErBzuB8D6wq/603moZc0IhrgBxFFDN+40LDUgqZJl+U9q
A+fWu794H217eDILiyoAYO+sQVuaXBPuYFWuWeT+iy0xYPH1Ie26JWdqkypVCC8GtUekAGCWwMcl
FhZL5KyV5kwcPZWoz6GodJ0KRJyZMA7r3cugIBfwMCtEehKwPxs1vWH+lVP5YpFsCS3RDn71a5ku
gyDHP1PW+eDmZO+XDauJz6L0shfhZ8gFBuEf0Kk0T25Sr09q9p8/iDq+Mg90PTJvRelHMTgmaYPv
FaY1Xe6yil+b2FF1wP/92ELc/YWs0YrC6VvgIDQ85jJ8Si7lNMzxZ1CwVMx2jEpeQ2/SVtBDjFRU
zZpPQA4WP46pkP/l590+s6rd/iSZ6CX7kBoVnJfnB/dBloVg8Q/q/KEm/Y/X5D+jRbsegR850U5Z
m1vbUvBlM7rRrmvPBjaYMfDZh/J4ED84yPgsVicHKpS817i3v1ezkzvr90VXIUKW2MuRe31aszdG
GOhKcZhABv+1ar4ULKYdtXK6F7Tk9HJ5vKgkLcmi0t5HNBLk4r1QnMhlm5sowWXNdzOXEjiFp5Fe
zvZs7xuexsZd1B/XvrXNUEB+8RMepcG29cw1QlIuYaEssd/jrW84h9A8roCLme1sdKu6ixB9TJtB
QIhvCmr/jLwk9cw0GU+EO/TAEbv3ytWhRmkkWGvks9lMG3RKUVDlusA+o9Uy1OUTux6Ey2FWwbPe
PFwbWjFMzRVIVH444b/F0RfAxlz5tZXjZtjh8hq63kBo4xnOzxuIQYDx6bsaQIJzsGPnBxS1pyFu
8dHzM5HKkXISCYqtk+osT7YYpqj4h0U2zPQ6hXVivFQStUmuYyRoqRBZkfp/6vQTsoHQ7QtWC21N
zYDSmohkC/Fg9mwP6NiQsB1LmK0UgsUDDwgmJgs6akukF8IgjxI9sEwb9QIMvQ037yCxhLMl3Vcn
PWmqR44DBG6oVBxreGhc8CE6K9a52+BWIux9ih1iV6aZ72OOnQJSzIUvz9iwMpza/vwOccMRM3YG
inaAyCUJ5LS3gdem34uPeoYeS6l96k8PqQ1KYBPaTPU+EWY1IvGM02fre+DV1sXAggJEie1r+o2V
JNmsvZ1xBq10zlFeFli8rjXz4Vqwc7GsMNYRkCqcBGS+2ZzDbhm5/A0tNNRCpZHDWYZmwcyjPtU8
YuMOoM2f9ecTYzo+4/6JfDtb8VES/YVem8UQDnMDxLMlL5smX5+t/+iEOW5PBqn3BjTMonaoQLU3
Wa3+AuysxXv1DyrpjsaVttu28/7NnlQNW+UWw4IG3A4oqxi99F7P0Yhxo39OGflkqaWIaPwHQuHg
uEUCCxrQrInYDzIDEQFb3lUKpY16uGBKnjwem83OH49hxkY9eg49QO4H7tJh1X3yebEbprUziwEl
1MQJMuW2qdc31C4DkMCJS7SS9mbkqKIdqT0c2yWtmOCGnuh13NFB9/Fp7OQStwEu9VxWV4gC21Q5
5nhoMpAxYRceQS5NfoCqDro2CCUo8rqqt4fXrNXLLgmisYEGSyHqBFWsB45aorlb98HGIOA3Dnx7
weerpfbY9Q45CwtGIn9lXafcjGGSj86xeFtqEWT230hbkZ/GEruKE3nY3qT5DBY/35gPBFQAC8Rx
Afw1W3Xu2/a6gTov11yCCCWuKXHpAEUG05R6NOtekvGmAw9O2M+9SS4Nz4VkX6ynYHaGhY6eN23N
78DK9kKLW2PaB2nqbb7TvHHFiHwgN+QxQzToG8OXUIuomiEssBE+dnSuTMWaxEJpuF+anZNigpUM
GNsYsDyuIQIZQamllLMeTTCCQBZiiPaeGSBgjOYJXSlQ8LsSaJBPayEolDvYsSjPDn2rz3jnGKV7
OxArRK2yM8VmwJy3AmsuD2EUyhOC27aICetExfO/RiTmjRtIhmfX+iIiKQyWa5UV3AqXzZiRpK+f
wgLNBv4oxlD7FPdyGJn3laP1m9o7rNBtAnu4SoUB+UNFlij04Yx9Q6dxOV6Jvm5OndRjJr5zu8GH
F/6BSFsagfqh+b9xJ0dIqbkOW+1x1Nr2x6BKvUxQJn4eUrm1M2p6r60aCE3NRm+rs1ZEdLAlkWLx
WO/FP8EzWK8VYSltd4+Sw5tyG/8apcocFTWdPKZAz5S6D0z8tyImIVoyQkB53l83Ij9tqI0MGsLt
CrhUR5woKNeLX/4ZbmzFAcufVolBzv+sUgtLjQS2BYxHfGz6R8X5LUVu7wbS1BHMCwxrVuXR5rlh
m839cHV8cBLokNcKthbmy3cuOivcisp96VwgsEEEAXKMgcMW1YUUJIyg52zdG9Tum+YF1AzbNveh
zrmQ4FXjauHcSwPvFEc3Be7Ppthce3bkQmGzgHs46NNS56O1lOQuKNa8VCEEH9liTFLHuAwOOmH5
Gzndj732x1UZORMh+6k9Po724KsT8xnqjwCmMdAwk/3aMBGovkqBpg5HMhjLgEMTFqjk9k3B+xjl
+u9HozoF7kHMrdFlhgbfQpnVSdmeYCB/wGLRzyxBjzU3aXLOLnWWN/KiBu/kQxh6FN2RoVdVni1B
Sxio0Vu+0jHRANCBVFPOQoqUJy+k6ZIIwD4QzURiVbWjvFPkLW17kcAurDdQg62ngvbPuMguBglb
HInAiKmoZk6kc1E4dKc8wb41CYcS/RiDbwugzusacoKAXh8XgKI6x0vmwj6rAbfWNmaYzVamPTNi
tVLddOTZrVzit92dWldUpkE9EBL0SItT5FwtF31gwQnL0ZEfcuPOXetwPhM/HK2agUxC+pk+FS7B
bQdleJ3qKEWFq4rGbfPS1X2lLiMrHj+d96JkNd1Brdi3BLN0Hp8zdD12SIGzGwpExs1XClISwX/0
fpxHRXOClDpTnNSKRbJTJ4wrMNjDZyjZbp9XKfAOvkEd4ceXw2BFbCkZ4kvxppbS8i5zVhQjWGaG
a5PE00G/rDWCOsewDXj3+XVyuJeZIdb15tOCroJrc9Kz1oQDraspxbODrziPKkXtXZu09EPREeYv
UC5/l1g2XJ7hq37oaWHL9QhbFobsM0n++LfahtYfUx24LWShbgJ0vVZMGEGMI2ZduZdiFoMpXA1c
ih+Se3UC9owNueBPR/EMqVbGLyN9Lw7cwRxUqZQXkTVM4tUie/sMi4wdNluQIzPUHdesiGjwa6w9
a9ylGNv+gjs/PyecglCExpYrWsS+FFwtmo+7qlKscD7MQwgOaw+uDXYYCz4h8CExY0wUis72z+5s
i6J2BofwwetmR4X2QdFGjY57OzX3AtDTir4gjUp1Hx/XDiEM2M+oDrpGiuJN6eHcSyirD8nwC1tc
UWlw7ADieVP0+yG+di8THAdPf1zvEf6wdD2gzbSYYhr/t6nyu1LZhdGY0Atm+b0Mjr1QSC2bF8h7
+PM0I981eUE0So0WwRDI6bg5qdc9Fg+oRIosaO9K2l2WuuxokLQpjRizMLnxj/2SWKaTadsgXzHr
WF0/01SrclF4uv8xHS2LuLCQOt+KRuWFO+cEw3caz57Bwu249OMaNctavHIBEi77kSwBUbj0C/K1
doiwOAOOLQBVVcJcxq2cEROw+QwiPxg87pmCtMfKkRsa2ZoiEIiwPuABMS58J9sz1d8MX7oUh5re
eaXTC6OOW+awoYGT6AaiaXmy/hBTnTOO9EdNFUG/mKrtf70Z4j1EhuPQ810ZY5hPEn2NRBVgLzTn
QMHYcFJsLeO7duNEEgif/fQMUi1sFtojLmDp7J7U+LNCRId4QyaWHMhJhbr28sb4fO88rTmc1pZb
G9hkAzh/p6DRBLsgp7FXnUthdoLkrNXmzDx46YgbvpbjaJYRgINCJRZODHlrEVLy5ni+uGSU9PWz
hMQDGMjrpXflZEMD1y6aAnDmoo8+rNc0G0iDWby7UBqvyJZw4X9rO5CqIViWqvcnivKAXKJMU0pS
S22DV6tUl1FUVyNVD0DPl0+YPPXWlRobjzt8LClYuDmuPFKpRp0iaiNTArlXqHg6sFpXr0wEeIZt
ZfcZCk0KihwUbKQX+7BY6qUrY/kwY5ZY9lwfZbk6H4rIpTAtglxAVa3uIhSEkNoSYuYMcBf8s3yd
5waJyAXVNyETvWpPjRpy2QHs8/zHykOQSoVoY/4L9JTflEcCaTzaCftMTBsVYkXif3OZCZXuyHIL
fEHJ7BbbPtvChoWjXY6WDDBAPxoBGquL+KiUxAEO0iE8sFCFlrkkCzbkyLonzuNPIsyAtyg5ly9K
Ii0k60ZOvomEz+UltHn0EJw2t/iukk7+TcYwOeCkUY92etPW/cUUrQ4hMPanPDv9gArtMjnBnc0p
MrCqr/MPc9aprQ7Eky1qJc72nSk8bqgXPFIrJlczyrghJ6DqJgUT249qrtQYjEI6olw4CySjzntv
pI5owfQfBEkztZePJyaeS/FdRX3Kwk2D5FY3CL6D5MnfbFpfKGq46V2RH5tMLNPHNKkmP4Pledre
mwYIwDPMl2BP0TBRcZCJ6da0NMdUcl0zk4Cjjnm8ftOBdiQadmOs7oaqK+qJ+M0sBk+kme0NOH2a
yHPcZQtuhRWxEf4iqc8vLbB/t+xl4kK8UhSXluyRM53YS18//uMUAWBItf1L0dk2lc2clWmHbIdR
fBjAf2r0iy0tSQRa8uyKSDyNujt8GpOiXIs57J1zqNgZU8kiqcqcCtj8oF2afs2I093STQFWEv6S
qyAW+CeoGmwEAuCaPxbP5mVoypm3qgVzoCUKE3CzPky0IQM9Wph8BcJcI8jn6Bt+ULHB09YeHjS3
73mD81/7fAutpEeDud0n1fu89uWaQWqtioH+9VPArtEoV+R6JxW/+RzO/d+btL8HubGokhXLnnxl
9z3vvOfOV37vQma+nPBEnzO06/wY8m6efVTtymeIgQoqvDFuDbYg+SmS+NMcDO4OVc9omLvxSLCX
Numd8yPGd27y4U/W+fbxyE+UfI7dm+rHEPzPPosUw+9XEosU+nmE7PIXYx4ybu+zZ53H+EhflE0l
i7mYQHyC68TeENNDMR0Nr0wSenfYTfsovrYN7i8IWLigjFINxJJZow25/MDxO0KYGH85HBi7Mnpp
qUMd++3hybS8T7jX1p8+sMQGd91+bH8M5r7OByfSd8sxf3JX0L8Kpf/09sK5phs1Zq1rRBILAkhg
jU6lA+q8vv7l3C9R/waAqVJw6vBztMJLAaDsB4iBhbTkhDuFV2UdNRYtzilTWgLfIW1XOfBZDL9G
hRdTbHuQXLhIFhXS4QmHWUoJUspMi5iIA1+sFm3j0iGvoxYEprr62xAWh57uus32/suS3gKsdzdM
7mFIjVmFOZ2J0tkcWRxweYyZS8nycc3Qd0GuxSGtjqixTfyMkMWY0ULRLkXkIhGJ8Iha2+yWlp6e
4F951m0MTjuflP3Re8Fj469OfjX6xZyQS2pp512VbDI7dFCv5oSqAtKOyl1BtQAbszaJMMx4jUiU
XBN2fCi+Ibif6jabj1Oi0LA9QT4A7e+gXOXLe0r4uc+vzHxOJM7PkxjnHAzixZFixmAYsO3G0mUV
IXWk1LY4gdGBWDmXFYsu+AQkVjeDw5jtXY4eA7D1jVT/TEmxltBqdxeNTdXUe35iyMEEhrOdzQ8/
lNgsj6GT+35D95QwVwnk1ntiamcNpMfoXhbmaie7eY8Wgf32p9hGfPcdEUjCZUa5jlUCIdVYsnQj
ykQy9fWCGXgqTj+V9buU6i6GaLQqN2Y6t2t4e7HEwhT5LTw8tfEU7xVDSXUfX7RuY6INR8qiVQKk
WYf41BqPjSm7VJpCIdDuOKJPIF1I5zfqIPkGpjkQN8xHbGbPICxYvep4mFrtBJdeDW9pgWxriWkw
MAh3Aa1Cw2QMPafcpSpJFffXVqOWsrkSd5hbeBKk3i+//J8lut+23iVcl090QP6fCxPK0q8eehG/
rv9dTFKid+CumXJ+qnQET7KTZF9gcxcb6EP8UzfqAIZVn+eOuzNK5rFjWI+KYlZOwReyqdSvR3+d
9K04Y58Co9Yo/e9OZTFxJe2erWSkLuL18gFGTIkyffGaUUl9ay+n0qct2SL1JGNhd6j/FlCdiYWF
iAy/5/qUBSzuMohnoWZrc91OKQqHrO8qx2p6OxzMuGXZ7Z6oJBtvKfKwwjAJ3AqeMTrKORFOlg/B
C5r2q1yiMsCwLfo6jW+Y8v/zVQ4oM7iJPcklQ3sc2hgKqHFWNsyQ88jzR/njsNq8XtAA0YGEZR+T
Jrjm+Bo84KnoHrrh4Pubkpd0MpRKEeexPsk99Yr0BZH486CYTJ21t3DnJgheQtZVALZJJcoA4JQI
kACoXTtL2SAKKiwkjzLaF87ONWzA/byKx27jG/wYav9BNT13qtNa7LjjlhDgTgOVQ/Ykgtp/TTuG
z8B9k0p/5FOa62vTaEkvr9WvWgLzt8s3ejqPqB+7/svjTSAZhRyhXqLeIe1Mf/vTsl5OeKFK0EB+
viZ75Q1tkww4vx+HYa+06gAQgv15CECS0MfbD2hW+TsjjMmclbPqkSUfoVFXSKTw1BqhphdOgEq2
CXAXLzmsc6NnfhV2UtnhvqJzK1e+j1+kYEXd4jCpr7GtrCeqDrzntEYhXNkEPAwwJDe3tzIXU9/S
b4z6CfuKF2yBFohTqV1uUHoCkG1mseUp5aLMMcTv/UpJsQygtWcMg21nGdw/6uNYGuERNtvO5og6
bs18PEX/YyzqD8UUd9YtR0lHOrwraDzSPUdXrYvNYh3xT4WCb8bFo6k8MZcLi4zTa10eC8LyUF18
tcHeGlNb/+wXUrTLmjTIydjPZ8ZEXq5a6UzC85LaWVS+lFXwHneeffumtFC1jIyNIP5zVTWyPq/i
/XyA0ghpSb8l3bJjcXsNVzz3KfMiSH5b3fqdyKZdY0PTPnTPj5zednemhADeD1F1H7xv7198U/sq
T7GGV+inNcC87t7idGdHTCvS/1z/L4oapmEpILPtKzdWp7dBF5iYuF0zWEcmNEcRsJkvqD/BW89L
cmitXBClx3BfppXZ6DBcRb8prOQPXjaGx8PjpLOPh7n41qW0rriuwMX2khVCSdLJgPU6HLiZVKRN
XlU3gdjgjC+CMdxkLfGkVN9wUxwIO1zadQ1t1fXMCexTcy9OwcKZuegzaUAJOZGyS0Jn946e50U3
gQ5pEa91vJ9PPiYhpTY1gkLiQUgSPzZJpZWrBOo8AvJ/Kgs/S9lLi/Hwl4cVlygYuxu6al1X+/j/
PYpBKnH5qGnJFpsvRP0XYi3Kni7jaNbsHhqiMzbIIve/Bo4Crq31nuYLEjx3Sxs0rWpVOPkRGXCU
4FFjK74iSXXgKPV75rCWkSom4mM4Z2E0kR/UKrUqGCO7kCFAmJJ6oI+Kn25KFtS1NNGmReOlRMyD
xl6DkJTOKBxiWtRUhkrrskBXmr2S0t55rH5Dr6GuQ1XzwlKYCSx0JC1y3gPw8dtHyuot0hWOA0gd
csYiLAIakzmE0ZtSxBYg3GLsRfTgQVVF2ExnBd0wlR0zigehKfaXqMTWaOGuuj4hN6nr4Deh8PNh
lqepjLr5MBcpG1/NiiYSyrnNAceWgP4+fnXzTWqjWaTqpY2KxTvVFyOTtMU+gqIftkcLcwH+BedJ
4+mltUzExNolrWvHcrbOuwTfV/b2j0imJhZL6HPcwF/qB6i32blh/2lBiO4Xx0RpF1jxepB6PL9U
TV2W4fOT83XKNQfG7PYVJlc5PAxk2Co+S3aEgXruOKfOSLOPZe5QRjXqx5mOXfddL26C/OjJ45Ms
J7Vawqq+OAwVD1FcUTTUsB1GgGLNbwtRvw7jToTu3KRDum5p067I5+s4WFRQ1LXR0uyEperszVKH
SFDxHV4snpK9UQuuYUByRf6vBP0uaU5ddLCNeMZ2naFlIZzpIp3cox1rmX8Ny12u+tWMUWKzYZ3D
V5rST17mYDqdQhtw6qwO23zuIQIM8sGRIQznonluvcr6NvbLn0lDN3OKurSba81dEPZMZJgPiAZ0
oEhvquI69ZfR48MTDA14LTm6CEzTLoqJ0TgSNJVSRhcV2zheJ1pb4Rwf/LZJgJwui4Tqe8aSIBoa
SIAk9vHOe3IEb9vaBGxjf7MlovSbKyqBEfrENGazQJLvkGDQxOVFQnLMq9BEDSKbOpl7D8jA4OPM
jwDt+qginidR8BiW8cZNwQVanNHNQyDLayG5OyiFwDQOVyG7P5A75hppWFEm3njzNynr8IG80yv+
TCxNopl1GIR5Zd5p4UxeBXlhdFQV77ppmYECKRgcG4d76SJkpCaENVJIi6EkfsAH420kCa9aaLM8
zBKyuJuDx8iOlL6C1SCzmPA1JHafdAK6dIaDsUigmMjFx8S9CupuxdqoThb40B6FYXPKfPe71Hd6
9xGpbypUzcBsmKkvHANzJZPgTQGZg3eUSpCO9CLr+Djx6hDhGuKxreBNruLoQ6Q1k5b/pXq0t1vw
xECENs2X+Fi13zPHxrjlb9Jpu5XYpEJaFhAfFJn2voegpMBa5sS1IqbG6W/byyRQKrQgYJiqVANF
ePZ+siwqpGu17DDu0tdpKWY7/oTglkzGZpr1GqlJHWLoHqT418xAyLLuokdgwlj9TR+5uusYmvLD
BJpXdCZ6VnrLqCTl8RKIqjQGqfKteO43fO//fGn4GSaW9b+ww09XCZPcJEWUvK0gdsMvTpg41ML5
cVHDaaYKl18Rnn5iovZSZT+tPwR1RjA7CSSpOOAcxOIAMdeyoBFZP36LLezBFFbjZJlf7IElBzra
ajdPRKJjcLrt8aPzSz2mQiOC7LnJ8ZZtWdLqaMSSSaJoooo5VtR8B2SrS4ub5xpzQrhEJT7EXKrj
aeknNJZQowfoqcuIMPLbDhHjKTbnq7iLsEKtQuDVEyZQ8S6+fnWdNFQQ47up1r1CdSDSuZBfcNu0
KWDNGfOJsTcGAjU58SeDF2IJ5/6lkNhji6fqs3yR903VWAf24suwTmSUjWN04trsP3/IYoxS308k
sNckHci7H61Fkn3VY5uUgL4dfGo5uXCtwdyXNQd/tXPd61RVoMoZxw6kfiYu+8gA624T555oBexb
v6GxgiBWB/NwTHRmmhNORm3pcoC+7a0dPHYKCtsIkdE+M2ft/TIZRWQE6VVAtvCHOaETMPlWjtjk
5l1cwVFBr0DyZS226EMbRhCOgEsZ8A/tJHv6h943a994014hnr97lR8ssyoY4Nj/dt2jdeFsONmv
0K/G8NHhN4tNBeVJHwaUg1u+WjcF1RQu2GKgmwAl/Z5NpanNxy/swkPXaB9oO/QlBavgki8eOm/b
r4Q4cOQqMqDbq5V/8trEckm+wEAUc/vkHQp9oTWBu/te72hYAMdEVC6cxKlWZq/Hgkd5MYmCeyjP
H9uWJo4WKfPvGpeMVo14wUB11NakvUjk73CBS7s9DyL7DxBtN9jks2Brg+2oOnZK31j4o05IItR/
txiV6HIDP4owank0uyB3ajNP8JGiUsIaGYq8ACxYtancOgmVaqOZOonChdqbgJSSoodTi40qWz4f
B3QsSe+AWkD+fWMaLfi0zsBgjBFbxo152cm5uHsK2GXLNHYSgb4jGMLOlubwIEtjDu3e3wiNpV46
KujIzcw+Zl4mmchEAHM8RZ00dsqnSPWCUt+2dwDN+jrwGKqSAAyqm3MBRL2rJ8zKmVXhd5yeasM0
+L8akMRPpVenlZYe6EWT4DohIvoUe8wAbe4SKrKa5kpOn5KMwiFV2uZo2lTP2ZylsMEBzBsAppgv
dgeOiTlH2aAbZZPVYAEB029m6XKGekrppxmFC3Iuw4n6FvOQ6RzbuO98WlI9eVKCzkpwqWs9OI2o
rmvZhx0Cm6IHWxvZQX+dQ+hY2l8m9i0+aVpalRfQO3zRHbndqE+MTdMoRHhmU+poqop4FDI7GZBI
wlzvg7qOUqL1pgLcbKLHuW6XWJX4XOaHC6z2fTlWeTJ1WRpwAMoEg7+EFNPQffPdtQMoj+/HzPyz
Q+flE/wXEACvZQVfbdkQAX/XF2KQiZbsCtzpMzleIhqnoAg+ywpqxKpud531b5SoAafUZ1HQvgGW
iPoKsugBYXn4S1vhXvrqkiZ2DwozO0Bq94Bv+E8KZOSvL/DkXIbymNy/q/eLOwImbzuP3Pik+gU7
ChWmgz08N+OSWLWstk5neLnIbr9gT9d1TVHFAmZSWLzqSwzS4c1rz2XK/faWUq/N+R5lhP/wZUOx
SeDOoGzDpSa/fjg5B3nnA8J70r/ZvXqDtcLs7aACsu7vh2H/54GlWGokg7yHMqvkauJ82w+ENObx
EOz5bTYuW9WeloQ9h0Oj1e26QwFWH4iTityPCoFmWbiKKbvzdHV/ujJbILElj3P8hYpsbnUCUnNo
u+0eVlv/ZEYCG1uI5ub2wGRkngmPRDQIpfFrXH4Pq4c9z2uX46LPZFTDoP/Z6QJfefoyCb4fV7vO
k+MfZ/wC2JI4eJ+2wKzwAzbOashMzeXafIEaDnd3egoeyMbZPVFVzxBtPEDhaksTnOsq0N+msXq1
lI0cYKiohJtAR5+qnKDMcD4tMifPBM4NkpL9UN7GKE/34EHy0epxKpJTHEpw1uX8VUwYDu9XFlIg
2RE+Hllp7d0EbocchvIEiZKY0FEkyRDnVN4jEeWzA2YBeihJgwPeOWRqotcmPZg+tWAEmLsqVUc2
WRkJumZCs5DydWOlesC67tk8UQk4xuAeup7YWAEUNSXltpyFCs1Wsd8biJLcng75xuAFtzype4Am
rN2BqGYINtZtaxQHIlSOvAq5BIx66DJKVbM3JT8z2CwPKtS61A8pPccx1mPnMPUa9Ci3szxJgXOl
5wKH9pw2F/SplrQyNf2L/kdPdOXnb/r/wMxgRL0+D6SKSIaanOP3b6XnO15oMgJRmckKETAmoU/C
k8sqSjo/b2vpWbxMVf3lJj2MvLHFJVU7D1RVRCBK4ZHVLqeSYbmj90LJmbLwFrpvVGQPup2YAc4/
RzyqfMOD9VE6WxYgvUM40bItotCrA3SVGUiNMhhC0jjn6Xb8KOZoFVu8/Q1EE/XqtEESYy1keLJa
UUi6RIpu4/N1NwjGsZqipLGROEhekV0skIy269scPRidT1GAgKgvn0MpPPsejwXkDCai/ICyyP9H
ySKVlv6yDfImHXa+KO1DEjpQvVPffRv6GbKinJoHE5JnJLiyqgDEI4QFqetrWzY3T4xTl9BaZ773
ad1MPFN+TmBxvP7XgzCZeJ5DlP+KYR+WulDXX98ErJW2/GEJmaMpc6mqj6wKXYZ2RIap4CZIaIqJ
eSVxFDAsSEcEatpoyermV6fmda/2U/tY229EkiTr/qI2AejOUIlgq2rL640RJzlmnQZUupmznaTV
hJAkKoUm0JiazZnTt6nTRLsYSwbF+nDFK/y+OqdknmOtMNdbNZjpekWn8VuYxAHOMntENzE5plOk
URKb2l2YO8wz4ukuqsVAih85A4H3+hH1lv0HWmMwCF6JCmPOT+8RDRAC08jLoH9wamUgYVteEVp2
rjJ0aqGrTMkJXN0ZtLPXGMGR/MBjdadpfDT237VsSa9oYXigFm6dzS4GZZBPzvmaJj7kR3+djR3Z
yxYR5pMwEBrB/RvVOCB43QfFm7lFkOApY9so3RT1Oy6VjezPNnRD+IEBbczfR0OIhfmDybaftpHt
9mc0LlsH93KlegdFV57SVlKe9glpcOjw+VnVcleGaMIOofVA3AAvSLpER21BEtRTGfM5hhvwhLtm
ZEzLun01wXWW2dIoA9sHBKdsAhiHBskPzncrPUAiuoOXVpj66N7uDws5iKC4775gvsmclDAnVYLr
WwvUDv4KjvGu10Pmow8tQuKOc4FqycsP7RbhrI0Fx3prqy8vnxuph7PY9YCSLz9E9c3pJgUgifBi
S+/z8sXxNZJ52GduyrvIK4U3+4js1C17uD4GfzvOoRzvkGmXRg5g+4MpsKGVcA4tEeZ4kg4nvuxE
H3sVZ2vnqGFx16vSnYImbvJm/xFKCbA6zbN2bgn4OVbB96opUC69JWaGCPA8t+1v58SvqxrLmHls
nP4b0yKdOkF1EU0DU0R/iWIKIN8NwOlA8YI+hUp5ROQDN9R7uQkBch3bVD+A9U2uFYK0jGySOVoc
XfkvnwECFx6zDZrKIKeHHchIaARErU09M8npx+VuW5EVa/U2xdnpnkXLl8kMiglUUjAWQKT/KHFd
4u+caev/BWYhV+LSaDAiQnZjTTmpql6G/sclDRZpbkRbcwSurctpTp3x01KdpqnKiQ4SgfI5YnOh
zEewpTGj46Edv0ZfPx2xVt2eVpU9QhTRXRLe7Ud3sCnB/smDirInxBcko1Jfe/7P3h1/nGUuE4fM
/oKptQELDXvLtEUBqKPHFJHibJYA5otxDxAzJVFIOxHeuAiODdEyjE3yzDSGx2Q6nAVIjc1xyRz5
IFqEwE9PFuZdWEpSAqvp1n21kqRndzTePW4vp5eZQHvpVvCGPP8PJA17XEDrCFDFkIyJ2Scr8/o1
EyN2s+Ociex68OIIg3nBxldid5ZTQxNjKCy5+Z3jDQKjR9R2h/2nLmwOCdBDXfbspcD4AiMAiiV4
YCQYT8+WZRqbnKR3E6lPBqpkOFH+BYt8TofFBWSRUhm1P+mblVGhkNG6SLXxncE+i5WqzXFdil5T
QOhtjxKY5EptPFamQGsbsKgwl6u6+jpgJt9jkO+IdeTd4nEbzdg3GrtTnbUsQtMWoGvQm+X7Q7E8
8YYsa/JuDPilYDUQ/lYbSzqIfyIGdDlFU//l+1dEwKT6FFUEqg+aJdJiv+KPX+gqxvj+kKsBTH/O
Q+gdATfsxBGvB1y5/ie+egCJSsGGn7fTIPauR7gw+a4TPBJHfFC9qjsTHRD3+Kt5X8A1m4RRwVS5
TKI0CQW3gi+edJmfmsiXDOVM6yjR0qGgtRJgkW7orKGTxvSFLiz7GabQvmPa6CZwcb05VXAMd+75
4CdXKEuShHGj+WCDyhrkCQSJrCn1x2PNPdNeXJCRn3i/Ol4qJeruyHtLjSSevI+ijPBJtVVNV4Af
W8t8h6xXSN9OK6sgmmQUNMkC6jV5ON8JsUUdh2XZ4HhnrFFPWuVh3IyZ+w2zpoVssBTqcHmVuqI3
Dv7qblVUxj4El/ql8kfmCvLa+CB2odvg6mlkIhGUaDdQsW3vxmBuG5iFlghMivoRtp/XTrYJQbgX
KvwbUbBF1WSICIii+Smbv0zviKFUevGNbCmErlyO6d5LnItw5xT/hDQHxyhJ8igcjOjvu5MryrzZ
xXX2PmaPtjnbfIRxBV41Qi5w4LxqOfasRevFHvSnSREK7YzO2DHpPP+SEHjHDZe/ISDvhwipIHlu
00FWE4ujaxRZxQwUPm0NimaNWFg+Z2TLMUXECkSEZY8r3ScLVs13Wd+67tUHd47e/ERrRYeVq+vW
rknL3WFgqJ/c2Q3XFg59hzxmKdwzjv8ILUa4wT+hmwdRZW6FUUqaJnw+2TBaLvh7dbpJvtCnRIEt
Me1/SjnaATXMTVhq6WNYWhYqS6sMumTpAFaDaOYIvsZp8CYii532P+n2eRKHfBnU7ccnHAPpJtL0
j0bdJCcoII3x17VagmBlU64z8mgtVm/yOnssTZ+pCW3K6cHnFqIZK4sIed1DiqSqvxQX+4raKJa0
GtfJoBRXRalQM2q4nPyPNcI818+nY4PyXjkHJVNzmtQEULpwUXu3k8VsGz/lx7A010JRTePPL9IE
eWdniYegsbv72tcaKCCrrnHY9kUDPUTlxx35174ctuu1s8QiQQ/XqLFaCvWme1jFWOGmofOF6Zy0
hLBS7wK98lkk8E12zPjONsso3DxpF27ApKnPfR1Qkbd2IUhge4mFI26j6/Mn/tNv377dc9MRHTf7
XVo23RRmbO06TAkpD00t647qE4hZTOTb8w4Lel2NkImyDCZliWMuawUMA/lZ38rSCei0oojMJBa/
Ijd2UIVdiIGEWjtBCSPGeyzJXwzxm67/5ldVKk5AsdwmYNna1VHTgMpq/1dyuIPJ7pIkY6LrURth
OI8rbLs3QDv92JesjwFRme1mMoILwsVF7cKCobpcajQrVW7mUfEUbvYEmCVShWXt19QasX80+w+K
14NAUa5mG+ZjLbTx6NmxtMwFVcmABBaoL05Qdw2R+Qc+lsLPUyIrF1CPZvY9wNVhSj5xwRnoLPip
eem4EtD/y4lR05aYpMpBVXPh71tB9MfRJ+okBq988DsSpHs/K6i6L8wnib7TJa1XPG5Cg7N3Mdi/
fjnSWufIYAW2T4gsjfo1JweJOjZKkIyNU6ILXql+OvkrJg8rR8nbIb7I04ENt6REXxiBQ5VFEAbf
B7gEgxYZv8PjwavTgLmHoPbYWjg09FLyA8IjjTfdch/MEcp+wHrinrPMxj6jE2PAVnfssvT8wE8V
S70eTGuELdS/JosPQ5eGA/5/EaWKzndHi2mNfb3ehNAeGh70FXfQE0ujJ8eVVQ87QFQr+Svjx2d9
vmU+xJcAse//eu23hilaUSEQZkyt5vmwQ0nBjgPo3BZzfoRZVljKEPmHhOnKMsp9BRchTafg0bLW
jJTGEdG6gRZceH+xJSeGmG3vXJaFv/Vy+4HlIwkH0iyJY4nL5GvCLDN9eoQb+1xodl7cBw2vflU1
ytNBFWb8J1KKfjUFBFTRJiBohWEowrV2X1NVZGGLOAOUGhVsR/YVjd929YAV7kAjBEnM9oE6bX0z
DKvI9qNTjl2Opiy0Q/JlIfpqEtlFv9D76mZ2x3a6lPr5CgOEdtKquaFhS4JoijroB2ueDngXubTc
O5M1qHEqlkWYnM2v1F0L41ZXouujp9ejjIXvmP9HBf7LkqbqE2p0eUflDHRx2TG++Pi02MrqsiBp
RKTMaHMHiYnoCqjCx2Z8DqLfnNAuv/smnBY4qulAGCdHho0xGMcYqQQNb3mIMRy4ynWgn2oIH6OI
2lbuOtxaIR9DjJsjqnEmuMVABy1U9OUoSR1gpZ+Q5e0MCFQ8v3QFQieV8cJCxy9Gl9M0c/MaXkBH
b3a4f5Fs5katwbmV3FwAYIlVzn7ooRru/N6f5lYPT3ctE/uITua3Lbg+bss7jUSqPDldg3oww82r
QRgg78QBkNMG8NkjPHQsWgm0RaKnZ7yeNhIC3gevbnezkM0/AmqHSDW5pnDeUvPjrzrrlR0DJOZ3
YpHfWsdf7P0D2Z5iKjSbYPVSBettQSCeMz+VwwKVJMGq7AkPfZTATcUsrKHeIdWJrV4UO0TWRvuG
PMHgHd+TYCLqGBuzJEth/0ut4ZL60qVLsqKkBA06gfOBjWS1MPc/b/ov+DLCKwsiaWVJ6NC4Qsyu
GhzQLLDoAFL8n3q63BUSINkQV3gYU5iPuEcaxZ0rPcR3w2eo26nvx2T9rIoer/RpRUElNUupFyKR
LSqWsjOp9v7pzjIpT/NOSih/SLYERK6/AUIcmAtlXWcABGihCmJWGI3k9IYVXetBk/ei08wEtjUS
3oVclVj6XBdOKxVj7KPIHrg2cmOfNRYseK2C6wAPwOxeEaC585R28InOH1dJkMG1RQZfx/00CtMz
KQqPY0Vpp3AIREVjPq6t6ylN4pzfUumH7piMEnOGeJp1QXf9NvMLaMcvc53venjsvteZc8hbj3Iu
q/SZ5h6XAdOUSPyTMZ2WTh1imGwus8lATpdsii8t8/jXGyKvOp5WBMnIE7RsFyfh5RhtgxUdpyHd
9sLPkfybnFBc0tzjV066X1lzpdzYoZpX9y1JWN2TKFZP08U6GHZaH/sS871sJqJLcNiycuoHuzAV
lekpJ5+GMHsmZPVaoerpbpefRjhnxJmlxveWg2Qf75X+YJf17jFSOsLjg/dU9Is5Bw9LAg3fg9AL
nN+QuSKEEYRc0l7avc3GinINkHjdYf9pyJDRtT6jjpWHkfKSFMDPoyBUQECfTQUqBuxASxTdzpLS
bh+cOPs+/KfvBaMMpVHZYbzJG35T/t5aHk+TESWWmXbYDLXLbICvZ1ElzG8ZB7lFltFVRafPxOm3
azqtZqKL0ZMNCDU2Zpof8Ae5dBCYnS5vZveIpWgZPB2zid+uT5alZ25513u8m+Q5rwZdOwRI2DWF
LSslChDguXS9U60UeSEMQ4lEKN/G/UNMOyetvYCXR9HXSgGwlwmx8YcFDsW388ORGWP6yAl7PNqd
mh9PBRxnoB4sWG8w+Xus5yKKbikbv/7aSZgROFJ4eDm4CKGXQ4pTYKZc9W9W7jPDKeh1+iNmWcPQ
uhqOVJbQ1kw/VMLKGQdgn4SbSdR3q0SaKxEnROr+jafTJ/7hktp7dC8TLydWkAlYQtuOvTQPqzdK
oVarYLTtWJxGHmMYlQNqFJciCX4XirZYQTq0kjHcFiV//cxdf2STJxqHEX4kldIIYMQO1bKjDOIP
/w9UNeI60YTmjEpxgIKuuTBZokfIrukJyAdAeAaZe2LuA+47q4w9QrwHKnvpBmPNnG34X9gh3ifH
ZXsCocjEFq5kHJZ5HH7/cob8FenN15zRfuJ+niPqIzGSqrIHJ6S482Ednr9KI5JNnGAGpuvb8LVZ
ONA+D9PglmynfqGXQjqKfUPvFNodmLtz7ya3M9EnEMcm0569r9eyYaNjg70Wy2Wj2qNhGebl+hd8
rL2stSTZEOzmc7HxMX6TQIvrctsGeIizqK/jwf1kPdaFEc0pLagOx3j+4X3z3Px99CHQOotyqD4Z
W+H5J58V7dyu47WkWIE0NBJesCVzuys14SFUAWGeOEdxN55ihZ6GfrEdVysiwM82J0vWLv28dSTZ
BMJMPAInFeA/XtPi1Mj+g3+EjHNxYMT8f/6Rj363/kucgSv6B19a7CCJEathwV6TzPI2TFZwDJ8g
5kR5RZiY2TvusEpsT60xGALVav3G6eJPT8pYtq0kuRZ1doYn/chJ2ZsUr/Xk5xfgtJ4Xk3XpWH2J
LZtGpF0Rsv22h3jG5YXUXwc9NK+E2ikGG2l3YC0sLLRaAnxYWALEdjYW64LxQWVd2dcJa4Fp7MXN
5DvOsdKRgpRGoY5NY1/A6BWN8vpe2cZzOjyRlNwQuZbb34BmjpgYvhZrETqWyJrDVIlnXdWMeofW
9mKWQd3+hxTCkSuviXZKxtCSH6e3t5EGk7uiEMTViEKXcyuTFU90UB4F0h/9hMAm1tVVTOZrviYi
baDcclUQM/vzSFt5pfZYdjFC3athT+jZTv8tV/8DA7mLogkWs4Ufm9W3AKIs54Jjx4fnVmFbA+bw
+ANLNe2pxPfRpx8uDfV2Nlp/3a9f7OJ0O6hglZpNhN2NZBAkREzeKlyud+XgHOxioNs0Pm9lZMLd
azZYEvi6sZ7nbiLPT1H6yXQlgkMM9fVY89ecoU2r39rseXTWVY/Ue7ktKKXHFOyO3z5vY0WKe7A/
hApyp+Yo++QJiR6nx9lA4QDZsWYK9T+mN+JpRFzWcYWQ8KWmru/8Jtur0RNCxSupe53zIMSPOuQw
h8lfnIxkcgtNuBfRAvad7Dl4F8VJoxTik9eI6OwzvQEsYUqOYC/AycGBP7ymsWbAinqTNpWCpQyv
qXKemIeyT8wqYRcFtDbudO4bjmzywCBPz047aDbc3SJWDEmCi6Fh04C6whk5knb6NLa44/VvNhvX
9ZPULW83gkQNP+TEDJFz6D+KxZRAVitkU4GGUe2xAUcsiMzR/BGKmFnshoB5o1rzDjB99EJL6IuJ
heNswl5N4CHiMjUZeV7RpGOMJ5ZlVVYFjH9p5vaU949VDIbUtgOnHPMHtX5LV1rSvgPlWloaMF+1
2MRXJV/l641o4wyN785MQ6HuGIpViGiNo7eoj3aBq2neXbeBAEEK04oN231gKqbrUj2uxBu2rbpK
McwFzNWluCDv5EbVqk3ld8U+7w4NN9zcwnKz3RIOKPfYztzImiqIyBVRO311Lrq6npde6J459G4l
TxXwu3JcldGJcQyGy1JhIF9a4oY3f6U7+cOHrUE4Ufdakb/voCFrnPr5UoXE4+2Dc0YS4qCXeVgy
/GvDhGXSPwNagl9vSGbWT9zADU+iVsnr3foMOZq3R1yoYv6emn8b84c7aopBHwnwZdNX96bAX0wc
NOj/jQUge2XwHajYRO9XA07bcsMRfYdiYqaat6KTwEhbP3r7U8T76QlDGVWxQ+UXqhwbMIbqbo4X
Z1e7ynXEbNlrMZdJdNCYeEQtfQRIBKJs4k2XTIMUsX4ZDe/jvkhMtd1kmSqiswHCxjLcIJOFcUVe
xnYVTmI/ofRF9mbhIWkSXWne5w7U5DFiziofyqCneJoTpLW2wwGXVMNUFWk72771ViXp/wFKsl9W
y2NlNnhdtE/NjHy1XWEGajBAMsYKpGsLzQ9mAKM7/jK9OkQs+Flb05BQYZ9EaIEntZrglR8sAoqO
3pQg5XIbHXEWOuRL5BgsfyqNMaoPdeOUyzS3UseJ/+mljUh94yqcQZRW+Y5NuF8toSgbWcqkd2aq
8CwFmf1oO6tzJdxTUVglQFLfYYkisO4PEWkLF4DSa34nnYtOepl3tUgbadfU77s2bXg13k9w20tp
MPjO9aJYzu0XEPFtDMmr9WmmJikTcdXfmYZzqHgUGToBMCQrRFNtkOxs+9T2FattjcXMrwd93NGo
3RBgvU+uf+vIrv+CCtQwxWdrZgsRsQUHydKK//tNn4QzFWwjnHe1GVKSZvfO23bJE9tB9RCIAfXV
W9MfRhP8gWOagIThbfo4FHLmpQ0QyqvuYk0Mo0qizSKtY9Uw+AJkQmkN6cABMKXull9W7pfX7BaQ
Fd8OAfBmylwOl9M9/+P02pzW5iMG4yqsKAq8+dGWbVguvmrmEHPSRnsOoXQsBHeJAl5hBcng1GWK
1W5zKUIne2+xOw4YpVVYL+yE4HsqeFWRcM8M5HnhyWkkY/Bz2VJAX3qc0aFr+QrWB4yWJts5HMCY
kct6obbsmUfUSukQiqg90DhPlv3ldh3YGYg+7r4qNJorW9ywcVf+HkOqloj7q4St7eQHlDjd2qbc
rAZdy+n2Y22KllPlaRe4UgXsX0i2+msUvyN1OvFEdeZ4UJ0ogSoDdDCc3D54GtP9Bz7p464b2oZI
gQUConJAfMx+qpxUxwc3rwrLAwtM+kmd53Q3sMrCPcHxLs4gg5frfAQa/kXAfMGYq8exEqJDyKYO
u6920Og+m7+rp8bcPzq781lqO2sViKncoy6a91vN4w3+NlY5vvag3ideEgrRdgah+Iio2GUfgLn8
5JJaG5S/pKIwjScGqJL+bMxuKCuQ3uMjxVmiG9GTPGk8X4NMaR9PDFo2akM+e1/cXz7qw6QIykk7
5bIpxRabwQcAhOCBqBAe38ka1A8rr4SfvaecLKCnfU4nuYOBWOb5lA6ahCdiTYp8LvZDXcU1wn3l
fdkVh17avhPc1rfdPcCnH03RrgfW8ciH87BRczxODYgXMU5wJePZGmB8PoDnLuoe6+ueG5NKAmhU
GfJBqOkeRF8qWVGR2yQlrxsqAEH3O/gyDcReX1ME2dbSUMa+jQ83XWfKciu7Y5+UyjWE2SPY3gIr
13FqZN3fZLceCMeaNffjLcUG80ynRw+i3crkssxwIVp77+ZCcTbzEuD+7OPIdrDwxoFASEM3uXXf
q2sfdOYxScvGb7VWB7BoGAfxihhDuKKrWLOs76lhCxAaYvCoO0D69aQRpYGv7OaP9LgMleaAX1DR
Y1q+OlZQ4zbVgVvE0QidS5IAP8QDVLc9r05VgRgd52+YtSBT+QxJALT9QOb8+422FfquGL1OrzVy
L+CyS6ki4qSlYaqdBniGP0Op172wyU0rOFxkJdaTTIdB0yZxxkArJXjITWN0/lCVtm2hf5mT6D5H
1lUEr3mkpN2Quul+/x8dEENwwY1hbEP1RpkJCTCMfkBbV7JIvbhV+Azz45mHv+R3q+Z23YjB74Wa
1Gt+wG6QGFognUEATo/L0ijO3PEN5uuC41U1ZHstmKWBC0OJ5panwVxmI8lihvA/ajWnM7yrC6nw
tIZKaZKjJw9xSa6pL9bYWxrCYNJa4jedQYmJdf4d/xGAO04jQW8ce5kBAULOKWSuhaWdwkUN66CM
wVtOwVzlWTHyTpAUaAeY6v5JJCA+u79L6+0pYIM/j81QL+e03uwkvi3KJgbRnF3Lk/Q7zfdU1XLi
sJKwdI8PI6Tw55AaLGr0d3oPiIZ1ZFf/a90iKtLHPc69P7g36T53kftLk5hphi4Lsxym+O0eoc/B
S6i6BkHkl3+C88zFtaMvcJza6bCx1u9VqdJbhh+8UmCWS55dY2S4760sInnelpjaLTYyXLmyCIM9
g+Hy/HddVrvEOBs/vj2UQQOa3FJvmjG3eLKFXWagOrsPnw3fB6YFiTeOlI4vTYUraEw5qdIVjttn
az/zz6dBrZ3FQJ3FspvGPMWgnp2JryQSAaWrGbrN3EEl0Pbvk896nldamZIu+/3lmJ4Eqd46E6Vo
K8jY1c3RK9F8oKpnxFc2MKcZ2tnZckA82Hqjc2N0aR111qijzkTawGo7wi19BBPJcHqdnMu0NYYj
+vrSdD/OuayvgNMqqHjZ7kSR2wm4voFFqoHNFU2BCj2JbNnSCtDn4oYWvdZXBn/i75VAti5o+kDI
9upzT5cRhSPNpUGGRwkp5F180ya+KD18UnFQzhkxuB4jAEV6X42IZ/hKIkJ0syOGoToE3f4HFR0P
XhYhdFFIdmglujpkSXPm0uNrF0tV7VruJ8pOHfL1qPdc+8fii7aqissNeaMvG3bsrv3Su45eEFPP
k17MHXCDOZx7pzzcJI+rLCly6TTGnZp7Vjd8BEH1rD1kGnwtiGUtuyeRXLzCVC4o6yZLkvejLrt8
LNZgzP7OzIXFU46LcGB2MZ166I4tVGx7ZEItW7rnk0rHly1bbbBFbUd3hcWMgOWQMZ0I/3a0zxII
ALYf6YnikVb3Kvmq1KXYirOJGjebYr4GJctk3XrQKBabmhBUpFd+xOVIc+J8Hr5hBOEG+Iz5Vctx
YZ98nPXkFcyevUJL0Tv+8+rfBn3/ClwW69BeSgB8uD2mp7Kuuup/myWG/xMLxmUJgekSBzx2pMn1
TqRxIiyB0MjuK4WiA7Tu5aVO8hMRdvMxROtbX5gftNK45gyfS4FAX/uT5zhz26dY9/aXEyuSIDJo
wK00F5aKPXBSb5I2o3n1dFLpeAS1sk57fv+kVJKviXj9fiTN6skgNx1ePK/TuFFaNJTuHd9Z9Fyt
Qx9m/2g92GpEnuMZ04OGq3Z/FvVwfA3wazTAnjiMc3rf4ocYRgIV7Igm/NKqXw2PIlWQ5WNqwyH1
VkOo2CFn/ZyJAPbOxRmD/C4y3DVhp7ltcDJ7sAZgMNx28aIhDmTCNJVewMvOparXmB0fhXOQZAts
ilNZcTv8P/b5cex9DgedzW8YwctceFSmc5iHesffe3N1Q6KjpyizmMupmTCi7F+5rzccglO+UYSZ
0Niy3L1BQYayCCVMo2WlmExV4UbxlrBU6UtA6iQFq4ciD1xNCFLmD9MX5tSd2X5Ntm8735Dveuut
B+z5K1fPFFFHsCuc+RF42S2dRXfRKR7g8oas8PQqF8eQEMZqydro4wZk1q/Q1YGjpZsXNFKFLgpM
2fmG+C5HYmnoqpkstL8CqKAXqgRFoxfaSAvtEc6kb7Prz/gp5ZK8Rv6nhaau0mve3MYYjIl+G0Ic
7ElfkYlMrtAEK5NldiKINg5l/tAc6z1yrs8NmX0dbNfjMMAagyRxEon3es75/pApDFhPj9xitup9
7nMdwmN3QwapomosFAisABi1ChKtuqEWuAVbtIV7ycogm/voYzVdRQ3V459p3ix+j4MKz9ykzKgR
FhhuDIWsMaNk89XLrR0xssTMr0WKpCZ+XyM9dBaoe59LRrbhiQKroboDRpapR8Cc23c5EDbaS5a/
x9XXhfMavypIwLw9TEErNVW6qinrqUE1vlPcTbv8mNqhjh65EmCwsq2R1gop64SapybWUcqLv0RW
xtuKrgmJuT+SLUfBdl2ZQQnZh8Q0BPlFQAXopyllipyzEj4euXzTKAcmmtvxKsrdVPGJEoea2KQN
PDJSsmrWuQ5JAS7/LIRXStxvdxspRiSb6W0F44dg1rUIPFkyHYdZTbsHzXpoEroKej/R/rAT/T5Z
rRxzDN38ihJn1q6Zuflsac/G1FZwiwqEopVDzz6joEpObxeRW7n+toWzMgalMbqSd9+iPvSnWRAf
QIVuTW8ZCm6GaLEchDy7cZmHcRvm+s/i8DHD4wieZvZbFjAw4iXU8ZlSuH0VbR0xo4D2aa2qX8zW
HA5E357nnf1Nd6y9BLWyBC/dk1NauXH7K9cmSQwWZCQQNRKiKI8X8RvePRljuvbX93f7nvjkff9l
1UOdVVjce9MXtJPbnC/SRQTY1yzSgIRSuaPaIizQPekfcuGYKyoUszz3erRfdhP9l2ivbc1zJYu9
MV7biGffOtA/lAYcvdJe2L4qeQhgdgxt8dczEjzdqoibxPok/9MK5fzeVYfBRWTJDhWLNDryCvRP
1Ltft7AWp24vQHO3RbvxCvKUnqeW4N/d720bh7HCn02R0KcQZbD8+gWr8Ln5xrb7ggpNalATc9LM
m8Cdd6OgPTAYPYwEwcpZ4u9lwI+xGe/eKq5W8+P0MCCJtV9zkPE8oqSpPSDXhIFNO/kTq9Fv21BH
GZgpqAuVlw4r4Gf2hHSPQY+qWGiWB8dj03nmH/U8gDFN1z4JklK+dK0eriR+JDv24zD6BWaM571T
iVgUWqL3cERrJaWTqS+aEKnoFS0edEfWpt+hVZjRhwzlCBON+PVw2rmLAvEPkSatynx1C5rDwzGw
LazKW0chYKNkaHpWVNVbYbVTjO1xXJ0a1RSfh3gxSIc5cXe9+/jpERqP6gvJoS77loeS/4cnyY9U
wxbouv56CzKFQgwh/j1+9l7h3+WEhV61/t2PW/kKXcftxuetzjlg55eFiB6dCBSWOcuuUZfxCzGK
EBgV1pgGAlRAu5K4o6qAHVMPLnWjqTN1wYK9V52UgaopEbzwJ4EuBNasislt5GbVeOZ/W9XoIA0L
3V+k+WYXVCgoriVcOHdcjqPYrX+0ejkw7SZCjXm9zMSbY05WATSRKS+RGyYFvOSG/pTWZkZHXhrv
X9wwbQBI/pKjTbSuabTWlCbmNj5FsZJSldOzn+9k7JSDhMkygor1rKklVeUZbEaC2AV8Q1yqYGaz
hPg959RNHFZOuTVocd1HWs46xe9atvz8dNtcnPQMk9xMtIO6n0UC02aN6pJDoTPgbq0VoZ/aWAxy
Cq2iRJaeiMFEAOmM3eIkFnESnW0/0APSi6GEjRnpp0BeqvKnYsCHZ+S4EyK4uVRBm7VsJuLLVkjN
81VZ+5F4aOXULuPWncEMiirZ/jbqKpPhHKw5crtmSTHFdMy4q0MD5KKPnvM3IJk37hpHlB3UIFE+
Sd/Shmu6O7j5NLimEGE5bRQ9QY5/BSKT+FEnBJ5ehGYicy2Q8dSwdDpkCAtaGGFeJ4ApWd+RvsTw
8M+7q56/oaUi22U4IdR0Hq0kXN27IlPU3Mu9QwobLPIX3t9YWb2LJqpxiub6riPx6xtbSbAxoBY/
EJdSWhIli24jdGgQf+G+QnKLA/JpTKilFSVK55ECx8VP85Vju0ncxwstJYzhmbZ7qsPf+h1PMj6f
L1oFN4NGJHBvbrXQoZxeDYmiJf9s/LLrWm87F0Tu9FGeQP674HhrxFC4witz/y0kgmj+UhYCphEk
Ei4exZwJqyelXzV3V+M2qoLljR+vklz78wiq6J0RDKXhsh/px/xU7udQErsaDTp0hSwvraKYfU92
nCVC/BEYhHjsmc9ZP2b1IfoSNi+DT7O5rEEWplsdVo7AKjqygmL3OMh/GYbYwTIA7jQtfn2i2ALc
myuaApy4MyQ7y9Avu9gz+9UotjdRjFyYBfLemuH+DsAB79MhoqShZPXIVhVFsjdTGNTuSueLVL1n
3QPVSOnk5b0N2R7ABi42Frl4tzxNfoiQNqo+HpBQxbrlCMJdfHUbutPDhFwRo6OlYeYkEddmIkzC
a7m/J71p+GCaJfYDfItye3Uy6iUAB/H4+As5RHX+L63tn/aLTzLpB+WUeGGCV577hb5G6K0tRBfa
Th8UiMXd0N/n+CX5S8OFCTIun/UclEi4+dp2ku7KGEU2Ct4r1u9bioLI7oUtIdOg0ue7wNBE1eyV
MyfFSdD3uypYe5aLEsOm9Rdevjlri08aXfg3qoO1seRcfobEmcLRn4aQDWQmq89BY/QJWhwAG3hK
UoQTvtmMedSYBj2dlUNEz8mtsrcPK60t1vU4b4q92wxFpvuUa2UpnQC6XqhlQb2ENNXUuV5I/xKt
hKSfKlmRVutnQSZYUGn15wmTG1rrTgLX9+5n5lMCUJUvdQFMMCnANDOKdik2zu4NJAw7Bj3wW0rq
aa35OUNFEL6uB+shFpdqJjbTp1a8N104z9r7V98oulYspU9KBQCR8/ilQxn+6QhDdrQochAeyxVX
rMHfOstnmWIP/H4HWHTOKBVlIR4UQBXlp50NrL/RX3J/iWd3uLJB2Td+bNSKgVFbPRJzA+ruxgkH
07wO+WI4dWMKtxIMeDpT7MvE04INSOmh2N9z+lu0gR5Q7M6hyeZ8Eiqew0MTQaFI9iAPeBeF5Clc
PqdVx0/jn9FG0fPOXblFysDYHX2VAdGdTD1BAskwQhS4oAoyQlDqHVf99f/QRLI3WWnoSuM3OBUc
MLyBVweGS2e1gyxN1NjwqgO+5GIPhbFDnNqG0n6GjL/nv8h0Du7QMYYBtLY8pSU9LC/6Kmn+hSfU
+NoI9s/mO27GrfZKWwHbKkA2dGBJ9Xp6+2YdxKRNBJYsQwWYTG7jSQOpEu2Y7Cs96iDjTHeTY6Of
P/sPJZRK95k1s/PwkFYFhkplIoh3rAZSIKJrSwhxsdKfsfytVgfWDnSGtUjc/9xqacph/jrUUA8n
+AKoYjZYxMg5LN5GDXgkoU1MK7u//+WkO6hGEU2aptACgMhPEGrHBYiYFqzqI2x2iMH7rTCq6iRb
AS7vvZYOEEPSyA7IzJ9rNFl/6HopRzdT83TZG+G7koxEUEEDBBGlvpGsfIzRaqsIZaDtbOCgEalN
gXjNF7UEB+P2Tjc8Ic2Jchab51rlgDJ8Xc3ViYSAZDw9h2cPB2rg2YhZfxeABDfB0wnUR9arLxZg
aA6EZNtdyXFJXJ3k6Xy9bTAA+XlyfOL4tHJu/RFEDmNN4TwI3sN9sXFkwl5YXMhBZkJ06hMjHXlV
znNvrWU3+o1M9ZOIbJPXeehL1cvvXRls4AmCmNNG3zuguQRrkcDdXDF0yWP4bhylg0v1SAKZIfGr
f/JazdteW0IaRnoFSJEb2Jr4HMIBi+cA97X97gPd9QKShPQQxfxPJtFP5j1XQCtYY4ZQ6rN3JrIU
f/0DOtFZh8lD0ilpUP4O1jDgV2bc8fUy5/HDMROw+K2FgWe7rQ6t55ztshnxsxhWkVOKdR2H4AsL
I2/jCAn4MuHip7AcSVkCDxRZbAVs1gUsFG18uniGl41BmB4XY/tCYY2QV4/+yAQKPL6zkq50GJT4
RLTL+ParlQYA/xrWCQhE003QMCeeZ1AisldO8dMTgZ/dQN1F9/Xzl59TtkleIA3IA13JXg3DlbkI
fZX4j6D8mlydV4OkLusrVGgNjAiR5xON2uUd1nNbYApOtJm04Izz1/pgmPYMn72LyYeHCEQPH3fX
HgBVEg9tU8awf+UdLRlNOV0sfd385OFeXldYxTFj0DV5kcoOEc7j3r1gH6Y4yEaNTvKXG1dRrPmK
dF9radCzLEJbEVBWPgExRbCfloklsdUl2GvLhUpyLXhbO+VKamtavv+dWrbMyiajFkWke/azukdK
rEShUBs7MLSOyXwzOVzyrgCAs2NOEEJIrA4dOBnWAIKVdcVR0hDGGvYG19LHb8C8GYInwaD6gLgS
20L0SPqxwLsz6U//n3jwFqyTdA3vhKu8r68i6XEq34TRDbEKnpSxOmwdJAWb9CWmxbKHrGL5rs9a
iJfgcqRNMJLrjpeXlXwM47iniXHfTEBCEHB0sCA7aJGLIEyTjJ73gWmH6RFhLzbCv5ZyrouQujCz
/iH9eogXAu77gtMwsgBzhaX9p/E1hxrTXOqGKA+2dE5UCtDpfgS1N33QtdIeHl86b18DLUm0aBqY
aWVgKZBFXip9DZO6W/xFLM5Ip2wX88F40lu7kDFGDVzP030jfYTLeHS0puSGnUcLNJXIRuYChNGC
zaIlSmwvRbD07joTcR5w8WBn3GXtaAZ0X9WvBwya+hNAy69bp8WjNAhvr0YXcnrXmY4CMreAhaBD
EuCmvob0wxOLmpNOgl+0wQrricAQNrI5ldg0nRa/yRy0hilvZnWwvr9/MvV/pYhO3mnsL49g1qn3
GDlIi6CsG+I2+Rx/jLkF7oR3if3sjLaEB5DlVLlJMflm/RHMdX4GwoNpUJcMvEILgNj1af++7723
j/hSxDOT35sLT10868QOwPeOuFnH/wKRajRv/MK9iNP8kwxG4+tgm3r8TjL3JRwI9LrSVAPB+jUW
aJcbeqluX/hAHy9kX0qZXV18Mgv76C7eNDUHDFdOuPlFk1JsyHe/9Wwun5Ql9c61pPAsKK7xmH4O
QpGCLrnbpas1oXj7JsWTxr1es3gN8dNkNQWoPdUlzjInLzs1HUARq3n3xIhIcL7nuRju2d4JPjRA
tpGjXQIzSKC/vXWmSxXrcQoUvqQhDW86gfnyYK7V1UwcBWM+SgMbm/7KaVfw73ERpQE03RNtX+y6
m8f6+sqDzDThUpsoLZFxK0iQzoQeP0k8ymH9kCtFd7LCXhmQAdZ0capiRZqp5+V553rCrDPeHMBa
kRoKI5F9KI/0sUgBYtTDr48mjbHRJBNDPlGn9KqkUa967aVmiGMYT+/6fN57hbvwRsqrKPNKL2YF
7O8FskP9KxjulRgylVDZ8daE2wI2Y8I7ovgz0RlLAobS5Z6t07kiGbk9OixYwb1x5nxWYCj1HZw8
5Rx+R0YRaCSrkiVxrI9DU0GuxrukUtBhUmNXd3J+WKKUl1dRawUwVHpMQPPP+8CEPCRGThH8n/98
o9TzECeE2E9lfvCqQOErTgR4RbKUaH58I1DkpAb1RHnFhhsZIgD5rXk+EFNfVOxIMFgwNdN9Ca03
WUHmDRh5CdtOrjkmdA6+dgor47UfoHs3q9dEDQL/4MH+guzn8Fuu15BJK6zkJ5kkiINKTUMF3mX6
RI5YNe9ocdfq7NRRKYxUkhofXDoWHqyb+K0cFQsgArDuEbNkv2jDXffqK5V2or3P9lBJeVgefTrc
XOWowhMd3rTrYThuqPIZ4WLgYIjf6HzP60Y5whirbQUoDbXdim2sNPLfy3MdqTODECCJHVTkSpce
a6HVnjGKxa6q2pLauwhvlO1PJoQnkalhgwHij+87eeHYQG5Fj1EJkTfbCRaC4a4hnfmPAbs6ZjQl
otOtvs8vuMLzFpNmhw65cJAeAhG6dzD5VnoKBPzGEFT84OUmSl4Q7HtUw03sTo6Lgd84KEQQV007
Ew7xPxWmVaEPHQMHIj6tEUNfYxCzeIQPtcjbAdbOk85Fz8fTeu3+WjmSncksUP+hNFDCoIXjnyGm
o+xyxZ3ieNbLuZHNQvs7dU1NYUsd4IIf9LF44tg4Qj5IHsBqmx2J1B5EzPH/cCge4PVM7oKMkVOy
i8TtjXV/7M6soQWXP2V5q58KifDjqMNF8GJjR4ijcjTcow1WM/TWYofEKBmM/xVXpEanKxMWlxBN
mUPs2F8k0S2BiPghFNAVVqhzHd9Ud2SbZZ41O5gTFLXJlump5NCFOenxHohb3NTPj2PSSXM0Pynt
hic3ggGHrkVo5Lm1ImnejjNzfeHrE70fWybsvEx/0iV/kPaUK9SmplIpclWMUkJe6an4b+yHK2gB
A8shGSFyAjlnJHsVBkGtOkiML50vJDm9Afi3706h+jkzl8JKYxfbwbCooWG6YmjHroqOcwAk0eHq
ycrTj4IJF/Km7qxM5G7AWbfPCajR4EW2a6FPdNFWL7CpupET2/A5qIsYJ3YCx+5zOElKgA20Q/E2
SA/Ej4JmQwG9REIzoJztb5VQvqRKqC5a0mEndHD5d1Pdb2pWBRtzUv8Q55fs9/WQNdGiNL2YgKra
eO/Ctn8Ixuz+0zwniuPqE50i7iUdUvcfJnAHNETEsf7pmfIZQZ2TNOc9oRSxH1NVyKJQ0xCSuMo8
W9cBkYT75OTZpGGlJe5j5VNF+OtqvWUJt6iq9VF2mIoFHmEgZCJ9dNIolJDi23eS7e6XLzH/OnxB
UV/ePTAIAZPEss/y27w92/xKQIORXA9W03u702FwXaXyhpLLPdu7vsYnR28qt4FXY8j5x5fulj/D
7E7jkw1xHDurQqbW1FwUe0YnWhY2hKkE2r65d8s6cMTCy8oKbsQ/1HdkoZafO6BeHfLF3QLA6po1
u2ekOAuASB1StbqTKwn5v1tEj9pRMz9zPkjYDih4u7YhcQQ3o2dXajAfTzvuYDjzjbF2aYsPhOzI
w64x+dmkb7FKffkF0dVYRVi1VX+ZuELmFIgdryS6z8MkY32vK3O/1qzK42RRYxmZ1080i/iapGyF
/H8ibUlWHXrYEytttsxU2pZFF4ZhodBEw4rsRuu0VeFq/J5pGJo5lz5KmdX7ja/+7ofsYr+FUwjt
f2ui44VyLKLbGpA3E9xfDKZ7j+0rKksQBWd56WhOwuByw41PuLhBU5SHSYrquQvf6saBobZgOzRC
azxv291fYDXX5FTivIh/OPfyAlLNaVbTsy8wR/AWMH71UEqJOtAz73EGa7DokhHyFt/rNLGGExqA
flDTYLI5+zRgNN3kQSiyq5UqYfePet6ZSW96Q2bptTgBEW4SmB4+cEbXLgVFbL32h4QGv7atzjre
2cgtK3rX7643wSY7BdX2GFQ18R8RXBDCZtSfqtrlik0QLaz+XdUO3EH2MUTnP4ZySSB/ExTtGrEA
DMSG/HD0XHYMRnO66IwGvxo3i5tkSfs9RJn4TbbazhET0vLmfevHWR+uV69skASKITsroBIhSg8r
ggXIcYbNiMrgjEMlkoGoixc1qm3OqdtAM+WLJZrgelZyXsnslbu9W4F9ulyjtk0i4phFNc8CDF2i
3E/bUIWuZlogry4/xM5CWbTWTlK+791YAbiM5rfO7k2X+o9Q+LRBye0vd/lZqlipiOyyiezOTN/d
mWIKe5Qnm2c3NjHlQyYUd5iQqq3LkRTCd1jodT3vqkFBtE8VIJJUXnzSgeDVUv8DON5XnGH3s7W2
oop1rz/3OYsCiLHQWgmi1xntYwOwGMmCnqzMdYiAMzfT/3tsKR95zeTslsVOMcCtiViPGVclFayy
gpmLUaM6p+O8yjCAk2I0QMQLLYpigZWDu6jNCij39rB5sVspd1sahcuipL97zgdrg5zN1qvGQEWv
BkDjjQ8VCveqU1YAu1wVL/LAobYPmsVDuLU/22ziJWDYeO+7wTa5Uwm/vPb6nrxpNoByDmtEFnwn
S+ihPl7HKk8ckq1flL6a+T5b32bC70Pa7XjWZllfNzJPSijIxKG6GFZTc0DlvIpb98EEnu6cMKzN
QQSUAdmv3DdOofMyUVAPrPfVZne7xYkIR2I9LVrHhLiAAJgqU8Au+22IGfhLLaJ354ehPcn3NnTr
jZEd4hCMpgMxpJoJU6lAUurB4nOs3FyAVxsm7wxMDYOyJ//DJAKphjYFSB4/zxX6ppJ2pa+tOJpj
NcoVtfSeaBSY0V7r1xV7k4Q5/JHxwJ3+5LzS1YA7qz6tPUBfLAXzPjMpQ2a3j4feDRI5CY16X9dz
33XJPartIj/jwG3st/zp+TWsfUvPQ/dCYWuZxt8PkN8kAHPutgql2dSAbW91Owbg9uOFlJsHK8Km
6MlkkGwBsC2N8Bgy1OTsntmedE5hv+CPPU8YvPQvyvBGNo49j5OEphf/kLfkz+Iu5pndc2piORfW
cia4Y9fFr/ziSj+xd85WUZfMnJo87DbG76CSyvG4meTsv84sqJ6WCD0A37ansHpGkyL+UEiont74
4BKiyp9sYaRXszaOphEcTVtqQcG1xC9kaH548AyWExQEr5/yqJiofhThWrjk/Lr/Db+c9Y/lULyp
3XbBFmrcteWDo0MyPLiGOVx3/TLZ0INp2PpceVjiDjUtDt72xOJPvUyxuPx9QXS3vFkdH1WzlOJ8
rFCbBrDf7Tv66UgMseCOpOGu7Lec8a1hyPCfjOADnywBuv6OlCRtjqD3FpG9RQs3Lb1DLgCJrs/d
jfKZq8h8RYnoQdMyxh8nB2wsY7uisS9EgrA3Y8T/Tpi7wver8lFOITnR/bJw64coWE/9KFeNXCWC
uBC//7qmUqM9SfIppQ/iUZuGEzbv0ykQ1AWbcpToyS9sKLme1P42JLVTTzbeegu5NwN2ZZdliGpI
dKWjuyYbEPfTFHJslnmif8CnUpG1jfvd9Nd/XgmDKCUd59UwhZgUq3MroU2kS9nUG7K2qKWygcts
VyQMrUYMjjuW428cBhlGScfck7ERLpavghmfbe0UQJE8Uz0GSkH9mIHAbJhrf917hBneuKNfn8Q5
AZIWgos0Tm/jsuKxoJTuYr0Cy4UUUbSn5dcoWyj3GMxV1bigDSHwXOb+BGNAwKdNz/KxnOcWb8CJ
0c9P7GislKbfSIKv7rGF3PDyiakUcbJ5cqAInemRhNGQJi9MUFmcKz79AY8T89Efbjz/Qd7ke5+o
yl8E0+2/adYJVHCnkr9GOhiNdiqm4B7WQBcBjjBim/CqFijxfXWOyv+QK3BdbluA4dvCd6Tni7Iv
BDC4Wme0ILjq93x0ughnV+kWJ3gh4xbFCyi3nmQUilUj4CN7DykUL/jzVgeMmtT1rIVBRBKuuQ63
Gj+HBRosnR8fFZmuh+er76j3LhpiKjP/XC+4MDBsJgEOXeqv3zEYW8spsXE6eXYSvEIvIZgXxER7
w7Y6ZH9+46l2BLCOIToBF+jOI/nGS02dNXgCrFdH7P508oHxvtXAbf9CAXnK0q1xzpfNLgQdEMB2
y7+Kh4gOh+Kbd0aLYf8UhegkIjiJtrM1taao4ZZMNMJFiH0SYR5Eo7UzQ3wWL7uMCTqRpQrVl8em
wTRXKu97+XZy1raZhyS2srgKnzLFtcB/K80w1AWKVc6km32T33ctMReRXJGOHfkiPxwAzNQl5iSz
FuP4dLj/rv+unGG5OXDWKtTNwuedcXm4OXTQqy5BsclYd5tpEdlQFdjTvUyoNHKNx5G8dgVK7ivu
yDRe+YeQV4YQkaDl6XTJIv8DYzRWki/JWNLUDbnJVr5pKIaSh+UuNexVE3y9WgPe9YVVNrGkGsJ3
WMlrJcBeTWYqM2rrxGuzughoVrpOqpwdOPU6LdnWokd5VjXYLlqGDOjwFfWxtBfWODQfzHjqUIL3
yIZNA5z3IF8sn0fned//pJz9zT6JIO8kgctH+ZRafFxJR3S7Woh10DAV/BEvqS+6tEQmcHMvsgs/
H3cbk0BgmJDKlQAckjDXr8LXsEZ2pSbLlVANJIW81rqBeR+qIKpU6ozIHMnWIJ9/HhaEAXPqvXW7
93LYBU+h5MIQeB/icJlDDh7bMPpDWXeWe1HLsvN0CUmkx7fxYfdOMtq1piGOVvNDhdayp9gZdz38
wBunBURSZV6lEESx4vB5OgIDM+uCPOcVhXhV8OTPTxM0Co4wyD1BYG3bhJDD+8gClV3+z5tcyqAF
H1xYDCnqsZyVFcCmqujbRwkpVdDPcjpA1FMWOxgk+RT9z7UF5IF2ILgJ4ijEY980y2MQ5X/4m56W
tybYP0ccWesOl2IPHfR2LfzjU9al0XdsRR9DJ/+t5CkfzvlaI0yOo6UeKdiZa5QV+6AUSljdNmuu
q6MCuW8GwIjd0MXV2AicdcBdM2mK87bP7lsfgUnr561V1HAssHdqE4ip6o7RR4If6yjwWTFmSpsB
6swZoyeyet9Z4HqzPV7JGjursyDGI/8Ndwchh7I4Xd45ZiB36ttm8d7MBuO62tgMhonuG7YDZ7CK
sLSr4SSjI3Vq+iYqUCPbUop8rWE8CtGKjUNid2YSRFOTOOjFgzM85T74aoVefzQHLl3Wxg7kGdO8
vbApzgiSdk006KzNikPT544Mu0JHLzhpt6kriu8nYgmdlzSRS0Pg4E2VxxW+RRMVWbDS8KZTn82/
KAwhiR7dNBGfQwiq5AkSyOpNfNbk1gBGsNP8JdAdezrffJol0y5tJ/33iCowr12zHvzgNRTFAIF/
x34snAM7I0CsYZQkxtxSdEr/dIP1aY5OYBM1EDgTx/ZIrPTpDHbjBB67QSjSzkKJFjM/O5mIuo3r
r2/2uR3QU4mInv7tIcW1IsiwmGcFuXNPXmuPxS9jsAWgytllESMWt9/D6a4tOCv1zJ4DMaVM29wh
qLsmG82xOWcHe8+T7W3MMz5t0GDv12yvNfDrKAYPoAfn7WSo3UUCjDDg5Is7P82mG2ulblN7EbcX
Y+xu7pUzuOWSbIZoFunki0gvRmLw6E9SWEbYdKzm9ZrMpu3M5toA4KJxBOPKOwYk8KeGn3xmuwqX
h8UjWalQmW8MBMZDvUZSAgqDJFasO88tKf7qYGEDbSzt3HvBVNwyrZO27F3RIc97zoWqUcn+9/RY
rfQ6LpLwlrk8s6BWuiIcmXtTD/k9vrXv48H82RuwB1XzTJSf7NaY9G1lXrDhuI6KqlQwKEmnnv3A
LtBYF0NgI3HqcRuUCA4mtoF1oE78a1l/3s7JlrDq9oRwrtCSBorGseRSYjPSwMhXi5eCn3GY5Ywf
6GOdBglAWjhrfROWoVInPHCTOIqzbnxqB7L4yX3tR3zdhuvwRhTsig/GGMamxWPqByjmQfFo1vAv
ss8tmeg3Xq4BlklxPBEbyQMI6pviCvn9NNcDGZX6eVe7uCrTrM166lgT8vnVYb8aVX/dkO4hV9Gg
82/3aonS4G32QTnhWXY0RYu5q6iMrlYzT9fam45iL72Adui7P3zWVQnYVySIZd1v+DVdw8w2gbNt
0B/jUpVxwhllhrlzgwFXt3AYak9axrWxwxepTkLDLxe7NEFfyFw/G0DNZPde1Ow6Rpg+dv1ucUPK
qkKvP4NIE9037qBcUPfIPTOtx42rt6AkAflYcoSBA7U5hYJ1oaJZ9AbvFHF6JOk1ELKHl81bHZ2a
IOt+XBiCX1XsW95+xeok7JKyi2qIOZrq1wFpKWjl/PnczurHYa1zHK9XYC7hHVq1reGFc0YLWZJE
CL+0KVkgjc6vpaRN9cUzDQ+88JXE407sFd2ulRnDAOZvhvBa1ES9uenjvrB7T6TUG1ZuYaSHgMOS
W8Kqjav8P+SIpM+4F1WtG2etQXZ2G5QFn1KP7i+xSeHV/77RwMz0lJXW8tTnq7Tw+u27RnpOpgSs
yqnaqIm3Btm/m1TaNxFTAl5kaEiCgXhXw1Mf3GeFMqR8w2UpYsesfc+QJHDW0Lr+z9yoD6rz+7C8
zdHjT1t7kBXtFEb+ZUKgDbxSEh3o37wUiItIT/v1SboilPkcYADWGpu8xglXRya9I550jP+//IW3
oeg7yVQHfhmbjkjMryHD/sPtXe4fGG4wKQo7WLWjCHfFkQvkmzIqxB6y8XoY8HB/+4hvvkDzEX/b
brYFZoAFsn5goI/jF0eOC/r8rlfnYFms6itLVL7Qe0rZ+j2nBMmZvbm7QV1fjhruXiOychZJaNTU
kH9ifs5y4Oe0o/Bv+VOxP7VPYsI7Nq7bvYVY/oQAUhJA/FCAXcKBdZd51eYSuSSRgX+vjnMHlYiM
KatoMYx1Ermzskj9sN8cO5374gCZl/OLrK1LN8VnpC/9Mg8ZhvrQbhl3sKk9kosyRObAVhsARNXQ
UrwT92RLsv5v0fHIA+RUv0EPAdtkrh3rn6H+K23TQZSMXCUnHHqe7w4l/W46SJGaTIEUUrT8H0Bp
XzdPDUWeLqMepKazW2dKFmJ9hyzrjNhmWiMm7xL3JpA7JYQsMhfrAGH3s2UJNNcRJL5tVfXao4Va
w8mVpzMdab6bmLLJg9gJkbrRgcHNqC++7quElKVU+v7YEwn05elZhIpBv4919WQyg1EoImGs1yIc
uNOSMPkxNCE3qimUWW/FHaWyk0wjFqihvFsw1BJ4jOpL7F9BrSzMvUp3vKw2/lNDAT/BFUodwq0/
QNySWkVOG+kGXoAB+Sibz3tegcPzmBfvEq//ncbRzZJJ/+jDQB6LzPzgq/89VhzXmgnOdhVfbjkZ
xxypxAmH+5ffD1VRUhW+J3BR3f7BVciGrl4yzTA0UbBqHx6sBPW7Ak7JDMxEwykBcbRgoH6/4nBg
Qij1OETjUEyGY/xQDAGJC+ZE1m3oNCH5Y0KwskOvCzawM2uqXR57yhaWgb2LzPfgRIkfQnGLGRZS
pvw/121S60Stwr0fOy+DEbCdlBEUSeuXbQJk6gOxrfVlISTp3tu5Li9K53GIBiPMMNKKptHPRfJf
2bQApTK77uNtg0orWl1Sqa87FyuH3wUOi2KNzNH/msd5ukVv/mOm2vwIzF+84ZAFyA9TEjhIxd2O
xE5vHO0vwLbox1mqHXYwuhByPN0TwMbLho4czH7t7eN5HSKAy36MXM8O9ZTxZ6DzdF52WsEA5tpI
Udn2n/3okpR5BC2LOC0E9Awm766LDrIKx/faEyL0w7dcoefYD6ytsSQLHh/fGGiMx5G5C5Dyp+8r
SyhfcavHIoR1dQqUDLdh1dDiMU7aAPVI9fR04/BwgoV8HYOHLGN/DGK+JZNa2sOD5yiGP9bDZgZ3
wUHvVYJEX+p1g1cG1yeosD56XEWfD/SMoCrG0fLOj+/auvn55hgj9lhmknK7zA+0LC771PP96U1T
L0Ygp1P7PMxHUOEicsFnqAWI7fJfAbhHvY8gwBylLgA3jEN01aBsJXrhT3v4fUAfQfHO+1Q4CTh7
BCmPtRWt6xtm0gJuPNABXp+Os09TMQE+Tv2Syc08HI0R6osrln/OXxcqbTtKvHrEf5rKz1zzCHxn
E6amHdG6PtpsVGudebyUussu2qZd46Wy4dS5ly4LVtQmM2Thb7GjyaFx05Q9TsaOpsqGK6KOMA/f
/unXLDASxhJdEE7M2zAZJRlnjt8zwVCaBlWz1SFaX8t3CrLtwVmpYhe5qI34lyTjy2qfdFCT/sv3
koO6B3zq+QUS0S1Qfz2gNVPQeu27GSgg+OiPwfRSdRmlTFFMoBOgl1QC0HQR0prbO7pNOTBTJX2d
7xsW9UPoN7704B+PAE87eou0qnumHJXeSU15yBxFToKbHG0CPeLU6f0VUwR1kwX9e0r8it4Hisc2
URS0PpJRMsS27rOmFvUtoce4JTIrFS898VqPiX1YsUn5HUGIeevQ7ce1cGh8QghfDCimFxZpWu0B
+kWVSh5wkxkq5vVm3fivfPeSkO0M7oGWmwyciaIByyr4BlD9Ywx1T9v9IWK/wiL+DrRaj8wji+ZB
pZr5GUDIhN9nPaL9wUBItrBmQCRIMS1lysAA6wKkXvPWR5bEmqbAJDIwtWzF6QQ/C8Q/zKJMfIzH
8Ovl7jDJX7IsRozBkhtcqaNEoTGCV+yzB3BESyn/izJJPpZufAdSGOcz8q+UiFQC30aJVEWDTWN4
ZEDAZSCJP9vg68/71qKvXgqb7acYhnTgUD/GJ/ydDGyPacfIz0w4LhKO1GYSx2uRGO0QNLQ8bR0H
f384P0zKKGQlaXwb5e8Pca4zE9BsBVMFrChjplqV7hc6GBT8XmDkQM6oq8ITBWawDuH6cpkmvBkW
wsKr1+C00yt0t7jNFXGpOGioPQz2AMtWxTl3wCca+v/zscvD57LaBD7ap1XleKTrCQDDklwY0pwm
aZ16qOsaMrH7FhNk4n/Gkt4oVQibx8uMDPOetS4ZDZhtjIFD1juFSE6QVoA8bJ5PIPYcyD2onbaT
1hFP0xtSMoBATr4L2V/8EGZDOERY9CUV0bZEw6e/9cvxEh13sbUYLvVIFioN0gDCYov50vO10dVY
I6c4UeOy7OhK52MGBJw2XjSSUSP26SiPoBSZAWt6ohDMTc/dlE91PEZpHLWMEzOTISGHm1+1WC9R
b4LKbK2R2LxcI3RiRAazPArBjUkjcOkOH3mFfHnsaFFb297hgdJuUW5RRPPD1HnpF/Qh2DkZZaxo
apVjbJEQdRXZkEYbRKc2NRRxHcYkOPeZnOs6lUuJFAuz3iisbc4nAG/SRyMXL2dnmVQJHyuDI0Uf
2v7lofq01L5nRgoagSuyNQPFjkQcWK572lkAe3ASFs43jaEA8gRCBqshatRAOw9Ge907zK7Ve9Gb
u3A7ri95VFrJfJe6J7s9xFV/Rvg3t4UnCdCEU491qIeaZKdrdys2MKNzPdeVVjmjGBcEtZZI8Yxp
7UzTZW4ToDrj+7jQgyZ+3RwsV8ZisIQF8r7paoldfEgP/d37Hvv79qZO/68ewQuJvUaNpJ76rDtI
rc/yQx1sY8Rb3x1Xq2MyBiDhjHdCwHTspU/ppFh0qrLdvzK9s7/K0BOogGRGOR8Ww/C/aFo/9bzD
sSb18qr7R3jgcuCOqgU8aLbR6LeDOqN2ywCdkTOU/+SEA/LVXfxAKKUUsuqWaq754xYXMDhIipdv
cypGjOubrMPJr4p9d/L7rM0iqMgInLPlLYWlyCR1Kstl1wiJT8dNci/QmF9aGqkM3O4GquYdgPQ5
hABPZ0qJLnETxck4Avqiz+wNiYSDoB8Mtkks9QKiWKG70ucHf1dnmHJYmWKTUX3olw7k2O15XLuk
RdvAmqYa6rIc04LTn/5qI0UYqa3Gbx4+KHUZcPJ2RFAGHv+DYA/0tQS9D7gcr3xyisc1J3Te6BBM
a5vH8Xj9No66qI7s5yxgwFXvAUNQYWmOrDBs6K5ZdUk9uXNUZ8b2Sk+fL+QnYGfwqsQ0hppWmPUj
s+HTqpu0yS6uphI6TMVAmQ1swmscbjD5MIDex3bvciYOyhy1EQpee0Bh9ui3POdI3PRCc087lNb6
dIvwpaar2cxE21Ouu8KMoPwIZ2XDiBnlzzFKvobQ+xKeEG3mLsvWt+XkL4vnbzJ9Zt0Cx9zyusc/
ctChtddvge0wqM1Of8J/291D1em2gY8NcYEXqjJF5BwCQTC5joRVW8ArmwqP9LZleTXjxjBIw7R+
ALp5sa+zOgCF79J4HMWHoosLycpwBZjZZysr2fXQ/rT2pWkHQrwnlMlVz9bvGncNjCD42VTsV6fo
lIhSw3dWh7Ff8Gch3V7Fg2vuk9l1yVlvfUUUznHTFjwdXyVJ0B3xtcNrfNMZGdN61H19I7BGy1Dd
pxRfVRoYuVzFwr86YRaE74TV1gclvUsvSv9ItdoEY+mze2STLa3vlAFdoxetDKTNrGgeWBaDDRoR
AWZwWG3bW46NOmS7iYKspaZlTVQPUCXGc8dl3mVqdiFEaf0WD45553I8AKrNPhcis8FE74XQDAw3
ZIuagMnQGcdFM6GUe/MZ0dt/JuZ7OgSRIz+lzcnZvS+/csiioqC4eUa3KwYc4wAruTB9Qq4sgAyF
Il4oWxQ0Lerwubx0lEr0xq+A/Ua+RTZUokl81mEWZpH5w9gOuwFnXUqtdESwPPEgFNoodRtLOyvT
PAZgdMNqkMDjNr0fymHricSYl3aobJVkfiaHomnJymr60OI6Dp0TIMGCYC7GIxLQgVuxsGW51xvR
xnttDEEiXPLslucEKNT7m/NXWuGaOs6MYw4dQg0yt54RdoH3a/GvwuayZcU1ftHMsdXlnIc31TRT
FthAxWhKjCjb9Sl2rQzLX5Uoq+T7QpfTZcQ24IUQlVx1zsiO2HFgSV5jZDZHxA6dMX+tcgOAMlzl
++QJ7UgxjrS4bucOFeeSgaCVc4GsJjhp/hvaSHWyPJt43fr6QV1UxAG/VtD1bmZoURt228XY/a2g
ysHTZxH6xfkq4jJjWXGclyQsvtYcB3jdBbazZo4D2ekpqd77uQ1LsukAFEmX2ezZIjqyTFkb1geV
t424xe/qVNwUWWf2dRiRuG2S37lughCTvVb7x6yhw8/ZWP1dpVxVOff3dnRuH7i9lY03e3qrjHAu
kmdfepSH88wojPZFwSEiSSh/psqzU/GjaLwpQPxmh94bANQUd1HsQQroag/dJ+N4v0d0JBXspXER
EpANr7KDEtnekkKO4+eMaDDOHOc2j9HtiNNUSL1Ls0FhFWKVj6lBi96yLAKPmYrT8jVOpgabcVEQ
giHGv7vPU+rqwoL582Zkwom99EaUqDiTHcKpJ1s2X2ds+r63MuflDZmP2Bf0Qpth/xxTvMhExqOo
ST3ayr6NdETKbj9KaXhtR4ktsZPKJugLh1VGCjNP+1RC/tla8HCnpm2RayJcHbeUlgZnfPwMWnp2
93OgpSuGNIq0MfLlrJy53L00joMnr9XB4zMizvRYunOhuMVpNWihadXhAtv3crX7E8xotGDf9hev
nkw5Tha4lj69U9IVTOEy8zdFbBssn9euEqsuwc8bhPkgNRvTN2O8trk9FhK27cGl/bzLT0ASmtME
2XAp0VFdPzUWySheOtAFC49Yed4jDq3HJCaNWAx/aqOFY4b5YPfirUKhr/xq1V7E4XfY9n2V/E+i
67JuKyO7kI7l4J5gbVc0FS/QOeVUYDdrcLC16rLyX/dYF34Tt35ev1DTUjZkP67qrK+pWn/ciGDv
uPYYlbzaZrCdM2vFi52qoXqYWSxEAO+RixLnmnOpI3X4giaXDIBGsqdLnXy/HcQC8SrPtsPbhvpW
YxXtruNN+2zXGHy2WnIDLVP3RNpstsyvvoop1VwR0GslKpP2yChP98B+vYCP2Z6xJ2kQnU6usw+z
gPDH8F/p6IuSTt43iyztztZl1LSL+0VhPia35RtnVKuZPv6MFG26tre9d1HpK5E/XkFMWtH/d5KA
13co+j8UuX39B3zTnDVgfrEujcyWEiCxyuKTevJOmXMQgQdo0j6mrBG+APV9SQElNDhXJHAnMoFO
9KdNJx3C/RkMwv2el9d7zyHA6EumU1gP83FGyMdEO06zTSDKODyUMi7Sn4iLRRv9XAL3XzakDghr
EX0a0SN233CSpXpYOu6qVYxjwt5dlP4I2jj9u8Yj/AkDfkn5pxzk+iCsGhYk+aVWmM/SjiFg/CDb
fAEuZUMHayooIPFVX7Q9V6KnfHfqoaXN4dhjH7R2jBmmE8QN5EcJ5+AP6Q1YHx0xMOp4NkQ7yHLc
koMTA1k6skXl6rSADtGDAVuPMWmgBg5P0fsb9Jf30ZG1d5dDJUCIYXA/EEcrI/wtO+VaEtQGoytk
IuVvlVU4yovTf8QI9siSehij9FiLAa1Kmc1TVdZCc63TStdwUx8ERN+5sOQP5TA+pKn+53vDQ0s4
8qSqS/I5FZkNKz9DWB4I8Jz+zTtzzlbM4WRnNFqLhYU/o6T5MsJ9Qaxf2J3/YVb4YR5c8DkhKjG7
9BnBujabZ3MZF65/7Cus1XH+uOE7ZNeedE6aQH3W6vKQ8EXe6uUnEGu50R7K/uwweSDV+9yxjLr0
kO9/rNy7GF4KeFyY7v9G3ETMOFjFbCQpqNtSnUKJbAXFu7zaMnPwFf3MpqiS4zWL9I+s1umfXl04
RPl3v89DVUPWyIq6pLCxWslN1wxvZBgIu13fkvl6oGFX2Yk5yvsDmhWkHy5k3OsuITc1C2oW4+e1
QFJbaoMHw8HJleK6/stkpdm1+FW9OhVK6OYbbPG1IGpUx6HsHX23gtgFnbCYOpeOdBCtEzTqx7DS
YoIkC1EmxKkJyma4p5U7Pzd0Yk0rchst5bXsewN++bjYLL5RfLrkHiNqczYDBgEs/KPVGwcI7gcy
OlfCexzleTWU0Y3GJYYajO+CjuiwmXfeq2MzrauOQAtDeljbb52W7iXUNpu/uVB5+l5NS8cmlNvu
AE08EY3JR9YS/YdvUhVsJyxfbJQhLbt89QhPERxVRS7gB1OfodAGdq2Zx9s/0AuAMIrExdqjQwO4
929oi6hNnWUUbi6wS9j/a8f64wKrCe+lWxapRegwgb0Ct1GA5HmIV6YMnYaJittL/h7dHWeZKP3b
J/SOPp210563IGEdnTCPnlehgKBvgMSVt4tQjKiILTZlfao3t7mKwcBmuxPpUxQpOmS8M3R2jgqH
UkH0HK4ke9i4hR3lihy+tTrRxeBO7bGA1ETZFJ24w/G2/JN3c4vtQPc4I8GxIoHQk+bImNNW8jHn
dfhtXOOUw0uCJTzBBmxu0jxryGLmGhxfCSQObMLvx3V1LSn98xb6Q7NB2FTsRyQjPICP5vL8D1Ng
8GQpFxhNj5nbD8qq9DP+YIztug/p4lUgcEcyfeFpz7XVwkvbApWHO/TWSBWDU46MYCSZWMxJWD+7
MblkuuWcHa5Hp9FwLZ8AcUmuPC9FUVC/nWgLWkULTCQgsmnlGuTcGwCQR2TIeALWQ4lo/e4i2RsR
RMeI7eNRvUIYkHDgOsipFT+bDwWbn4WAbCq4/8U+r8bBFLh2d25Q0qRdIQ+RhTcZKhxnW4VEai65
V3N4FVDPyqsogippxsKoSMFDcotH1sHDfweM5kaCv1pNVqVywmwLI7YnlONvnoTplNwVN1vPg3Y9
bU4i26Nh2WdC8um807hjxgyOVeyVlNYjpqqEQ/iS4aVdgAQexUX2ZyztPQozUZUPf4/Xms/wtYv1
c/UH7Axo2KTTfOhguxCFsWimpAe6f6eBQ3ZYtjaibju1hEMpnRY6KG15E4L9D30PhhSZD4EtSIwA
ku6h3bU1R2ObwZ6R54vMjuQ4KE3ubw4XDB5BSD/AhoJp6wL33w9f7+K3LdrBt5MF3DH1YHVbSrjZ
E193dvwgHZ0nKlF0hOX9CoUfFw5owSJO/Jlm8fCSNsT5BkALQqKDXWv2z2Q1/9+sxTGBhsMyNbCL
qnx//NO+X0crtPVTKS9dyYofN8LdI0b4pNHeeUzV5GrzHfkyPRL/ogqMKEtLLVoIA/RPv2DM4w93
mjPhQk+3TQdeLOu3szI0zeTKyhsuPjjeq8MgZKXtZ1J2KDAuUamEU8wFxebi0F1a4dwt6LhF987X
bkNHR7kwHjfBNP7WJTUHwJk200uZoYQuHZ8xV33F/k5B5lL+Y+57a8EafsPX6izPorVrz4uGy7Kw
tHGs6SGYn/VhgapyqRd7CFsoHy7437mZi7LwAxI69ZPrd7i4rD4tlsPUCXrGWYzmmVmKpRaTswfj
5LOXdUFy4L0UfOu+tDOtuvXDxEt+Y+ZlXOLmWPUoopzJxpaHM4budblJnNPrCYFxrEfFYCpYmaOs
upO+XyLrAq3MVMjZUR2WKCwA2XgK70NDnYQMKOml+dfLWGj921iovxLiMSMOkokii5t+h+yd39CA
t0+0aWsB+c3DnG8MaJlEiNQAx805TGa5EjlsdNiRBjPgRUSiE/czN7/MpgZKMWNxmh3nVs4L9OBm
GcGhVolqHluyQXj+tdJhdzaNdfXpbi6JltHfNdgqGaC/5TljRMrJyEaUflAi2/DvUyYo9gLP2NDS
9T8Vn+0J48YI2tfk6B7LUhvdrqXc7itHMznyMrJ+u8U2jsP+ucpBQDFkQoxNtk4NPPTN8XtCWS0J
mHbFRB0wuJu1kuqVr0u0BQlFEoo/SnO19n/Vy7OgeMLkLOKg36rnV5kzOUF5necj+y4l/xE6OMnL
G9m7l/VJPMf0bqVqLqepyTgQ7wfF0bq46j4UVPlJxL+U2Kl2ZIEZ0Jz7AeRYyM4S1U2ACyzbw17t
Dmrei0prYRdYQS81V2q7ZZLK6CniMaRCWmFwc5vyTndbv//IFKfpkJGlPRggt5Q9Rtcv6LlT2lK0
h2gwRe0D3BY8d+hfIe4rDV8f+FE7Bn+XYKWy6oGtxOtj5b6FSbm4cLFj0XZDO1NRYBsxnzhN/+9g
QyvJQ8AlcA5DqfwOw13VeN+H6auNDm1K5wkdWjXa+5dWQXS9tmYhOSAuLLtmONR1JmCh+hI4s4ZG
lBD9i0y3O0xPNh3GQhaz8YyCbm9AlaLxrhPQzQYHkG5x3+evhpwUWJAghWbdY+UnhCl2hoMY8UP8
FV8c+JH+NPbYACgfWylwm7RC2/HFr8Fpg6unPJ+cuwCPnpr+qNY4QWUaguKVMpx55fVnDZtt2wEu
S1+IU6SEnC3p2BT52p0afuOTTS1/ajo/4Fa7tJmz7iWftWPkgCbCzUvGhLoQgr0ZABmznjSnmsOd
ECXSQlpkqc12CARuX+Ol7OUdakaon6t41I++H1/do4OicJ4OwjJK0INz2pxRIILJgCrprJgEQcNP
ULFiT9+C3SlndNvgq/h+PmfxzkdEQWrRTHeLFiodJZm6jy4FrCG/5mdNiFGKRA4aKsY6vdNEKg4Z
aAaa7Wtb/UPqkpM+ehp/ydyIVnnYj6ne5j9WGT4IDPRrGml9FE3i43WTkuZACOI+Fd4GVp9bIza3
2MYphrR0w3d99OnTxoAiws0OhEcEbG471o51u3ZQ/ITdILyri5FmyDihaXDRPFskhruovMOSf4on
D1c6g1p9/sYqUciY7c0ZqpjGK6MbFraaVdwxJodrYQ9mLDfmpJNSSgDVzxz5THHgJlnNw8oV9DtT
LVyMHHNYapiXSZf1bASHxEJGstRrv58uWvvLC9qgO8wPLNLcjZODESs1hi+/Gt6K+LO0M4TKjwSb
XmQMl1yd9E/lDA2ytyKS+PdLBsstxiOFJq/dxWK9jquE1211cE+Y/bt61cr52JBwOyK6HPWLyRVS
eFF6B6gPmKjzLqhDJ+HWYSEgugwwTWe9n5N7VKwGkdI+hD+fHApLKXfC+odgEJCjuYIRz6FiLIyy
KSHLkEI+qc7csUJPjUB4sES3tsdIZd3Daujf050l5IHIeJydOiQ6yKpLpU3fLaVXavJPmXW9xRWN
bUbjSmiU1bp4xdmJz4ZAe8fpAYWsE8g3lnI0iy9DF+cULDX6dMtU/S+F7YiMqnGPeX9o7HxRbDqH
SGULA9554DO7GiCfxTEjunfRNYrkEpJDBCHXD7d3yspmVTUqd8yVpviP0pf7hvJ1vOKIDLYnyL4F
OPyaTNP7/9AG+iNPdfUduQ5TtI18IvcPA6x5WB8sdMwK1WgppHSWOAQ84ujonnmkoUFuiV5xgJ1r
REHMXixrAdLYP2YKobyT4Ogx2wJktH4wKWqc/eNO0XlZ0gc+lpr2uq6+SaNBinlzsr0kOTqp/a57
YOXiSPlxDMFIPVnOF0RavknTdNwbWd1mGQSQZ9lvvcs4fqfo1n1GKIM7r1nVJxG5kUihYbpI5DL7
oJhax4tl/NOZJf2LQSrR+92KLleitAfBz/zYWUTKS3VAJxG3Es3z6jOLNZ5vsIgRw4Tl/DCkoRQi
twaD2GDT2l/B27suiNGDv/erJvMOmxt557XYDxLR73YHH8xE7R2ZUivMYY/d1X5YkoyVllKeg0pq
/Wj1CXSzTtLp0RVIuqtvRJA+i3DeVbCVqoLdXVHCgOZPcEsugGtW1RhqIMeP1I4/Y/S9kwNLK78W
44VymrmeuWhnhnj2pUBtr5wsojh1DK6KO4q/TuyQve9bd1Xa6GTarnifgeUnaXrHWk643R3k+fLA
KmhNWpfiTC0WE+clU2CGqD3h3XP3XjOxr7yay21QSn5LYFcOK2uVtm6MreCNDy+MopEsqxe42gOu
QL5znkE9cFqlg6Wc8f8aPBZb2PKccCOxLrpvctEiyvTWo9unEE+kjtjCh5/FQvS0NOvMiZYW9C3M
Tyry2IUbcRM7I4FhSNKoDC9WxbmJ/zHH2lEj7Bhk52SRMFhJ2tXT1ulFQLzbLhZXytol0VfOEmW+
K+Wv/frLrvuZ1P3EayYjO/oa9gWiLxBPc6MqqaksyA5D63KGU/5v09Z1uCHAvHtqduDFt6FnY2Bn
X2cxcaNvlweXS3nHaLeLwxW3BQd4UkUr4zQ8KkPJWx1vJe0GTmHkzgvCePi+3NWGV6JkdOFETNl5
Roaf2gWnUkYLvlhmKBo22ECO2UQhSJ7nQ45YDxsm44Mo4HN7Bs1BRP7p7mf43uLJI5JrC/1ddWfI
RVK0psBDwSw8x1sbozvz/STharWVm7sbAytLEXnoCUcJbENZGLdEKv8oQE4avN25BM+5giNRvaQ6
/paJPw19JAmjBS5y6+ntlV+fTnSqHuAuyqInvDWUX8PxxRKfBqjVU0y2HGKwU0Dh0SgpQyH5iQUs
HVJttINZ8CE+YiZRFeJ9wDbaA1sCnswRTAmA44v+Mm3g21SC2H2T3fvEQ5p7lIHwNs0lLOyhfvCN
Myyt1sMV2fDIfX8v+BCrP0PND/DaZruxxACC2xWw0nhOwnVvf12ur6TNDm3smdZgUC3sh/i7yuNU
DeMaPF/Ov0wcIKRjo14wcw6Z36NGVuhef15Q0/SmN92HzU0NRz1I09jFmtM3jZF+p6Sw/YpVn0jD
O1rH1N6dqCscA8UTqDRUGKEJNWjRHVzXfKlQZdOS8bpuVR30gbnrYJz5jik0K83NTTgbBl2MTTNt
fZf+ioDnKEbYccW0GQQjDw1oOSQKWdJCu0KRiqnYsZaWM/kIayttV3STkUGaHWuo0Co3OsfarkYL
GPEW8468Qhiq3q0OxsqKNG2eBJ4NEEDg9PxD+XW7+GlEVPLX7RuP4oqvsDkSAK8ZfX5DlNNlLyLZ
20W6ZwTNJBudK6MfbCGRPlqA30ij4hMpZYg1oqY4Ux5oMU+eGwqgto/fvC4COZbeIVeH4m3qvH3O
lv5tT32ttVCtGK2hKrR7mjba39+XY0F/bSOGqhe4/gcJYQyGkv6l9Dm9JV6aeE3V0QnrYfL+K/6q
x316TrkciDnDTAz65yRnKPEq0azyOcDTaR7sTSF0wItDBXIqNKnLkJWofwqKrEgFcoREUlMhCWYq
+yDPonYiKKHIrdtvcEQ5jJXXtv8Ly6+NNEFCfnAznaP5yLqt6f0hkOcqoJk7SIbUEpxNujZ0kBSE
7OxnvN4LzLM2DgOiKYmzuiKw9YFpKzCdvlwSBHuG7JaKHzSVRs9o9J49RlURF4ip6vXlkWRixl0k
pXa+5eQkopP36ozeUFF1sXr8XtezTdpkUMamLRWTNtJFdkbZYpLVzyrn9z/YoUvRUoND7S8jHSKz
9RxeXvuZSW4Kb/piIpufa2FPyeopjBasiLszaNggIaxxGrF5S6BVxYZ7yd0+ohxBdY+foHIRcFDy
xlMHHZ/QRST4ZerbW1wzDNPfyS5yfN9Zml+U0mBDYW6LLWUUiYgMsAo6lXxsnzUf+NpHdD4RbqPr
Wv12cBPq5NKBazVdaKwBS7Pov34sk5tzTer87sX6mXtUjObTZNRXIYEY6gkYfADJ8A4HXWiqKLHf
G0T+gm+zg6sJKKOUAtAuZ+rvQcDXS3akCSxdDxL7tDzddEjT6rxYUig3KGSmcC1KstyButB5g4GL
o+u3iYNFaj2MnnUo0CRz6PjXHVPxsyKkuHvXXkQkfe9OXN+nMujteQIYS9fRreznZdudesFV6AEb
xdBNbf691+vhLgZ4bb39vBBRpHd6wUxKnYMGnxzkE00kHcx1ORNlubSZxNauh6rReoxDloIgUBje
Em20cXXGVTaQzUVC7YDCO1KP4s047+AbXrEIIlvdnHnxAUfPn3fNIcG86EQ96klE8+oTRMt6fz7I
FZ22CEA0OzS6K2nC7H3OjJzfhtgFnbwNTn/hcU9qIfaP15dhs5M51cdWso9kfL+A/MzabND6PteG
6rpNMQ9iHW0ztRspoTj8nMUsRFQmQ3tWFKAY45h0FIHJAcUfBNezheitdZxkj9/EVj+qn/rngYzM
NtEm4ywvktVUSeXmH4vhrLff/XOURNurqVBKw3CLmcsBuO2/MvDQZTvW0EhylKGUEbsQd0bPztLi
fSC4xh6rvWwo8cz87Ka8T0M7n8YB6AbkKqfkzSdWQTc3/vYr4N8Lpq0uGd2+VDUDkuzqAMdWd4M1
rq4pMfHd6gQuVXvw/eu2BNUlE1LTLYGihl5icXY/8GMeJqDJHoeYTg3Aid2rxdo5MXvmLEqzBhsc
bKT6x/a8XwQNNSn1xyCT6pNlLyiKQEk91mrDhPjIX5Kt3IY8qiOuna9ccw3fl3By9nnciikjA/cA
fCEVQQRa0sunpnoavoWO3jriI/Ka7d63BYKttwmsNGPo1FFDdm5Ue0VmYr2R1+Jx2JiNFlTsMeYd
HogmlDRRIIMMayFcA+pyqGs2Hq7yoqu73KJYoA/wqcJsbRYJxiro1Zn/k4c1e2U+15gT6oQXhw8n
/u+5ai/SuIsW8hgUBd6hHVOO1jbygNrqJDCQWPsWLLIFllQyUWVb6yekQPM5TUddGRv6ovdBvtfi
xY4f6BQn0a5DMwomeHvZY7TmaJ6IDwP+0QEwxd+DDX66IPgYQsWm6xwPvXNyyIDmV+mTmyFLeC3O
euhG6STT34pS1ONwpR2jOooXYfhmT8v+eXxbu+x28GqiNHGCeBMrkFaOkI25UBJAY/uQ93XxdM3g
kXW4jcVW4APS/B9zMd7L0RPzjrxqXhdxznpLT8kB1kEOsya0nN+i1+qXSH6cPrOZSvuxdUO1uTq1
86PM7twk/EaDAGQiRM6u7+6b/0SQS9nz9ThK1Q23lLyAPqA7yDxlEIVkr6+Zkfw3ZOm6Fk8w3LYd
2hwdZPZmKy7fKIX51MCf+TPBkYCcIL5gwcWDE4Iq+g5Tfhn5v8DwA8Dyipjz0c/3XiAB1EyjPbR4
6nAU9+hMsuEUju7uKwlx9q1ai2CES81UiCPaRKSg9GYCjJiwQnhk9VDZqI+GC3JMk/TKoxg4XM0R
6F/019PT21GcJu0m6anL6cxqAzHE9TkjxHbyaE265TX+wHiFZDR9I1j8uyDxEuaHZiOwvOsoXq1/
W3/aNJaDy7Z/TneYpablz1L9cRHvSCaPjNx7oKLhp/csBshGitC6KLYN9V+wf8SyeHwtAyOOqaHW
+WSTEin8rsEhgjU4wYcC6DDtDQ5xJD2M6I5cl/Hac2g6ZMYSabXCs5gp0HF1Jlbgov1cTqoByc70
r1xKTJYbimufEgD/ZdIVcX0GziC1F/GrJuoNdqsA160yH70YMphEuWMCtVE+jTbYTJ/NEsFjmLEA
DcrXm794+GG1uuKMtz3ZqFwdccP73CRpBekaOwc7/wrKvFbmMGRCyqoSjEHAHLVkumq3/5d3u2/M
rtxJ1SJGpc4Gqzq6tfWW/k+/CF5S6egsyumkcg8d3SgKSkh+seZR0VXI3SvWBMX7S/y6pQBL1J5V
HPxmZJMpQLMTh6R6UDGPrLGM7tXfIATwuezbf8zFW+n/ztk0NFYXMKJIo7E8FSlT1zWf+IUiwM7W
tVZIaMAydolkOrhHXqvoJmSPY5NKS/DrOPqS/RY++pjeaK1t9P/39Wr/KpYXBVVa9OsDfpf2wtz7
7SG5zRqaxlrRtARZAST+s3srKcr/5t6TTj+m+Eb1UPxkpZ8dX/2LrRwHWTs4lMpNsKGgvKFLbEns
e6NluT5ws3AsGqM8xDGiBdUCZmU789iNMmZ/ivLHvNxaMnc0xUs0lLmHnakaso2RBX/u21Ir6bYX
NzaICNEniQDiRINvXVJ1l5pZFiPmY7bglLo+ygq1/T2C/YigDngDaAyzgg9zp0C1MD4ss+k9Fkgp
1jIXXxVFMZsxv1zigQl6RaqD9kWn+2xtO0FeAzojJHggj2h1WEls4HxPK/sEsRrOR7bHNk5WraYH
cj5ppCA1fQBBg3BTG1/FQfVwkTRJph49IbOK29zSGtQnKmLA27vIYsCliwft0o9v3XH8G24WOb+i
I4ZP5z04eh0jRSxm65Nhn+R0xcAVU0mZHvu6gBPX91aCwe3dDhXXMDrS38ZAYTmSr07WfKIXumIE
o0dyQoHZqtOBUZmQ5HYlmYNn529HFe80RXMigCiBX10u0Ancn9djK4zZ+YKN/9qQBku7qqY8r+HR
n74S/XZ3Eco09a/7cWk6I7jROiLDYN6KrEM/BM/laGtNMsNUlhlyyTeeJbaMIhgRll10eg0w0sHw
5w5ODgRfmG/gedB/sWx45X3EKSe78p9L6F3UgWD3kRdnhQb+XNDdHrbH/E3EgDAqUI6vHpCJGj7Z
jl+4IVRZRV3ANhgbSMoLc3D48DYRAOkYaz5NSVBlZbOQ9Ju3vehzSz0mkV8zIXX9u3HC9QEz/c72
y7swDCY4lU/BL7U+gqUV+ezmd0A6j8ctE7XaoeDJKoPmN/geu899kjfs9WKWEXUJvddQIcUI5wTT
EKdaNKzrYZgt+BH3z2LbWTjto0x99fFmW0YD8JVa2Mmf3kSUf7npv2MMg1Yt4qV1Eb7/26VfTEBl
zXTIv1QcwKJHJ3YEtMgdmZFjFjLiVzE8C76kuNRIkV8YJQ2ZbEQZQJeUkYGeTZuqqGYqq84lU+5C
bJ+UDoRA6cU8CFf9Oh+Y0uLz6nVXbo8cJPrzYWO8pKNd64EN7vyaCqd1rt2lMUUZEyYT80r4DfLi
VwLHJ+iBDh8vIZoNzKUj4O2uAfUWufVJp5fvksDqopnKjQGkJyHYhb7G3DqlpG3T2TTI4f+v+jqq
s3XZpjvL3sMRp/Pnwu9R1OBCAWWCfiS3YlqCGaeOzh588Y9WeMxxv42J/2CDWz659BP6wGI9p5Vd
Z7GEoWZ/b0t+j3WN7ToNi+ZIq97nVZtRsyQadXyboh7mdvqtMetTP3eo6C/EEkHXc59Ht5CTzY9G
Y+1Bx7zHTsL3x3c50kpG2nNCtqMPrV36N292WpoxWUWESEsCAVnTKPtsV2LtTlG7WKuGh78vyJ5W
n2hzs9dEwwyZDPMTT9b+v+Z8lesn+gebd7X5IiX/fvqY7cSBpr4xZwJzRR+TLNKEEQzciqVF/XlW
Fze/1mJRRCzuOcxIouRjjyEqH6SWcNWNFZd0Vh+236oqT4+i0titG0Addd1aDWQpiFAsTEB3CLch
VOJ4ubcBTYbuCcmQfc9+K9qLaWyG4D9Y9HbTrCKAGyrCaxuKmqSX+CQehwADg1ntR/+N/ZbtmD1T
g4PAnmUA2j3cQKH/wRJMdxMZSsFYZ0QPQCSdondyyj1Jyo7CTOXZHtJAdvJ80kL98KUyI8jlHs9q
3td3dd2eoKGOPrkiVQvzjmxIxAXxShAsWA5/uIevNF3yAYkSIACUbPcba3b7RVG3iK0MJgDznPc/
s7ekUL4QmoC0cQ+WO9gwEfoYwy2WO7m0wwO2VPZ+jkNb2Ykzmc+5weUlWfgL9IZLvV3rwQ7HTobg
nSeEoM4US/rDfoJlM+ztbPq/wcQKp4vEl1ij5gUj0VSaWuEF+tlfLvda2YNkvskP1nCCxH7og7pt
sRzTjC23GVHm7G+XOxnr1IPC0GXeuD/5ESyRoGW50JNlMk6V9lp0C945D+Om7NmjrX1yZEk55KZr
k7f6gd5Ty5hwvWOtLFqQcQjZFev3bhljNsHSrxJTxl66smDOgMfs50smRASSuJotfghR7pfAi/Sq
OEo3JQaQ+5+10Ej1PG73BDeQDV0kwu5J+YY+CevNs8yuRg8l/+zuX2XaqzWxUUobnaWHTCXIv83u
FiSxnNUqViPwHdDuJTkiEt54PaNi2dPK5kFYZVzw0P9jr3ZY0q9sLRKcWJ01/+ADN3DpMCi+zZ2f
ppyfPUZNnK1rBOEbUs+pBvXr4ZdXk9x+AOazqXmGA49fI3ppSZ1bu4ZFQv09+fpidtbrXWKCi3Xj
pZhKQBv20ItYwGCQv66Z6lvgFFKzAZFmxTTE6kdGPoqh0Vw5XsqrSCUCb3+cWDL3Ein2NlCDg90Z
VmZvGfDXCl1eHMbidL8z6sJVOT4EVoQbmfWBDz57+FRZ09+fW/4lLbKgYV3h+gUwMnE4KoD3azVc
r/D7TNM2F9M1YKOOGxnT/ejKRr8YEOuAdmMJlqnCIoOA4gBc0x2lKuSKy9ro1QpQgDCRm9yIz8if
VkZnTBARarcGvYMc6L8Tdu06znKEb3+gojuIrX4XIhZWIqBpDtyZ3St7jPMIiCpnvL0GcKRgliUp
aaw2Oym7GjKK7rmvxUiS4ONv3/ny984SQP2ssatBEI5+wVsGDYFrPdt7V11E1cTz/gIQqgeqkc20
qhwWMOivG9VSmMhgiw3K8xB7r/uKdf3fsVVtxGZqoY+Lt/mx9mzIn3tP7hqcBg4fSNB+VVxzLr8i
fm1TAOnc3kNVIZ6c7TMTkv2OY4XUeTDQUe0IliI41y/V0mVgmCnRhAa4OsV8s4F46R5qKE097fSM
WHMCENXPPFC9NZH7PWuIJrL7JaMLHImj3NzvUcTL6Kkwe5SzLjpz+NUb5i8wlQYzHqO6nQTsbAZb
YqZMYcyTe52ptH1+VLdxMjDSLc3ULIeDwM2OZJbXUMvwCSTkH14KYmGMhULmJnlKplJUKtDPC4Sy
acE5pyuWN0FcRMApjnGKT0/teohLQT/N1oe1/o7iKywaOrFGu/82IAzAiGfoM6sFI0e69e3I0geN
7C+G0wrgV/jS9/eK1fVj5/Fg8NkDhFBbBQ8AcSqE48tVHvcImxygGisJhajpZfeuvCHraEr8DuuJ
EBnQ6EBaqa8JjURzgv5E5S6bZLw54NgItiXMcljNA5+4C7w28myM1C9czhsnSVq4u/v88FxEOE6U
AXhIVXuI4FZ0YknhTqmiW5kIGTphveybAyZhLveV15OT401ISDkhVyM7QHrdVeKuk83UzNxyV/Lf
kEsN6js/tUm0lUqZrx3KJ/DBNhhNRMVoSiyK35joct/rCCqZxazqAsHqoOiSxk5+gYBQ9Pc9edm3
b2/mFPdZN1iYJCndza8k1yrPXDZExPS6J5F9gBc+sW5Ik06TrP50ZAmLvmB7A5ccZO0slAHKmtaE
XNqsnADxJbN0r6q7X044Q1QGzyjMKzkNuzX+kLcmhHOaaYzZ6CRk7wly+0W+R87aJELwoPwQg38C
zvPhhGMQkFNCMJpT0uqHe5rf7Leh3Rw0v04l2m6AzoOadGvdsTm7xudTP26QDU+agXKRlv/htOqP
xRfcR/i/vo8k1EibYvwAKGqo+MirUQ/5QTICoob87lUNq9r1ZdglGhRapp5u8noeIlpaRVJ/P5dE
bSn6523umwbuEgkGTuodZEEGqHG78zI/HZBbps2m+5tRigYmeKS25EWxxMFM5xY9qBNL6yDG2Pvx
Zs4eLZX/BeOoN9g8tPzGT6LJQTh/uFGeQZxoAv14yX/squ5DhMERUQW+87QW22L2Uv3/keoOLIVT
oc0BtrtnZ6WQoCUFAaOJHU5xBzFFC3snrsa3OrLdroAT8iXVJ7RbWLvmX8kPdzmrtLd/fkatLStg
EZSyAf7glzhHDxCA/KpcB8yeAJVv3v8zvzPqKCRSoB0O1JkXykprisZ5i1omjaWwtqqQmk5KdyAZ
ZHykrl3Q0t2RqfIdiudVbUtCBN+xzKcyv4cUfqUlnzNQCztpvRnxWM4iwj/M4c95q3MIaL1SF435
brF3e2BwirgvkSgSvDVWAwmlADqu1TR3641nrMQvMiD5Di3srSH5q90qP+7wIvL2MVfB+Zo9e9Zs
Zhqi4Z2Snq577GuD1X8G47nf+0wB4nx8qXowjfiT5tLW/Kkhy4eMVgvppZssnWh9/GliOTofYx0v
F/2LfIEKJXHenx2U70lt8sLNhsZJ8tYTeG7BCS075p/YIpITfmAZLgMczStRA33w6Vnr8HYaDGwc
TT+441QHueNkPjUqI6tH1pG4OsnyEsph3PbBW+/fmGPgQfgepV+xn3cWNo5xGQovQXELnYq4Q5c5
7fC6ObZwm8UGA09CTunf9C4YNki5Pf1Gkb2ct5YNp6vmvuZVWXGT4s9SRP0Vd4rIWDZpU3TeON9H
Xcro6MbngNxF+90xLEwOnxv7ut90wXFfDgoosQT+bed1uRNJuNnKiI/BTquTdhpO/jmdQbiOs4Z+
7S1lYoQw/b4RdUhI9Wk8MLt+RomO8pJ7k+stBP5Xw6wTeGr2Rhi6epHhwnuW/o1LjR4r/1SLFE+G
r64Z93i2+1wuI6duyoOme0EbtlqLd4wBhxazH1Z4VLDhxy3eXlXT++uulzOFju0Nfm5vV8BD01Wx
N3GnYUtyy/W9o8HOJb8dyKyaopTFOH86G3OAsLdHC6CVZ6cA+uK3+U59HzBB3BVDRToVtnpq9sGd
7k21TkD2pQ428R/zVOilkf0eMJzb2TNTRCYpejF7yncg6hQ61plQoAMvC9gtHJ7ac4C5WLJlwmru
3R5NNgOC4JQrENg9b0MtK4YQeEG/sRwaZXYmRr6cr6f8JFniTpPbCNARensDtslNTQIbYkeFVMl2
5DJ3aQOAEqjoQcMAH33ibSI6zFPSboG2Ze91BqVMIw4BVnsYGYzEw6EVCJiXoYF5linUUOyVYpOD
gC/K1OtF2ER+hmrnhGrgFQNQ+MYWjyLL1a7e3tCE70nGfeJisrPiMYr7lBaODRYNmMIw1C6ngZpN
3hS/5euTA7uj3TuvqohNXJz6uY6tRCnBj5Ue9AT4PPvPkZVhSPWrFvfp/JQInHLEQpWikeYEcOHG
TcXBolCM1itv1twyGBF4gkdYSlGD0xFNclyya6ztwsNh7YenpQB9quYWgDSishVhd6hoS0n8D5Xr
6zFDj79OnvE/oLuWzxVXpms39fzU/ehXFAf7K3B8OgTtfgcQario4sXIgZmMXioLBj8/l0eeFQDB
s6hjnNUcGZMQCOWQE6bFKBvGNSgFL0NMYTbUYmIraNFqNpvc+65DL7lRuKlqNSQsORtQNNJphtT3
4bwkjxCPCQDloLzmmsQzbCDMb0ItW8WJsmArYWE5nRbw6GcBDtiIHKwuI8wCLlUw5EqMuNDqoB7G
aAadtZNBhlRUcxwLYCzgNJIzUEiXLRzoMVxG60oENL6mN8ufVkdKM/hHsMFC0l78IRj6Jdsh0NjW
o6Q0Bp8PRfNw+bC5HVLsn6ar3Z2EoJmaYVzaOyHpDwE9HOoYVgp6pLl7JW9SMiC4XAwq8578nUjd
K/t2NOtzAOIdMDUlQ0HKYSUBSvMTBH3ReZoHB02whzciQ3oBNFfPbEZJD4pGBzUggDeWLVtwdCNW
Jwbd0SuEb4KyadT8ABdLoAsduDYOY7MVyUsjJOEmY+ReW8yCIANQjXetYIvWKP/6BuaOP/Fm/Q8t
ra0jeVZPANKbZNkKPCoJ1dHpvfV+Y+mT/1l9HS86qdftqO35qRv1HZqII+T/H7kkJAKf3LjPPAmj
tJ7lOT6IeFCxlwuWlBoYRZRlFTlTh8DKp7FIbrAvgzbUIOqtKp4COJuyd6TFAhr7G/N8x2ywcxol
Ku1G8OZ8ATQri+M6fM/9KVEQ8V1o8h9s84h77R0HCNnMT6jsTkN+KjUtfS7sA464yZrsy2IWuJJ+
R82HiGlE0QmsJSdVgu1l0elcJPulA6sNABGNtisD9VsZuPHxCSCEzX0JoP2SIhoHFkJ0CjQOyqIN
cWDgR4wskH4wCK7muwhs+H8QYoEUhx8BrxhY4NSRNgobAqTilzVfncytt8im5tMFJFBbhslr/c1f
zpxfR+WLKFb+M+kTrzFkh6dvmXwqZaZLRZvfJVG9yhduBTxPh8Q8jgmE1jUtDqjmZIZgsi+VxQmz
h16rcD/LAkKKPZRkyGkSxTOiAUA98MlfB+OpFO4KfQthWQJWflzj+MV3598MaiGb5d9JLrLYsxoR
vnp1Kr96cqyUIGiYb5U8wOkCTxAfukgWTlC9kwMZI6OzGZ7kFLy7Vy/4gXweIHZwY0EuymhTxisE
+qH07x5Tzq6CuudQJEYw6RGJ25OL7suQw/h5BbHx9AT3qMRv0Qdyo0M0FcO9K/fboezh8RaEbHiV
3qMSq5EKyFj8P/99lqflNFUbU2Wd2MV+D+3wEuzfnitGJjLpQC2CDEcbHzLmK/QGp/4MZqwKBtBv
YUVSxAfkjZKSmfPDFlJzXWOuxmBD5mQo23GsMM2qLptPfXToxoZJQ1kOtqCY1iwDAiayS1S1H3CX
a6NB5NvduCo+RAyTszLSLwGzPmfd67LoulCkZh41PvgBqVwPdOCEABcdDqR81LiYamrwyFDdoLrc
MJrARpUoAsCQ2YtzUKMVrFtllsHXfTzuT76SKy5bYgkm4Z9vhQda8XHz8uvp3DPN9vNjRJwLcXUf
zBBkRzbfex4cL9zBdoQTDHIFAUtsBiGjI4WQTMjnP4gpNyZ61ZXj+wO56gb26ouPY8xv2BLdM8L+
qMKVjC3K0RHz5mfp19IczIeUBkpoE0f65ybZkLOJ/A3EA19odY6adqYYg18v9BVEjkIiTZW9Entb
lOMoNBy0Y9EEUnCGlZshT1Vy1wDv0PxSZWJXmdPHWwJPv+pvYcMWKe7dBXAfFfQATSBt+Wi4Soo7
xvHukbSQPlHr9uyVE8cgjLZ8RfR+aDtJDwT1869gz+Kr9y7IdKMJUwyof2/EWMHjh7ef3c6nXoZG
Q0WQlWOQDORcZQZEwqHuN1nD16i3myF58DBwAy5vmgq1zFfXQOhp+8W9pu8F0hVrNntjpo3D2MNq
0rnYCgsPsLrluiQejVQaBlVS5/SoPtQxkQrUot04/O+pk4svp22KZ5itvNNiIO8ruEXvFbgdn+4o
BJiJz+IWUxpontOUPLbc2acA6yf0VI4K1hoMWloTnce7LDSwTEtAbxxDcD09AkBYQv8xRzH9NqFt
3xdlEgbE2tQ4HW4D1iD2g0dGosukVhIXerMuZU2zudJjdnDrN/2RqmeNMKqC6SCpujNOdiA4maH4
q8Mv4DZve+pcbhOHqe3ZPZ3biG1O0prsNiOD39jlTGIpGN1owpwINueQ5Cq2TGJuN6HVA9etjfKF
hU5Jm04677m6mCgXcuU6Cxm2s4CvMfFq4ali3RMhHTAgLBZUcs9wrU5oJe7HORfnfdexbwVwDgca
aXzZGePV4WrqnCUDMdIMVC4KZKZHkHB3eXFSpxuEbgMvwlkTxDhR2biaOhgbq54LPCNzuEwEEnhR
Mvl5ulZK0pBvuw61DbTkKkYMQkAsFrJUPapb9VoE7ey9wq60t/xNSfTyJvQ+qQHOveUOgw80mu28
2zffCe1+9RLVfc3RqeubbzkxnMhYbVG0hQPgCtDUVdhUxxmsXWg3NUJuAHOigNIxc/rJnHQz+G8V
sOF0Wk5ga+m6/XLGo6Xicak1lws6frc4ouyNEEha+V85aAZhA3yI7tb2eWVxWa7Hs+647T2Oymeo
BHvnfpBl1URD0TgnOxk0pRCkN07VaMaAYjdas67VScRJcAg/hsJqnNx/2/axWay1UGtN5+qw82/i
FuPG65G3kyHIMTt5SpV7SwYnjIwv1XKgAAJdfCLnkUyewQUCVIBm6G4Tu/rU4hy1kkO18SZjaIyr
HA/zaChz7B3Da8+ZliTUX44MRMTaCIgOrKcI7gg30lNaMSK2KCjK8e+MP3YzaDqItBOLbm+08Il8
ATYRC7ExIx2Yt0MCppykDP7n5TXteEyeag4kNS1fc/8mWXN544axG549w/W24ikmH3qemDfPuF0G
WCdCwxmcQ7SrFwPylJsDRBcUrzRdm8z9YAv1XusBfJ8/Sw9sB8PJWuKElVgGGUOvyZt9WIVAEV0a
EPkdvKoJFW2InIPZ9TrxE6Mc3MdGACks0B/7F0OV28nASZDXxaDeIVTQnAFszx1Q7UltDlkW8lEh
imn3kKgD2GCi3sgTVwo8pfAaXooyJt8f+ijRAe4dxJxccCuKKaDE28JryVPTHIl8XgjkBb0IfBHz
SpSrBvOHSQu/Q2kANQtLs+ln3C/GaHe8cT/Go3nRfhkP3Y0P1vCw92MlY1ZTLAA7QvPMrb+MesRy
YVn/3fwq5E6cIA4uo6RtTKSvKPROjRQU/4C/eLPg+LE5L6+mPzNe6CrQcjfe5StkPRD3rdvCdP1p
yPBTdUBJmOUgzQgi+Ynv5yKyT+ev5yVb53fx+sWQSu6CZo85QAv02ycJcXu0pOWYfOn0gmXQtN/3
NdpAKVEkVJ22i8QWdqegOwafK2zp8Wh765toT7Bd6o1kfBGAi+fVA7OMRnI6dykN//TEjr9f899I
jG9T+i/ll4q1M5L/41hmflmXN7adNkoY0jr35gu2nlaPp+4Mx6JJZwZpdfY0G1WIJQNviLbFiG9Q
2Q1HEiOK+ezrqQcf9Ie/lTKyU4L8rp/G3GSx07fqKwqyvBGsfTbnnV5qEc5XkJcA8l7WGqTcIlT6
Rn5FjKZcV4jbHNQVwbPKrSfUMlmngrYBhez84GoUDo3T7+Q3jnv7j62VAuRURM5Vkih/bNMd+aQv
fENXCjKf3SNZWXtqzxYNq8mNpVQIEUgRxU3VKbxcYOGhktQEnSJOHDrHtfDBP3OKJAN5Uj35UIqy
p8cPiv9F+Jn462xOHOEWyJI6Kr+UXKkk2R7gt0kXYdFUwFPbX159XqXWnhqyyjLA62DRRDHNBXtt
SdzkDOT6bNpQF6Hno4cdaTIcmujyvXJmz+49KXXccrK1uWQV9hWXfXr5BbKzGBKLRUwYteupRVq4
vwHKQS6kJ+BBd9QluzwFw6IPbc7YAZed/vt81/WIAcie7XnagzgP01w0w3WZ6Ow0I5fuxj3YQsWX
sesnOQiWztEQsBu6944Uz0erb9ysF/N6Ca90C2Gf7ooPoHLTYVEm9udmB0p1+RmxgmpS0A4CHvVl
7IPeemPkEhjiLtffvQo6Z2ct3sQBCd3ZLRco1eRVZsE0q+hsYCP4yFbKMOJPTFWx3xOlDJT/B9QN
WeqXGLvyI9R3KisvH9/MkG8Z4VcNn35eGETe5R91s4ngZuI2eMJ9B/DO6AMq1wlxJU2xxOoS+N7o
Unf9x91IGq9H6haxD3S8U7C70yOa20OrbiiqCj7Phtvc2/HrBxXZONPJIaK81NDzqSJ+3c2qUP8l
pKu7Q2GA0qIRN4BcZhUNNgKA6YEHhbg0Izsw6npZBEjvTWZP50NtGvOIhcVBQB83vTR1Gi1BBlo8
3aojmcXR9mO1xJw/NiJNdnx2gOkLmqfIVHsa3JyLZmvCF5q6pSzBRdAoBD8YtZcW92DXKWMVXAjH
Qo0FKx4Nz0X8UEDrexiIogQnSerx30YGtBpGIYJc2w8ob0nhBo4n3UfVdfYpgHSEDQJ6QHPP5z2I
1u3/nODLzaUgj80kkb/5nBmmydnUAITTsBp6YQ3LnqPMSLmQspTqPgX7xy7wJaYCv8FGsCl8lUsF
wjNLgTZyiwA0SJDB0WOsn7gocDfFJRPTqDVA/JVAODiDx/scUt+3KrMTElgt4UPvMymJCwac9P+E
QUxWE3TOyCfzpM8u1juTO2sIq6djy91EFyN1wJ9YUtMhFKY1FqmbWpEji5RsVN8PVb9IZHJ1JOAm
ckPcD+MKVUHOhF9ybvvXIhSmKe5eKyyZWbmpzGFD1/X23Q1cToVafF/AdXpmBzDNJOU5obWL5F9s
yETg3eZ+lzmuNkKFfN8+s6VFVFO4V2WcVojxpHZPilWva0EDJsHtj3DUGeBU6BhHhtYVVUNAqlJL
UxSuVYLi8fYAiFgYuI1TCYY6Ueq6ektmding/Nqi/NxRd8dtT6cgVc5RNXBDCYMzM5JSDefoFY2j
N7TDt+Ur9pRrUNajHFicq8lorLtnbY+NxESAAsOMl7GypZeef7MCMClPQQeHb3cA1WCqCaVRF/cx
5kY5n+5gkN4ZAi6GnZV04Q/VevorUd/CRf3PSr3jROrSh/HDoMz3O9qRPnJqMn5rEFZrwI9bFP1o
3qmUSr4OuSPbTPjhy52TmVdRSWy0aubD77BZOMh514ifThyuW0HK+9jrwJAwCNrJMNm/HUawMx4M
6HvPSwu7OddDRYSEd7Cue3lcAzwM/zGb3Emy9/cLcpgzsGEPxDqtOcLbqCqu6BLJPnaXs9XUW+Jw
Si+164RJCsPE+N13ELJPT4eX3fPUKomoCc43glxS/AXBewo8fZU4EbMxIphDnkrKzva1i3bR7UfF
sGAVrdCUitHeBJATIZPX/+JcIkahCK3gTlEVRs4vetI6oQ1axaJ6UtuSUTFaEK/WpSjmtCFMs3yy
p+H6WKuL199gzHGhaHWW8kHGpwLA+oIJ0Pl6azNJrgt2z3wb3ky0BJoSTG9NOffnVp5ohUICywhU
vneP8IL0Wr0K0tHW8HRkOCC0PwmvozTPDVgRwn7C31uwJC67xgidjCI2g4FTbec9ewqFhPP1foa1
DbnM8fhq36gMFGC0Ch1ifWwNWrdY8+ppOijSqH8p6OhIYPlCQZdMVu5aX0jK2ewfFzWvTi5bEtGW
L1ATA7uso5w9i2JMnAckfnTKFpCOpEp2ESJSyoCcVkhhmRwa1w4gjURxF5xR3B9hJ+3C+IixEE1Q
0Q/wuLYOMP4hn/hNeX710WLkgol0BdgizQIdzArKxiDOEQrSq7TompBIetMqF3pXn7uh/338TC5k
aVPpHslJWNlP8jSo+16nGfKbncxcgr30BDNQ/eBjgGpUdldAre+2zIlBOtcIww0CArtHyx2BLsN6
ONKBxoTQmv5Vb5HeFvVTLsjzSaFXpxbiFaxYPBb0Rvhny6H9A0ETt6hGULb3DJnDRPN+7sS2tHLL
+PzFR076CG2JYLIWE2Awul62koabtJIgo9Xp+nZMT0SBfglHd3OMUtbEJ63qcI6+3xbxNYfKZNCw
SmuNb48PhMJ8GPqc9G7/ig4OlYdSQSWt6fM4ER4SEhkTb+DZaXmwMyTD794Ui9H4gdBzdNBFwvY0
cbuLhm9Ie7N9ExzjO/NuJ0IBWg4oWIvSaJrim0tyxtDUoRWBrcrwYr0QuXcFphQFEGYFP9dGrL8u
JPFv79FYUngwmnlzx7KmCLohvSB7uoqEefe5v0UlTWFRniZO7BmsvmExepmGSzj3+jGY0Kl4+kh7
/+kjNDFsF35NGzh1Zb8v0AzHJ2LxqN37q6wKeYYMR/9NNb7yyYk1JIBFwUd82gfa3RmdHr5PZibf
shuBquP2WgWFSz01uCFwHW15Pbb0OgjBNcs/7Bss7C9zV1uMAGnZqgSuREfq+xAvlUQvH7Ff0NUR
kpuKD7k6cGRQJAITlxqR7PMq4CNykAMvPw4jU025739i2iALyT79agCD49eHVMKGKCkd3GCU2PKa
i7idsJnF+NN0EMv1hX3X7gBZbiZ0rKDCVCnOnx7ugadIDDgdcZYtk56Jbf0pQFKmtfcMphtWQ5uc
jZkYPljfvQdFfxaK/hKdHP2W8jRSsCPE5FidlUnI599OXHC0XXEaqx+N9WxGTuGFF0fet/f8Y5oq
oNYqKJg52BKSjJBKRUZ500vnl2iaoBGtnKU/8aUijlLL/tZzzKv+b1s6DSgGR30mObqwvMZYnMLW
XCVpBzinHatQVyZAsIJ5IqvgabgVcuP68A2PfJvy8EL3aPBESm0nNOwvic33eoeoVXNAQJjpzX7r
40uZC6pOXyIRo3wrU0U8KAFMNhg5u5PRDDEM8ZmK21cySYx2FNei1IeYO7TeZyPJM71LQqTLaYQe
9eHIc0wvbzE02knZhJNlCw/NSsKGhAJw1Q++5mtMnVCQEMmHm+Ownrv0OAynflc/XsMsE54WoKVl
PPoFAnjlI1MDeqMBdapyTmhThLpGN0IS4q8YI4TExBLSfwq2xR2YG2CtUr+u5ZsCOUFphmCDW2nQ
6PETI/bZfhOpyMntUyDDDCTesgyJpLnHeVS6dJYgC1oLCvVCHYNgJh1exiPq3gIYCmtY5GfZVsCu
DFzCWaQSZr/tFTqgkWOovB4R/LRfXKCZeGcwjIsWxm+a5pG2Kkb5dcxw3/WWRxMy4OigwhwewDyC
64vpzF2pzLUo3eFVB8fOSy7y3yefu+89u4Yf7pqqiJb3jtQ+pSUoQux4dXysL8Yibn+Hgw/hOsJM
XN/tW5L6MoDlWWodpYhgv/nnTlWlPGbeg7OfuSQ0YPdZXO+fxqx98Xem16QsUDBp0Twf8a4FWzdF
+RAi0vpq1ZYVwyWzwjuOJkN1RJ1JQu5BdUks/3DOgZygwTObA8JzBZpfl4NFXe6Rn6Q9t7K67pF3
/4Ht+SMSQX0an3ch+p8WIi5ZhUpJjtsYdrPagnN8CcFUOwtn4Fhu4+WNX8y0twpYA/WlTuXTJRLJ
kEbmintTX1DPKxBkPlR88SMKFvOCFHzHC9+vfox91A7HH5OybPbT0cnspGIzFRCxySjdY+5/eJ3J
mcWa6lBMe3F9vR94NVDqZYsqVU/7kZr66L6rPLL3Ea86KId1mQyMx6vWNRLY0G6qe7UmxC8Gx/FS
rxPhZ0kyTzFFxYMNp+5y+Z1x1DaTgVyg8mQygUwW21EHUTUeJluRmzHMR7/9Y4306IcoXiJJUxnd
IixcVQW5R8Dp0fIb7l+yReBr0yFo5Qp4Jf+u+zBhsIxOW3i4MKO7YoTX/xh2Xuf15Lq35WpSz5pM
MvNlH3ZVwJlWU+xw9XokWDwZ1aEBJ30gtqJ74KUSeQpaImQqaqulztCctZhifitYNieUprp5q3Pe
YQaoHs1rgDVJYYBXSGtQrOcVwIs4sDj059EHKtho2ODz3YYIVY+uZoC8o8oDdJF+ZsL3lo2Nh9CO
kkUamY4XqSFFoq8bh0OyH6yxd0ZzSoQrultC5pUhcBQpxrRSlUJteJt0JJyb+k27NNUeMUaXapNL
6ytcJ8N/cLrT+zlE0jmbk8yvnbGWtuYq028KWdIUQ6sqak0yLHbVHnHSrwiRLR6F0kpPzRzGNgOO
/stUX26uVpUPGeNCoXUXRbmvxjPiELKJ1G2/x/UPyAzyJx06grzAFfkNngDpt7ICec0zMm1+olDr
MogS4UMl37eKF1BPBv4MBIVrOaJq1ucXZunyTgtkmxbYgpxiw+7F9nI4OedSNs9G0MqjM4ZFkEOI
9gbF3ewHnoHJDAvcCSuv5xsUbsEamruVBuR1bCWxLAnwef4Lvkq6zhpePVYPPwOz1n7FUBaOOqEx
qnCMWD+ljajpf/+Z1hfm6s7WC3OtF1CrC4vNfQ4ah3YjF8Nfy7sWLy1jUVX0gNiiEBYLYdzJuHVw
i+naV3DNhTbOttwJPhKSI4Bik+GkKxJH5jEnP2RkRS3J9Le6JuO268FYiF8GzQN3Yx8Ol8Bcnp7W
wee9HsabuVUAC+yv499fk8Qe9z25j+10A3X0DDDV2oObXgRGIEm32QUdeOm5N82dJKJ0hPM59Viz
/U03P67NB6k4quhXFJ+ZO/1aVluAzbW8n4pZCJvdgUYHVjUtaUJ+V9Aj9HmWHLN56cznp0A4WcIW
uSqEM3678tRSlvNEkRyW/2nmLTNC5edT4+ju9ANdwV/dG83LpccZRWTW0X2khwOOB+3Zx8ksSrvy
3v48NtXViK3YPc8RfBHtnPV3+OMTtnR26nWYxidg3YgrKQjGxMwaVABk4qkxXTkztkbpl9/6aqar
Obc/BevytRxLjUrkcJHZiG4+7FjdH6qzCsyfYK4UO5M96+jae/CR2/+7HASjoIGk1Mz0UHQioldE
OfTV+zJ7XeTbckXXsvCf+6S/zTnDsRCsfs0SLrjChdN3tHrgPlJZC7alyeTaSz96H7m2M278Uwsh
wtgg6lLJP+lh/nWeuGAqTh7ddYYN08x2moSg4jl2DmILY/CY0pmxW4ed300YT6MN58Zc882gRvck
whFNdbgIb2Q18Y7QOiPNuguVr61rK6+MZ9xMbqbOiSIOL6AGgO8ZiKd1GfOECsM+cfF4Na2PBKy6
mt/4kCNBO+nfgNLKZaxWIocenlI2+FtphOs3IHaO9MxtQS9rDbF/XomVk2jqvFqoqTN1TlLmMITX
g+0P1Q7x7/DYH3DEoIo0RyVy7CeAYrK/7PFfritwiVje+4nrIbJCGoUTnBWl06lshcDtz/ytyOt1
24n7OJMOYK+NvLUexCF/3yOc4IkcbQs0MOvfrPFKAIIO+2oHlf9h9PbYvUD7AT0kjE0JsVBCsNcq
xjJsUKL2OP1V/QjI6WptgBfYJRUXLlmKtfAMRi3SuPIxCbQK2XGhQUmk9DyW/3sD0rJ8hN81MkE4
picE0449ZMuhP1onTLo4AJ8xVtPbyZsisJvVo72SJSzSR0ODyfG+IaMrpfGBlPr9Ow2wqf6BbE1Q
/Xn6Yc8LUOwHnQ7NMIj3i/FtSCd+JYcxWPkrwR3GqjDyO7avPixi/K/dFDCO7dO5tnoKoYcBLNEx
evoeIaDqHce6cY7b5OlaY6hWtElxG+G/0TLYtV8ACVSQwYdCjU42W9Yt4dsPNm4QyKu7XVuWXnm3
XL+UqG6HXpK8ZsFDVgvMmXsh7tVCPO44n01DiIZXVZvhwmnyif+ZtrmWuHcy7PWaSKy+u8seMQrl
jJrunKlw7dML59yasbk4FPFVczh9wb2fm0nIh/x7kJvHdq2IWL7os3vGKsoFXsRE5fIxw3+t4RPh
64BsVAKdFkFKe206aRjRH2ZoaYn8s5qFIOLLY/9UKR3D4uUGqfCpmTv5dDEFPOBFp3096BviXhw7
57i8/T8LdNjZ2Q5Ax+Qqo9G7b/oKAUJL5wfQce3meY5faMWELK/3OpNxHmsHtdH6gXI4Ge/kMCdV
2SwCHP0AayRjpBNCpB3xmA4+473G9i2UNd/RT55oTINHaMwxVaalUu7DJZUAbUghtSmKOpavs0dz
zbcDuLvDmz9MoUI05DeEv392WgVw34feE3n1favtupYDyLGsnNBAaQi74YKazLe2bMUBeo5PwxG0
+2wG+v6EcHCIqdR/BtFtgSjxFL3Foy+G9bY2Wk/U66eZu5s0q1CADLvXlxEjxzjjlWdPvEWzHi58
KNzOtmxmo8/vzn+Lo7KJSWYPxwmruIokgJJPnLaZwfJu8x9r/sTxklPQ5WbsF22VlpMhkOh2Q+Z8
h6JTbqWDcJh6cItS64nKfUEhBigNPpSNcQOiwKsB4GsNvBAZSOca16o4IpsJ/te7/iMi9uA+db8K
8JJuSZDgxDjQZHh3iwvJ1+/QNrFIa5LutHzOHbJ1oX94/KEcXqSWk7ivX5Z1lPhITClR9fiMMaRC
9eB77pj4yui0HucLQqVGMuzneU8ttIHTnDut63saVEI0Ay27oiLqckmpNmU8D1yL67NJPHh2g4LA
IoSPlVOKE4j0tQigPOsKFkiaZghqM1dyU1sbbp19buLoBNgYTKsKjHwAxEzze82SXSwTpufiDFqL
lVVIDC52zJ3vuuO6wU5HxObvFIyrXmTF0e1j6UaScOUhVlCpWA4W24bxlq7WpeatDGr7fz3lo7rL
472jenWaPLemr6QI4HRMI5hXIgIMm20MHXvxcAz6iZHaHAaXqTg40wrtK2s4B9nKGktWDhjh9CDl
fDAOvlc1N49FWlml1VlqeZg9gmmKRvyjFQjAsNI2XOn+QRB0yIAAHbmu4RJDCn2VshY3/Ym13TLm
pF4UUc1B6cF+osjwWwmlF4wJ8aSgLL7VO3rUGrX90ZwRLhANajUFV4LHGdoe18W0D2pWXOT+fXde
8hJv3XwrKI0dM0ROPOdve/r200pqsNObxYohRfglD2T+roZHg2DDJ3mso6xJ4MNfHyB+8pyFHZr5
AvRDcallgQDJOKtE/OzSj9D6NLk/eh+GSzOTBbYXIim4rVSUZd/hMNRCTfr27u7OwDaX4u2cjvBk
tdF6+aHkB66aK2EyRovhyn/xmMwiC9GKZ0qI/0+bFoLSeUW6YiJYE9M8ZFYvV3L9Dzm5FA5RoMa3
mLuUHOUg4YBxn/0qaa1wSqwz4sptqobc/y92ewF3pJy9zWt0FUZdy0f3cpz0OHE094W2kDx4xchL
jbdAYOQUzi9BQbwUwm3OFeRShMh6RK5M0NE+1GF/EjxzFIAIQXGHGpxSdiUGrSwHSIaP0cv2OJX/
HUUdL8+X6gSSwMSVRkKVAxx1Pl7M29U43dEi9Fb7hvMUTbMjJ61pApdIR+W8PNYCTEtJwDMs8Mkf
CLHrReSvIGBGK5TIdhIRaQV76hkwK4VC/Zhh9pdjl8e+UnDmL81GWMqpuVHkpa1ceXl6uOv0e5e0
uR5LgqPwl4IFeryHY9qjjmdsMs6KSpAO/x0yIF7pYTz++JrsX6q5N7N07SKe5HIJr8d7s8tN7Cqt
MOG+L8/OJRwTVB2/X0taiQ/E2wMyfpyZesk8vVa9oaXUJUCXIhLMEFvnsoOlM04oTP8+OLEBcKIZ
W2I+p1HA1NIeU9f2lhjwsoUTJrUl/A++TCiz21xsDRxIHJLCBrCrJ+TBWgt4+cvJUSrMZOlbprb8
uckkqeU3JkPHYarTL6//mUgFAme/rvlaWdydfcDBIcSJErLmrcnGqEEGlPByg2u37kuA8QfgWmIW
HqN8+xda2nG8HjTfKGvemBog5M2OD1k93qPaz5KXpN2jGw8xcf6w8tukcjWN5HLJWVXPPoG5raC6
9LiDKnPA9IRD7aLJEI/HavJAWfni5Po+wvKMiPUAmioxeDdefQnH4leUp1bn4m8ei38l8yBOKm9L
rQ5q3vofHwUJnXVFv7F22Fgvk4xyIn0qJff5CwqW0amH3b8k79Yhf/sOmkOD7aRWk1prbffYHYFZ
Ba2PrGMrO81Rop3hBVp50GpdzEWEjX9d5lbFileDlZNwo4IcFclgYlxuRruFqP8u7Krsoe9fJVXW
euUCreOdL1I/156bJbJHhE6cerCdKg11ELHLz4zzRGxDpvA/fHYYawqSU3rHsipjjCq+Dv7Vi+nv
uu00D4Sm5cRKO/4n4xULlJtAIm4/8GGz+/IaUY0krnAMe5vCF5qX7AifdlahtSYuNUMZjQgpGQPv
Ur/pSZKYtppbcp8EYzyvYItLmuP+CcvIsYVbBl6pS/dQv6uoDmuQDfnFUUxGEhsrAuwJesx1xpRb
6uSF10a/2Ep/qgR2rkrPiImELAZ5O53lc0DtPDWJcEaQa0pPjHE0pUbkzlTJ0SwES7B6cdklQ/6e
lSDqzZIsdRDGB+7C1mOVQr+Px/0PYC6tARKMdKuwcydbuWuduqFgiC8QpDdxeCFnmVCvVy3qUEJr
Unf2ATHBJiQ+6VbM9Y55TwrOTcoIoEODQsL/9M7Pko/AjZo0ZntWrx+hN0hqDeuU1RsCqV/5mUxi
zXIDcdz+tmqAr16z5r/KrLOJ6f3LCftnSQoFrqcnieN48PY32B56ySueJP9LucR7ZoV0P6oeD+Ve
VdOkluQgOJQO+QVta6YmrZX2xvmfrefPI3epRE5SVvIWfvTxtL/nLB5CRBbVGdknPEskOZYFfVXA
n6IVTi2UvQXnAxyT22ze9gGMeA0MX/tYdvdpPC3/zqLMPWz1v85z0JHRiJtO83TSCH3dzYG8q+4z
lAjuGzPOlozV81PjzYQFtlRGQ2Sh1a7Ladz0f0X9n5iGI0/SZyU7mI0SNNvYDQhKEmMA0aKlJnsG
O1mcBKchNHZbvLgT3gvT8aruFcUK0KkVs0VIzM1XRqlSsMj0xCmMXBXA7VCDPXG4DzTGHoTBrndv
X1FGImF1wy7qKPRsvnQq1xz06EpI6UhQeAzuy2AZMdhDNuzWk8JXnqlSI9sJ1TOTmYgCcEN1zjd3
c7DJ1/GgyA10nVq+yxVsWI1J2zyrXMDcefSdIYp1Bve0zw7ByAWYOq+jqyXodJEbg2gLDglDP7oH
He7uM3KUDx0JCDmRchlpCwjvT4EFrk/Hjwo8vyq/e6L8Fa1z0wVQ/SiAj4WcKGyKiAQdrnOclVin
4kz7+ZcMiwX+jpCXcyYGJMRiNEmUan+gCV0CPeykt8lWCcVRAJuu7qChh35VrLMPebuiemkpEYAZ
PiUBqitXX9wmasX9qBxHiv0mOhm0uo8Nwchj/rbsir9QUYOB+yxj1VfodpHnPhVO876Ff54sHbs6
BnR8f5PnGcYDoxVOfzFdimT17RSCWb0C+VIEfwWIhEVRLGJrsffQtr1+rV2sfHIBpRbMf66XY6JY
2ch/mcQpJxMjxWX7xrIho7wIwF2Qs1fZla8UrcqpDhtcxL6rnRqhCif1KEZrbQFVsLN0FaF1JM9s
G0qjGKkgLcBrrjL2yEBM6bRTmNWhQX061kgiZvdECx+8UGPU7huTrMDjQQDX2lUGeQKmLL0o9qP2
wPebfw6JHz5Y8CGkkq3kVdi2hb7tZJcO97uB1sKRwEzU6LS1V0BcMBv+rs/T80pmaeGsjiQLEJNH
rMRXk1cugdxCSRnxYJjFIPDZR4qMQ3OtAy8aAocRx3XrOQQ7ICjj3vKqubRTN/S+PMSF1FIjQ2v9
nGo52XVeHKYp+H2lnIfjTfREZAOmD4hWiU1A2p/GyNxG0zMqi/1LQSeKFU1Oq8jDHtAp6QQxapYR
sePtrzdh5taaupYxP3JpmXZ2NtgW8j24o8N0gzdKelS+EpQG/hmrLJht83b9rfgQLAXZEvfK4c+E
sBcxfy1YpBqZOEgTHooeSipwUaeHUqsxbgqpJoM7DXPxbcG/cHNva1nkACNPG66NjTb0ggWLmVou
M0SGjPM3jAAwhnY0s8B2ILW71G+1CG6chn3Aa2jHUQ3T2Jqp1gWA74a9BnpFf0Lr3xKc5u7UpUIV
LLcbQBq5PE0z+nApEpsA2zoSJd30XUHYGi/KZ0r6c/fyYoBZ5yQ3aGdvT3XrU5f+lSpH5FPns5//
PFxX/PPPNUxXkbDK/95NkFhSFrNIauS4DRadw1TGy55xX26pNBApzi1FPEsWFHCpxxfWS3qEwN+a
rKsroLVYfTT9NF4d37WlGf7N9vUXSe+GA9t1lbW2IXAi6XBZ9Y8WVvSOuJ1cMkCYqoOmIZtYAPSE
6y1X0quA31ZmKtr/HlQBoUFhmwAsyQJ/6cU1PS5CYcjGyjppG4bkKUT+h4Rfigh577QpFxTyNCpU
cnr90/yZsm6mlA5Pr6zVrUljlOPewY09ciOKWpXm767yDVzeHbQESkPjTeX0HGb7KmMNWfSsVOWw
a+pwupg25Vnpx5z6zDl685J7qNTa0s2h1DaXsgFg84l9Bkmdr3gMmromfZUQ9XaZoLw9EvErANRL
Ypt1PfhJgTNOYA4/rpM2+qNVuvMXP3trk61Y+ehNZOUJtzrvi2l0hdR4aJAXngQ2xOzHM/VVJfhZ
x5FEHV9ibKXoN/YqjFBljpbgli388UnZho4nBkCd8oIAkcb5txjJm2AJbq2EuOaJ0ZDzSmqlDN86
28Cyjr2ayjWqw2310o/3JkeJcnR1PDZwpvbeNdb0QLOXw/N2qiTh74mCobm7zAocuAwJtenftiBP
tcKdB+sXV0kEOaJrDxR60r7MthvIoC/mag1BsQF4/A/dtFNqTw7+sb3PtihMP2HS82mQemOoKTps
ZsbOme4qjkiPrefBWs1G+7VsOWA+WweZQldKWfmSnvnAdwXezRhx+9B6ksSVH8oD7MESGpZeY7/S
YQs2shd9QzyxjIuV1Ab1kdSzP1d3j9/r0k0bHsFdhszba3fbj422paWIDbOsgTm75jCRIP7QwbiR
tnTJMviF/qKyJSo6CQqPsAqeMTwPDI5cRWcnrYG7HyVZ/RC9mrBPRVd9hpSA2W1oG3jNDElSSnXC
ozQxWEAzAs0DOzcaQPe9hExbkmgwiH2W01S+Xo0N+szZKnEk973ol/Ygvf1LQ81QmtfMejfbVXWq
8MWFWNzKzCrLGC1AWoElLPh2NjVntQkuIMwTpKGL54rqLMokFGxMk0UCBRSYOKLBTlMaY/RQV3Bi
lK75UCEAarwjRXcha6Y9jfcZiWkdQy/uqXjKszrrvQ0K+miT5F8k9N6Z+aA68bRbT5/aU3T3M5gP
Se1cpPe71fYY8XvP9Q1FO9Xm+nMDwcCRb/xwXTY/L5F5fxblGMCNLCfpwDzqZFUWnRpasngPB1kA
UzdvRPihSVmjZjn6isFd/LfS+OAINFQ8+1pZMF9qXwoLD82Z14hpdxT0Aq2cAWnCX5+VTMt2EnIT
X11ViXb7gauPOl7Kel5CyCfqdafv9qy9+hdCmAjde1iwT25qUw02OTtAIbxRoW1kPB7/HOpj/Jaf
gE5p5AR6R4X062iJgk1T9WIqpsj7gJR07mj2d1IY9JXAvdhnpA9dfpSreet6FGBGw8/vBjJTE22i
JBf0su9i1SRgesLF9bTAfN7bxQivGZFBWeN1YqQZbu9JFubBs+6rzDbMqnPWUu8WoCIP9AeTFuIU
tJdIys7ldU7EtWW5HNMnXAUJQ5lMYI0Q741QrF/TeJiWV5tytKSrhfmQzgwu2j4krtxeuui70XJW
oiiOG58oC0zY88XQEUyTmYTvhKiG1JBMtREHD/jEArMlug10716uwglRT/QyMAysGEUTz0Q/bZLx
1bp48Bx6D9IWjgJXdFqutnX7ijKmEj55bM02vm3ZECqlbpUzYaBN2PVZo22SFoJ/dGJyPvXFf+N1
NVGs8His83kow/4J/v2QIpmnflXFDAPRm1XtadMPCvUQYKpvJ87eQIPZwwkqssem4d6AvQSfBnpQ
qofQaviVlNNm9+60OPtOvAGi8Ql9xR+8rceYekEQFUuCb3qZ7lpux47JFBsWCqtLoC/hl5pDEsVY
WgLG46mhuoNn7d2sf+gIHKsgCN98VEJNgnnKalZZ2jclbCrRPnaDW5Xp+ikSc/YHlBgyLYODVOA2
F+s/6NEmohz2din0y68U/j5AcQjt7U0UQ0DTpqnDs8GTT9r8rxmzTqNdRgq5N0XUaZKno4mdAneg
8aYBZ18RRQScHllBYvVbpAojJnZHsDY+8Un3DIXx3Q77FyaGcmdjH6YTW/1dYMj8o+eUuwPK2CbO
1k92Y0xE/arq8E1+GMnEKe82vIEv5mA0/eE6AqqXESHi2IOvNt7cTmK01VoDGX80V8TFklgLRfZ0
GWYZg+TyQXKE7m8w6+XQeP3cKtKqSh73qXXXvUSkFEv2P03LAUnQobdx0CT9/BMflblPkpioyHtX
D2L/ex9wpuKnp7aSxJ1TtO4XaSbUaPSR2RKYXbWbJBbs34ag7cXgEgzgejhgl6q+MG4tOIzodxeg
Hi4Ebmh35dDL1hIhOYpxstKdRrxb2UZm8kNB+9bXmzsYwOj08BkkAn/f0QT+yhb2mEKloDtXVH76
GtOhzWw0yRYHMqLEaA+AfNLk03TK9G+MEeN7JKES9LDL+m6bCOEEh1ZMp3qioxRG2AjTqY2wYYb5
o5vZgUJp5rVagKUPBEYGAIJN7vNuhkUkQg2PUK95Xc4E9cp1M5tcCI2P2qBtDTQIBhbSgW75dfRg
ENVitlpJzBP8qUuThyFBmcG5P87v+jhjA26/4aVtYzo5Oh6x8FGt7ZPBIQpwPaOUlauCeFeNk3g/
QLtUlV6kKVyd65fdaiV2niGD2IEXXNIClcg3wk1G4KpVwEhkmNJ7bjyednWNJKpk5lFGDNd6918d
n4bUmfCdPKpiG+YoqB2SOx0Ryre5dTSwWGvvDXpBdTxTqpGYFQDdCx/FdImpz+h5Zo/SWwFmr75B
sCE6Do0DWg6oqefsiNzv09H0y0aZcf6IJ1sCNAjf2w/9r3uhLRU+Vkw6pbw3BGD7fMM4EY0Tmdsb
0a4x0gMt+aDNePKCiQmV21t7yUiTV5ESwxskNn4aRTu7GLQzzOAAonYzhn8QLHdca0+/Yem3J7wQ
v6J6iJt3Qi2fGO6fWCvKPgvIJGwxLHbYx7p1o4atuGmsCMZEncv1WVE9mSQekfST11Qt0gSV9msw
NTQGR6WWcFEBJQMUT8yd5gX90R7JXWv4+W9T9Kr902iL9866mLLPNA3T0sZTwWMmXrTgN1CGWFNZ
91Ej9pl9wEdCq9EQdUPkdc+jsf8d0z0lqG9lnYt7FyjaBtmSeesySgqkDGuFBusAT5+Z41WaJdnu
lPECesG2l2N4+PvP1XCwOhzBn7qII0b+wwTLJLLY++B0XTl445OHB6vFGpkAaWzM+VDCw31sQk8U
eZ0uhxrc+98Q1o/2U0a//cIMdkwV/47tncTh5MKliUr4Mn7Nu55fSVILYGJ8PzYidL8BpOt7bBJZ
+om+T10z+RC0bmsz2G1+h+lbCZprSgpldcdgnP8lJUCrWMq6lj7hmWNC8X4bFgdOcR+GPfkT++lO
PUmP4RXiL3sUqXN/80ac2tYpQ+NQvKi/GhjsrbGssuL7LfKcibYYa+zNU7+tDgxau00ADmTNo0Xm
hQ5urXPW9nGNKFziwraiwMFQSenuOOtQi1nXzrG5y0dkyVT7JCPEhxZakR4+622/z/TouUGtByQ4
khEVktd8EGE52t5zkFjd1WHtuYk3LL7W9JDDGx+PfyyTScBNyrQfnF3bsWGEzGBjhjruPFrZPuog
a8b6W0XmPDKJQlRc741qSBw/dn6liQ/cYDmpgVTgiN9s8nq+rMYaOaOpvj7kI6CBb8AHYU0syRar
N0MrRt55r9ZAQQKB7D729lrDInPAxAjRWgZt4CXGtksREPdKctENEM6n9jJT8JSVIrK9/U1t6idl
jc2D3WWcnxIs8EmEmEKLn00Hz3PBFxewGkDeZ2EutNMC9lt61742owp3hIftxPhoM9u7W9qbZ9YL
6WkbLA7TGyb5xMBgklyyVh5OIu/U32sD6Rck6E1q0NCdmCufEX2XQYc6wqcBi96Py6YLae5RahU4
e3i2Z8CtA2fKa82KlXNHVFKfUf83gBTcGv7kwerS4JkfLOkOUNZ0jXft47a+LNaEfzvTBITDHOr8
pRjYjhGqdJOgwu/plwZw7zz9LjHhX4p3t/Lji/K26WaWNJm7iinCJXHH7gDn6gcOeueS6KgBJrGr
36mWj1j2perxfkWbv/MMam+SICFny+vYgaDodGdQrAVjCoISuGJ1BwafV7PzSCe3KPObtm6MoLOL
x4TXIYznTS4Fb03X1ehNJAQjKsOqEwHg337MyMvFWefgFBC1Ipdo8BWttJq6b3IyYCT7GhOtM5Yc
i65bOFW2OCefptQWM4pSRlUujdxoCsSGk3DAaWJfMvVhLUyyZ3JUon/w5433wkQ+fLg/Q+K4yKW5
SKsmM6z/f+mxcIp9LVdwIsVAzelg/0j9ktUjcjuCoCmSBEYmaMqkv/0aOFnnzCEKlyJBghBLY5Z8
vAU0fGHrnkm0EhSboIfT5iv2Sbl8Dbw0aC+VWM/1fepPbmC5ExhrwpsdQBig27VWtxsAz2cf4sID
m45jNYPEQ379+nR3+xfbmGKoSWJtPdsLgsUZkFbcIoDMmf5SOx91tMvdVvsOT8K9/b1rGp7yke+8
8Bsl5j+mfINX5NJvggILW8wfQw62xHvHP19/IzcnOHhhuZnhdKtKDoV7A9tbJNd8SKmLKhmGQSlV
If/lMs+OyZo3CRnSqaHmWG1LtL1wifsED4OhsWDohom1FdR8GiJmC/5AGEjC6wHwj+uuc6h0WdFJ
9AQW2JyUKuTwqreJ4n19IKwuKJDZOc03OnesT8ReX+S5F/+JtoTcVi9xErVvvhEtLCpqh0SAkHYq
MS4WJOf8+cE2AbpxPXttCSeDtMczz/iJSr2UuIeDgjALGDivcGCAVZem4DLjOEoSe7qmqlBY34rC
m6D8LOYaqzzG+rv8LDmrKBggJpPYXZQvrehHVAIMOHMocvsBefG8xnF0iXlWUSMLsPyjq10sjprG
r+7jrwneC+R8Pk5FKa6Tzp6CcD602LhcBiJi+QNNofLRVFdNb04eCfOv/Bdmn/hHjPUaODgs6IZZ
ApQZpPoPrcgWIC/nXXXGexL5qYEmA94GqDowpCf+eGdWCP75S3Ns0lq8teysV4F/hXij0rEh532h
n03YLSfm8LAbjqMSDAFukg1wzN6wYsr6gdga3GmHtDdpPfWlE/hpl9nqKn5jlG1PghYR9UPpY9y8
zXNVIp60VuPmMFfTVqlfVjcUfB2DLe9nUC8PFqCZOVB1HDnS7TLwfNvCm25kwDes51zSz5K5qvTP
2GPoLmAF/sWi8JcuEHFaCbcWBDla89RiHcQMvvYuv7KImcxh7cjFbbQBXMtEkDZGON4vVHJ/OYdC
AdJnynwE9Mq+AvbfT+Bh1G8wAb72tz3iTqv/honZvg95UqZ+bkE6F+z0V/i9jO+KlW26HB95RLc0
2wGrx3O5f+02mab4fNtBvvEEwqOhVjRTMTvvsx97EJCFKe73FNEYlKXGIU+87xSyrp/pFo3EZGmD
xfz4+IUhWuVNH9QWe6Sm2a8g3KdvgVFRFWNpO98tLguEKSe/hTztkFI4WGK3GDzclWron70l4yZH
FR5/09CR8u9obSJvGq5KnjgLmP6iy/If4tA/P8km8kax2aJ6kvIHLY4X71LcMRaVvWRB+sNdcDAR
GGHyKeAkbXrout69JDJ5k+7B7iEqnF3YTecHeaasDr2nV6CtPD+O0SzJzU6XMkx5lW0fKXBeUDDX
O2pdHrZczIlgjzC4rLW/3ikMGfUXxB/f20/Q3BIRHuw7PqKSQwnOQ3dKkiqZ9TJe3tbCiq6lspm9
J1BEODJtg75Yigy/ozqcBXu0eAowwAORzkSJA/TnQc3zyA6lsTeyZoayuY5mZr21RVY8FmQkk4CG
EQmP16oQBy5QUydP91QeG4NbakiUqwA3uNx779OPZzulRFmnmv6BvfGkXzXqT7QsZMMRnqao/NeJ
uPeQIq12ieWvajMYKoD1Mib83GLYu8u6xTGPbOTCXFKwANUdFIXNdsaplVpF6W7zayKNcTLRY6wE
PYp2ck04BvEkzIqvTO1QZ1xgOzOCssTWrwyNfE0PeW5oxHxE7tU/vkawuAqcAZ42yGhCHq5MPlI7
a7+BaUJuaKMFnNxMEmQHJlowrB8tEWcDErF2CwdM59bilir+SD6um6+sLxCj3JUt74YJxnQ2O3rY
Y7Wdv8p6pl8lWdJRTuswcKw1Un4tHHIJWSMC5Oi9ecmHz9Gy1UR4kXVP0kqmD4bUieK2M3o+gEEN
q/KhE6/E/WnzS56rcBLphM1/7CtGB/+1qGpHMzopzRwtfrApQpC2uLiLcUbWO+OTQ3A8j1wg/hnu
eGUeTYahkNlUlrk7IYde18qkU8zI4mtb0rmxZhyiu0JjnJXCSQCPyW8WdU7C2qxghpXb1xhNu7Cv
+ZsX2CPnyBhH+1CoZpoJcFkGZewMnfZbtB0TxqO5QTxIfbLDquUrEK3cz8gPVpywJ/5InOfgfNdM
f2E9TzbIg49Sv8g+Ny6AnyJ7ngJkg8uH4bRyiW3vDc61fQTfGkjj/xFv7Jh+juqjncMq1g4VePYZ
pkxgbiRNSE/5AfW0+vRROaMM3u0fYTARniFMb3mG5+Jc/yd4NXSQWhhKpBfRoYdbRMzKXLcpy7ie
5ChxC5zCO70iFN51aQ7daB4cWapgX5Jm46Ifr3bGXv6nTLh5rPu0xryKYxDCDIblLlGDrzmdyjpu
on0MyRPuVjbYk8BU+nW1E/bBp/jZxl+G3R8Fe29yA+Vv3lWnuSCSVfEQyZi8cYXxElRNUK8hJxDd
SuUQc8srRO4HcCZfsaiAl44XV9x4lYDDM3ZiVv3d/zsGlkStx9epBNewLGzVWXAi/ucsD4DPb6VV
XVsF53u4s2Ma9TnUqNSJ9NSnarqyFqI3nJJRhg+bQVvn7MQS1K2bYOOV190eXUpITNLKUhILDcpo
0UyYPGl2RZl77kBX6IGXSESYsqwRBlnmyHp481cyLDljXkGaZ+GEK+nOJ/sgmv5I5sQGor6STWC7
3RuQ4sjNlhQbMuovowyhvR5s/sS6CJbWoJkB5y4xqyWQy5FxZ1GqR0tGco0zMkru6sBKzjv4uYfS
D94djQsxquvionc42ZQQm41oZGPBJWCeDiZHWsvXkrNnOgtQ0bfrlv+JNGPYyiwIv0UEPFOpJ71Y
/FKLdrEABzwGU3M22f3QTr2tmqQsNiOGSKp9W2BPBRE2OIf7Rm4fQwbfKV9mJ5YKHJi2Xvn3+wnv
HTIZi5jBijnIAvSq9N2i2pMlg2sYLQMOEWceBRNyuKP8aDxIXsBEo317SmglhvX4rmKG5Q6BPvtH
YR5S1L7N+ySWFSIVSqH2MmHor9XsaRwyKWT7Lcp8PLyLkCP3uh5C/7FnNSNgB8z3QcwXn/p13JzL
Mkj6i8TvcKzZuhQiwvXxDK1lNVBB6VyZ4bZ0FJ9IZ+1NE5XRZTdhKZtgj1AKecSVJA7b7gy6AiZ/
NBidWZYozQqfPOKe1rpqZoaGUKTIfNdslljDvwHeAyhpBo8vxBpY+NnKWx4RPUMROQBbn4c9jp83
0RAF0tv5G/hwtPIbUmeunt+SoJhretV7GYKTv4ooCSzpM3KTbKSJZxC7VmDcijUhWPMJthKlpm+X
YyNpdnjmNUaq6XI6rTfyutr+yzrhNPsAS50Xz54cVIaJhR6bQIE99O7Hb+25xqRjIzvNTgHWW+7P
wWOoxI9wEPQ1pDC7A7R8fn7H+SJeqsCqpWvp+VEPII30P0aIUuQbdqznG2aNWnWqJJWi42vygZg9
bPdYnBkIu2rPtpEwSLE+v7pNwBVGkL4qwGxOV+LGfo3dU18dIJQb9QDzGS4vKBvbY8aAIQY2ZLz/
jyvZfjz9/9bS1QI+6s89Rqx8V7gk7gm9Q7tjIYiDfO45l1XxV4PFKu2Bd096IRdz8P/dVA8OaNLY
qxLBCS9tMpJUbdwNc4HixBVdw/kbVb8yf1aPaDoSCUWHpC5epUKYtko4WC55xuF4zoGC2/xczaju
n2NSSpSfqPVmD2Y+Z/QyD8/qtiX2a8US/DNpqDyLGoq++ksSrJjlhGcR0yxl1QCi7PZd4i17T1sx
WXV5f5TE9UQRHDv51MDWzx4oCABUGSNHh3aFwKIOuldZSgIpvr0Varc6LhOH5o6kgbpxyAKzM71Y
diGdRwRAAQSTDSupERyYbZOmP3QlAWQeHL6QZqkkjP2r5l8JSgJ3W3lmJMHxknTC4jWinIVZsmR6
5oWTIWKUlNTc511TpFQKxgwW0NyJmreFFPQOH67W6ux38fiRTieiAaqiiCgUvbB/bvJ/RQdnXMen
TFX/GJpExNtGcZwQzyoLNQd6d0tMituCsIyD0nXRQaCJSi4aBz8QctlvicArCcN9a8Twlb6+Zi2G
cEQTZURKAv0/w1+onpcNXNIxpAoGsUPyGSEmusr98cx7Kt8tsiuD8sFHJ1HigBshOLcZ+zL/MVA3
RgrgTGUrBeJi214mW+zS2pO4T8MMIZLJVktyqbPX3mrZU/U7NyD10LncEXrr292YHGrYe0ZBVb1V
lXv8bUIbmw4bD8O40CvvESoYDpFI1yaosj6uqmZ0RwDolpF+WkYra+bsBuC1ny6D/X6iYX+RIsoX
mkekI5EE1aP+TLGmUGhTgJPmGSaFeT9pZis+k436eRwx/tg+FOkdPcv4QSPNGZkfBbaiOkPm9r0I
8jdNJW0oTGP/d5exTPPuE78X5rQGWJidO1DcHgH0bIkCgzbCzCElgFhhQDLxynnVm0eQ1ExDiaPF
xDM5/W4/dhNrlqHJ6Vf/0s2Wh+cEkJDqGyRvVGZQRVowz7fCziAgjGlTYSIOqn8jQHBHCg6RhhvA
n/Wx7WTkxKisfzXDq6hnnPn2ToREvX60/Ku2PZ3wqpk2xM5T+LCIVndzKz2oU67sUd6vWW25HV9K
9Tit7kLkseAq/epF21R+2V9j+jmVgbIzYRMEbw3NqX9sm/zZNxg13zRyW37bm2lALBje4UiOMDPG
RI6f57StEKx+Jf1DMQmLoBEMYCTeWcDK+qq4WvE/m1ONXDWtFAIcnvrQOhGyTxADCe69XbE0wPmz
dmtK6lSO6y+dhlI7C8pZNYFDZYXMtpcEImFdB9azli2xWE0WVVSyzS8g5JMwuhsQgsy+wVSk6jy9
6rN2URTiiTVmM5rTgQWMw5FaJItnB1atr2pOCZb4VYpAy0Bft2qMyXFDvlU/feNuTx/xsTG5cWVX
wmV8bSZf7d1Oh870LBcQjhKiHPAesGyWJLZeOqmFzuF9bSPilF4yB8Yqjn9aUnorVZS2GxsdKzCO
saI5fivl650WuFoUhF7DI/vaWZuNavQh6W0J//0EvlBfWtW4DLtJM4Cq1Hv9uFaQkn6dbWmsgMZT
UkYfvmLn7ZygfEibChB021wbd1QuoO7GEr23rm5zJYl+Y1SPql3svCXErvRXeWHqqKUdCIPEtVHi
FJmbDN8vaLxa1rdbm0w595+Uf9UYuewmxk2wcpBVme5tgMHXQ4W8YzU5u8KCQrNlbMXSTaDoBZzd
xf6dMChtp9PNTugI8JDRhvo5vZR1TnmlpZOfgxGG7eq2BwHabQoKbHt6IMFrQIibGt3a9QjLghDN
/MPHHFM8WouQM4+MMegxg1CTPgRm+ivQpsLQ1CNZMPESDFaG45/ZzJBOf3s5nBIZxXfP5nhwYN4g
zbxHRFmDoI+fKbPd4d6GSgRKd/kDtgdi1P+qo7Y10riyPqyAN59w3Ybi28hfUPVya332bfDFFWFh
kZ1uC84bjhJ8v1k2js6balmZKJKkiPn2r/FUi4eqxDO686WvM9pKCcFuYX6PK/TX5zs8YkPOrgGM
PxSpUDBgLhwt/sarhR5+BtylpCaNaZyrCdYiuOjz8c6B+gLTXsWOe2/mvot6WGzSKFr9lqo+JQTf
Sn1jYlg2yIlOmpU+IMyLLcuzx/CuSModSyqg9/Gq/kOA3T5+4jVhAjRrNk4M5jTBtgrDOO1b+PuY
wT2SI+1icXNWQ9oItKOnNIQ5/5wDE+P8t2jZRDmygRSuCkdAfObqhJNLpVz1U0oafYqnXNfQkemH
9ChCPk3e4DPrrqNgAwh/nbl6MfHeGfF2VM5ny0y9djQmsdKGCYD2Tr1zbqh1C2ElWyjBbsCIyXyQ
C6z7oNA64eIYfx0YJ6nv14Oe8ONwxnJT7/LulKdKEMAV507CRASCCNJlnUUkdzBRUoXg8TIe2zB0
AODqaIU6zB3prM+4G354E8QeLtsLHh+ro3oY9jzGw42VwHqrsEa3mT5jHjsj+I3CMjJFGVTj+CXn
33e0jq90C4e8XkvXH3q3ImQdo4udBjcy7tbNked2Rs73H1IOaKtBgWAlR4S0YaGcTwXPoVFCbk6Z
hIYNGQN2RcPy7FoF+bAFV8FcsbQJWVhFJdaGdCDPkuQo8hMy0qond9rkv6TTXTn1c/Y3iRZzYb4I
kCGsZZrkMJ+XT0GY8BJyM3L/Inx0VAqNqfYlTupOTPStF4nDBW600MtaZKrh1WHfaWep/i0DT5sp
+0VMLzW1NnkKtPjGGPsYybI6kxyLFOsjpQ+RPF2QB6Wz4ubRs9FyFOjGqOtZv6Bd6r6nlwL9esE6
8BS9QIjv2wMe60VwM54Cz9st4RGgTjsoCwiqJHi5LjUUzHSdOTxS7cxVKhSixRu4OgnjqK3MyTSZ
FqKW2etykaoqcEPxU6tq9Y0DDEGsOO0rBgVLJ7/j+b2fTN+YETRCBkY51M4dtevvT2muE5mTS13F
n8uYCZffGCCvX4d5yzEOtm5UpFVmhxg5ltZavMRLyQ6c+s9lfbmma+J2ViWeTofNZKK1gBwrWGx6
xZPn+R85WB0ukyvblJ7YKnbjqW3gSs/w90wrPhZOTPMbTVuIDA7Lev+tphvY/wWcUxDQIBCCekAm
KcMPoChNrebj8Awttb8CHFoAGf8K1EbfUxxpvxSjk01hcXiFidWLeWZ5VvoRG+ylashcuMYUMSJJ
w7w9Wr7lsDifDk7p6Pgo+O8aR2jJtCx+Az4FS070Xm48URtqBZGoz3ZtUi/rv2pBouJbLOV/svMD
+mD5D4xoEmrfFyIQ+ljjawYoiTjhfJ/pNoGr4Wi3PlJmA8TU9qaj/IEUUhqebvM8DatrT9x5rQEa
lmXCNWpFyyOYd6cYd1JjklAATvPC1A7a2eWZk0skkByPFQBppqYMiM7fa2Yv3M5MVwg1A8r4V8Tu
11MycAgyg9oyx7tD4714rKkwyX3rinaE+4SbsGOIDQcBAH3IOlhRNcM5C0fvMTCFU3HCFttJW9TC
IqT4Z65RTgVk94VtMYTXu3xUKvgZzQPDGc1TBmLHN+789sQtHfVyndandRZRJ+YwWOV2bQ318Uam
+eTnrN7LNZo/ynAPJHo9axOM5ZFgaASWvL3WYgMZhLsy3kZu9HZR2ozcKynrwaFGuTiBAX6r+w8I
P48Uod2ryvOWe+OTsxfTyyaTOvKBZSAxoa0VsTJC1ZGYa6Ry/RlYFvDPKtRsTdVou/gTik+lJh9D
SQisoFyF2gVANzIel4EucsA1IBTrFHOpqwOn4esOmSFSaUyN/VFz7PgQZXIk4ck+lJxLfuMUBnFF
luxq65zffWF+dOGDi+EdXjHzjDQmljgtUaxeyUmkrPaVIrt7NHy+J43JQNFedyBignx682OQL59V
OOShjCmDNBVHw0uuQnrDmfgj1XQzAyoJKAKgq5AIPxhnwBSbT6DahuGD6lglhy0tYLIm939WQ9ad
6OXQgpV2PTN3aEtyb86+MFgYhTtbO7UvGKgIoOzuPbxG1cB6VrMccidlOkdXebxcWIkg4iYCP2ef
631cNt3rMEezw1CkzZx4/6iZXR35djg962uZxseew62A6BYdiX8Lb9LWRJfCpE/gHriXu9HB3NYl
L0k3A5/L3Y/yXPGw3IgsGDwjo6A90fQCaHDOZxRYnQGtIs1LISuNFO3iX6S84TpgrdcprqNACj8+
hu08CPirGhqfuc7TOCRVeWx/p2ZJ0BS5Rg8LDUUTunas3aFFczqwfeu5Cyguu4m6F/ftN6WTAmff
9J/XynkeqsXGxpljybEL1U8DY3+TyVnr1abODx1Osz1zpy1o5yoOueCGhr6bDKhWhSDuQoYPW5w9
Jq1l1SMLGsnOxD4syXnxenwJrHSq4i8+AmfhsLjeu+3xlufZwB8TozKj+wR9gVcZV1lG8cvkoBGQ
2rAnYzoEZtXuM+Vgn+SWQsvMEloqFO2loTcPFo2KNoth0PwK0k6iV0H+EBlEUm9VKffhAnvfgB1u
X2ofm9Biegxm90T7OZtm+DFDu876VuomZF0waP9aWDQq060+X+4GDHybFekH8ESnMGAsVKzhNx97
TeaGqcJjX3qMsx5lIcYspsDbiCrmBoMTKQQ7vbWKtnWqITug2C2TuJcqxsCQqgJlamAv1g1SGmO5
5Nm74up/Xww2LhUOn6KmsJad7r/qJWdJgbGnmnaLpBNv8QlXSxlBv+ltOgzwTe+w6jvotyoKNnQK
EyGNY8j/cB14KIRvvhw9022yLTPAcqirmRXDO7o+iWNdPqaTz94JqM3A2LS+rmBaC3od92s0MvyI
mvf9fYIogmkXMT9bDWOVCdk5sjDlzehHK2zQu2zVvGc5xAAzXv81Ofi17F4w4Qdi2i8T9IY0FHCx
/DEZ98ogKlP09Ehe/YyIj9n7oytVfDmrcgrVe2v6085ckAck7RlFysXch70BbHodQCeXfDyFioU/
9KLftsvW0HTBsIztgqv+Sww6frvE+pf7SkzHxEFBeEhjpAvmYCbQLP0IJ13yVD19C+nZHtnXB2ZX
5NnRUIhROzH6QlozQqKrijhoVHk6DOaBdohYzi0xtbHVYrMxFSTiqTrNYpAADPLq1nKyQJO10GYy
W8koqQagZPnADda1GNYeclnzjw6B4JCk0DRQ1i8UiMX7X0R95SlF5V6AIOL9uYy5rBeyNCIPbAAq
Cvke7tXskYoW5Pyeneuhiu1P5LXXd48kqxWq0CAmreMJilFgr2IucrX6E03tDzxXrQrHxfjLCSTr
0nqZTfzXRT73eWhF608YjjPNrCkSqjPtItOYDpm36dYKJYpuKrcE/K1IY4ezjTsHNYCSGGmevlGh
zoSvEqWPyHQKfrKQKxNJmyt3iwb8thsRUGGHHkQqtj4Wd2urnW8VRtapmpPmBQYRUzKDLt360B8j
Pg9FT+EcWXyi0GfogPH66u0dWHJB9iryqQglFVxspmBUuj4UHhIYbQUT9imiUvzMSwHoT0pkTljX
M7VjnQ7zmdjxFUfggz1h3PBN+1xldekmBEf8oBO9r8lkq+UyyLrLOcFsk36RV0Rc/ykhPjHB8ko7
Fncij9TK/Q1bCClEhQ0u6UBECkNyml+iMXx5H1jjOY+R2jU4LW84l3cqfzqlPatkx9CTaDQSz1u2
wAQzMsUqo8lmWYj4/4f4XNl99OPDVmD9k5W6i3KcmkZ9Bk+eygWdC2w4WjEnajohXjKQjiRgpQBg
e4boXXt/I+10OUL9i8LiO+cnK+gxeOG1ce7KrZpi4XIldtDadIUvhxkIBd4ELhPTdjcycSyhU3v4
L85vdJwUf+BQJZIchAh24bPqQhwfWrrUb3plGISl19ZJSsUlTadedbu5zzCzGNj0LCsrpCC5diBW
bbLAjHkoJHL4KjK/AB21cL3DYAaKI159ptmg7JIHeDvyBJ/KbdYa3xHc9XeZUlMkq6XFjbZvwBgP
0/9pNSsrzAXadE9uuqfQuyYOnZBTDV+3O2as0UV/HLeyJecOE6V0Lm+2NY0hMSPiLvpCjVO1uCl5
5cJcrGoDiCd5xrbPa44Qk48z5HAp9HYXfTsY0V9v8xnMpOdCvIQ21DtPD0W92gLVBtZRCSKLzYOq
IQDe27s2CDp/JXNMbR14w1R+41GWwcX94nb6J5R3kcvi+3TkGj4KpQWixskRgThYhc4hwaKZsqHW
b+yDmY6jQPNNDrhnPgVXelrMQSN5gSN67kLw9NF5arXabHzqzWi3IxdITpAQvWcyAsKWMP5xBno8
j/39JwTPFGK3tCo6Hn4FeXnNJ2RfDuvqPiLTWnfdEMvDiggihCCL25nqboSgl8kncaJoIW8tnRkj
RfBvGLVXO388yXWw+S/aK74xwof/01qJLMcFgWGu0q+tIOPwexS1XBRJr7571uNC0sC0YG3IhiBy
GZTufH9BOBrIpTg7Ik8G5wDUkvlmjRDvlTv5asmnFLgGdxtjLpONFqVjUwD7mnS6YdxSSRDCgzgs
AVxTmO/3R039mhnv1Atw1XIKsB1gn7pbvdn0bhViBCvS897Mqik07WVQshB08HDKJGfxGUxZWXRH
XLDC59m4FnzJmIqGKNO9hdyTNsQsE8IWS7H2NkhLXleqdEEoUHe55edL2BsE9EE24RfMvYVPt3H6
ZuaelG8TQseq6FVcGzQvMIxd+PaEufrjry7FboWRL/0FBO0BPXx9c5wJiz5F0HjlX9wxAsQ4v5eV
xG3YBQJhYtjkFASJRGKS+uIB4c01x6Bwvfw7xbtFRt8qfuTwb8bkhDwPUXeQntUFOJVOHSaiYkuv
NuRuE0wqbdnqUsWkHgRfWSUmCPK1NiuVfA724C4Lc2Em+LOP3Y4/FlWbiVFHc13f+VvzKJHvDINx
Aa638GW+JmPr01iXkKSy270JAtc6iiUy0g1Cb+t217FhiNYZy8ylJ8KB4isiNlCJ684+MQamqGBN
cIomVHTVEifl29vzlYH8tfpIeG/zKzOHLi8oi0TGzM02yNSGGtAzk3SrMfI4rV5ozmuapQHBMRFr
hdmYdUmh8vpqV1OZqsa9xH1bpupuBAKJVjQ03wXkOa18HK6ZvOL8qfldQ6yguf1AQ0aNB6N8krNB
tsyA8lQCV7rzcwtdS2MBsseyGx4mqgAxXAoC83nO8pISz3fO3W36+NJjnbYTQOChbpG+S2NoGd47
LDCiEFWHvXAr003f0HT/ZY67vvQv1yBfSz0kBndc7IT3+c0EtPRRJlo9qDQ7H+sKOWhZKVm+Ov14
NWxsnPjzzlDpMQGlUeKH6Vd6GaoDztvrUkgmBGy6d879PrlWQJJq66RUZi43WR0VAw1DvEaWWnxr
x94dfF/cjCGIbpGbYwlRp4TgN8VppE9WNajCku7mhWz4X8hMGho8yKyOoVbkm1bWaNMg8i7saczP
M0QipEwpHWPJa4onBoXa9YUmZF8fOWYwOxpbIAlqFP3K/I3Q+n9hOLmBunQq0Oz/eetsVMV2eM+1
9dtwJveKvg7xwcY0IKsroWtrZvuPfBw5WYyZKQNYZ/bo2hrEfHo5G+8W9R55Gcq6echpjm37Lhov
tZ9RYIiB9wHP1vlV7WBnJjcfq7kGkmxr/zfN6wGjNC56WNXchoKT2K9A5x5xYfe0Io0jeNL7KThO
qPY8iGTQN0WkuAMIyx7Or6YCtbGUriRyqBMlX5MO+IxHA1wVzd7g2br+AId/3XQKyHTWiYM/eB9V
UywkTllgwq2Sdekzy888yspSkL5oooLNvSf0FK3OzkaAme2Ip87s28/RP25DbA5lkGlDhrFnC0t/
0wvWfIHxBlJOXFB9QvIs8IopdD1O+2dr5Ly8dfacu9c7ziyWC6ZH5AlPxqnfFMeFv4ryrsjuR0uP
5FvZPDc3IenlKMdXSEf1u79o48hmJv9wflzjyrvvEDkSKITJzIF9dED5X8F8+qncA9qZQyU717N8
zR4TAwA+cpPh+EVsKY6Uq7exYBih+xIt22Xz9DD0D6TGPAvm4qUPaqyVN3FzT7hVLg+NUkS0wHDZ
n2QZuvf+T3s0rX2mT03ApWxwVskN5G2Dq6Qm/1YttT4uY/Q5NDjiglKv9h0NnRpskXM14rq4YbZc
djnIqJXWFCADLikfZubAs/4anZfJQbxSvyMGQ28tl5Liwol7KgE2sOToxzP3zUZNoF+5Zu4vKZ61
FWti+J2Xqfii+QR5jH+77bqwV5rZ09+EqQ8iydBBvbN5yL4Mk08E6Ssl2G6E2UGdFNkUxx+wnAVN
xi3E7s4dSIDdNJZ6hIJKrDIoA/T+oS8YDGpUYO2wcmAMOulV8VAEz5MpYfFl/Hp2cf6Xly0BYXhY
g+y2AQ/hsAFDYcghDSImSK8pJFLcojMg2c5RWvWc5acGrHeFNo+FY4S305gZfopoK0dLI9p/slYc
8/4YFJ8PtvciRvrwzNUqonC5lPEMpJMxvqCjKB3cXyrSj+pniPfWHirdra7UDf6C/PJKBgK04r5t
AQSnaoE/VfLleVmVmicKvquOCbOkDnVGPqB1tvoh8QQIWBEghVcmyFJ9pwg9RjuZyut6AeBaopD7
PAOu0jPZfdgSRT2dPcvBL5GDW+xSr3enm5H/DhN90s5xND/W2+ahG0nI1bK85lyTf1jtRtAlLvdB
sqpu7CsO0xcEY1ZCO6I1U5JBn1F3GbcHVXi8l8duQsoYSQOiLk8Hp5jthcSZYCliab6kFZYUYCau
GYaw8CVlw1aNn41Fp7FiV9poPoNrKTv3P2ILwBeVUeHOgZM3A5AK9URdho2hzfXH/5x2NAiU0rf2
K3JatkIdeC2DQeVBzxNwZBNQKje98J4R4eKwHuQFOpYFRLJrHsEaBEng575OG0jv9NaLMM78KGis
1RCduBicnXqkX8tPSLdVxGYpA/CrqRPG7R7M0PmnvegaXYIO1Mqxr3kFqcNxkVmAH4tZtRB5t0Ys
v+ZAE4SPlJCqqGxZeuJ0lhNtu+K9jMa3+VCrSrqvy+Au4RFAvJDLuU1TrN0xXcNHwrZU0VGlixzJ
QVb2s/IrRw0PkzGtw7uctjiVkkmo7YUhkTQ6HAa/IUQIzyOiKCAXukFAo7/nOgaR/1TFcRy3JhE2
Q97jNqjhovTUbuVYVJCJT3NA6kYrFoiuVBM1zMnxCTPBAZPQOb5X3fejSYD/ExUKRSLAPFnlDXs5
H9kRMTd8bRXi4LfuYpFvAp2T31fvhwqopGPE2txYr7jo0czmUc2/ve6clyDECROlx+hbp9jmoZho
ppuLJk99YTw8D6Tm8s77Xf2TM1jTt1BJZg5fCHIqp1LNq5m5Cgko+JTBMYJvQbl5SjG3was4hkR9
wNkB7t9BOHOSobYemjQUbT0tPefb3hvRTlw3Voo2aCGNxYZuYotWv0MmxQMLL8HeMNbA6IKsTNZJ
AhP/NqcLzH+a4tdhv54McuXk9Yt/TLmGqmWIWvE/uKHDOcD8osvA+6wRd+G2zzfk9nchJd3qzarF
LeZIdhOK8KZ8WqgKfnc4j8JrRVfwiCUR1XP9EGdIv5nyXIUfNjFtBtCbKySsnJu366d04WqS9G1M
2cySDgCDpkQlS0/KRcV4UgL2jX/B59RmzJ0yenDSJnXJGw4Z9WK8oEbRvj5luj/o94jiysIQHusR
9KOVipjlMzldbiWqMVUTYbrR0WPEtX/l+YDKHGJZ4dcXo9sX73HGV/6pclDGgQlQuNXC94oaUc8Y
RI2cZT1gP0noVHIiY1EB4pC4R29tq2tHTOMy8atFmC3Xs/kHM/shCZcMXJghx5qa62Xuxi48eS4Q
Rq3ez220SywAtvJ679IFLHrkcVaJfQ7a34kJtK3w+BIPBinpPChvuOdP3yaAlKW5XBeF4SlaTR7y
RmWP87hjG9Z2P9ENthJo4AEawof0TogeQLuooW6zrYNZj5InDlQPCeeX5G/67Ow/9D3+w2OEZAoc
a+m3ijNGbTtViMES03o60j7Y3nl3cFs4OhD6XXbL4Cl+ItSiEhZAq+9x3mpu04NwfgahtsvSSDNm
NSfFsiLEjm16Y3p1B//vsCmQmjMD0eQRdcFVDWuP2zSM5CBCCuQuIVj9Yu00rftwo5Hmpjo2pAcT
8oxXeVfT5wzjQ8n52uyU9dp54X/ywysVqaFidzjoTzqCb5wvFfuu1+E/P72p0D1hd8JwJYg0090G
WBrFM2Opzb4/RrkJIGzmHSVZ1o5/M10rIekrC/JwqSNNHBWwAdpuICUeqjhvKo6tQAQ9fnuP8l6/
RIkwRGo36kH0LllNP0Twrgrad5Px99PNfG1B0l3+6VgVk91gbIzKmTHR+OsOnVGDkZETMf3AH21b
QRCOMSUnlVkvXy+LeucoNBBYP0TVpDX/yyWywIgYCK1p2SoGJd9AnL2feU2vxGsFkfY6mauntk7e
1vP6T5PMiT3YTDHM82+9RgL4w3lBDgQSfIZkshfyZVV4xuaPffw2PRWCF5Ni6JhChZut4n9OKOxL
6PmzCMmWRqWJ1d3OobAaljrD7c83wuqCU7fAe6vqSGNbMdZOogU/Psb2N441NIDnbC05xnGVmMsX
Rsind/Al01eiA5HYhjW/VKifzEPjuywo5XgiwW6OKZ3CVS2b5QCTMDEfoGwZ1GEMBSHDerWU3UFR
2/dtuIngsulmmi3/S1OJpv0Ed4JTS9zRboZz1ggi5YuSz+fx7FbE21P3dbx44IlzEXJfQnbsu9w4
ZY95pMa8Ale/+D2cMoLUQ9dLPSu4diCo1v121BTz+Um2AC2PPlz7Lde8Y3wm6Uiq9F7W2EJSdlI5
8crVQhlZIIGFSCtRicq3MBbNbgucjPaT/p+b13pvqUR89ycrT8W1o/aCnpNiO9JmNbMp91NDLZP5
zjLVR2bmc6fHHLQvDLyuzEbhN8ZMgNTKhDwn84rJZ50njVoYqDnEMR+b2Z/zTw9NrrJnuHrhoQU5
KKXn/zo5fKo+tUoVWaUorP7yLwltWpPUsZ54S1OHh39lwzseyn9Na0lwmLa4r3WOKOWmaFQTyVlU
9J560Ij1yZjRQ5110wM4bVpDi/tCGdtxKckZw23unROg8xAzE7CaJ2CA4h5m2XJ/pHUzivVL16qZ
6BT4Sf/nxjoNqx2nAUDadJOfDt9sfbXMDPRVgLdx5zr+GUIoNnzJiwiGW7/Exi/U8uOZHHA0MxbQ
wzMOQmgmvx8jY240/RLdFcmZjgfYFRGnJWTxI63fx3OE3fB7lkpC4KQRQ0wS2bHb6grRyW0tYmHa
Fapnk5ZHkgsT5Ey4d1C1hvNUzOlpUGAgXkOnUjWLN5/CO1Vw59T6oeBcYFnXnZhyuyQZPeJUE3+Y
rfB5PRxcx2yqhMa8+yqLSPVEs9xTgzVf5G7lfikSFUOCqU5qBNnx5xsepdyz/vnrwxtGgFsLXz4T
zVZgYV6iyP0ZB/IPmyXTDgleXUyrSsGmxUlA8WJ1KpSfROBWM68Wv8ReGFPF9n0lDvj6Il5OOXTk
lCy4VzxnVTIkrOJ1P7ETVFOxTWojnYXwseTNKtDW/ZSH4iSMaN4zIwmX12Ur1VX4BMzq3qO6ZGIS
AKq131DVtCIdTSftitMbZx92m9ssQFN401UaKZAPGKuCt6DOaMW0UhpHWJGURNTNnjzh4wT+x0ms
0Ha+UUdv0aYHOYq1LkvF21mrB0dMTcXgFNT/FibmkrwC4fw4UOfntnxjYNmYEu2Ep5eKAzzMv1Pl
x8xraK5MVn/dM7MkL1fU1dHe+btPTNQ7Vh4nQpI+pzZNiwbHa5ytG2NUmX1eSbC5zBYvsGUiCpO9
s17GjuyLWdwJlCeyUkMP6IytjXNpK7qiYFmjh8OdxBnzV136+pemqaAwn0OnBVevE0PIR8Iogb0C
CJ+YY3rtQjXh6pnL2W1AV05HjTZgCfTQa0XhgEb5dAuO/1e4A1yZhSNcV1661h3OSiCIgHj6BB1I
F+5myDAR69sIrDPqWPa5AnT2DkU1OZAtVOuYrMPGh9IQvV5bpp5ruuK87oLY8J5VrVJ80XowW3kp
/mVShmsfzMLmHYEUITTmekjOr54NVatVDfcFI8Y4/AQBhnpejs0CASuy/QMNfigmXP7cnZUvEWfw
eq4dIoTAa39gWiePT+VLHz8HW59SYgaFRL7kqe+Fu7Nc0rAEuhG6+IOPbkb7elRizo4ytX0fQSIR
At/9rPsJE0OAsFsKF697RdCBgigta60borGu6aOeGrlKeDD5uqnq5H65B7RTLFvqB0zKM+4/2Ztd
nNQHIM2NzM6DM8j/sw6VOvLgZduLJoKNCBOwN+gZLZ6KW+6G36ZYbDqLOhZviXRUf/4TewkSj+pv
jjC13Shr3eDqsCvC5rbIe3qazQf3ZaA8cQjT1gFG4qMsR7X1ghNZr1F2ujFXLrJq6ze4vj0TbSVx
T/mHL0SFFKY/NtRqpFf8Sq+5Nk9UkcypfkjBGZnOe8CJY88xz2FQE/ZStIxK0IUjGTFio+iYWOkc
LFtrZuqwulghCVI1q3O6KwVPwx5kOqQAdoDSHN6GxYmvRWM1GhH0Bbn0lhVFHqQUrRg3sxpUMvS9
95UowO9ifiy6CCfJIveEZTW2XEsvRw6mMbi3x+SLmfF0kVylQO09g2TkVxsFhDQgT3pQQIG5aRYk
1aC30+kjd80APrGpuL3/dBRimAFmDcQZ4ZofyLZoTmv9w2r+0wQccQGFHMGPsnFDS+eyD6ECgfWb
jt2n71CjY1KdN1vYFET+MVj2GtdRHlZ44Sz2VYOagDEnFTq/IOvAaM3uAJfYZqeSyBVKIPvVoEPM
LgIevQ8rnLqEhz7HcnJqgcEgayljMkyLDd7X3NSfzCTsndL/s+16iqVo5+od65IywoARTz3sNhsd
2ZTXoB3HhMdEx7Y5D5Qz/8P0L/qANrcvPw1ZP+EprifJqQ4mF884TD9ZngnR/4jdttSlpc2vjnEv
ffFmGl9vOty30yqm7c4hoQ86K5ZIB9/dZ2Aea9r8Wo8qbyDBTI2HzQA84CJYmuJSRUS4SdCznS6o
IYF6ZwGEec9KvecIemYoeTPxJalx57o0IKouyK1oVUJgVOdSuUZT5aBNGdQUhQLR7gGO+7rHJJfr
1tmwDly+hxB+heVTGPD1PLw0+6Wzfd+oZbOn7dbTordso4dz1VBi7XIVFlrXJxp9rjADUIlnq+Z+
U0gJozBAw4M66csX10eWbNsF5qn7UAv2/u28fbspSjIOxxtr3u5kGdhlcX5HJSHcTc2F+hzlk2o3
VjYa63B1oii5uDCkawszGsYZhytYy2YiikofvdLpgeFXvCNihWrkrxhmbNtya3OtsyfEmBMecGvv
XnNwyhRZfrI6TS0hVHiWo0zNVuwvabEKhZYGsfIFbU71+eYLtmqWD4iMcVDwPvYBHxRD4E9yHyqV
p17Bb9b4FsWh9+pwWy+/Wtvi9j8RFgycQlAoGUoB8IjRYq0DB8R/wX9+Z6uefmj7pKbUYYVikgJE
g8149Cc8m2fFVyKQX1vOsFH46PrJd/1YZj5HDHvzItgQY3hdjCfPcfSPWhzxbgt02C8d01a78CCt
gJBe5uC9Aoj5B8P5+7gx7Twz7/9RbJxCnb0XWZLeIe81G12iKfzgj2ByDu3AYlkDcH7cZW8vwWGp
TzijqG9Ymk6AS7ZMpz018zTB2VIHK/WfxPcsBTvdG8MYQ/pqFMTxMg76MhgFaK/ImyELGEWMFMfO
yI4ChqYk2W5JOjzke1MOPr6JPlW0rkjlu3msxepJJRa7PSB+yYJtKhGPysnXHGJOH1MW2J9W7g6p
hfJujkcKyDTzitqZwMu4kb8j/qmE02aeAZyoqcUXE+cCvZiJLM8ekp6zZSco+Fs5PJPfkQbMurjo
5vBxDF0RkXFHgJMytHpmRA9kPMuX3LBe9l+HBYz9o9qVMDb+gk00KnX0yr7q8Wz0pOSTLU6MYP8r
zLT32dxS2IYS3qPGMP/pW14X64bWy71SquwjhQ5vbaPkdi1nJGqf9ln2lt2Jqb1DAHwUrk26dQT0
PxDtds98m7+6gr6MmB3RfRGFvxmxybY4UCakL95Yn2gw4QR4L667mcYHgiiJROLAXts1FDrxCkc/
e5e+BwogagprnjTTy/NuNlDEnuCykFWgnLsN50Z0sfppDVQm6UQn1RBbHb7e128Wl/m03obYHDpF
2Oe3FrbMoB8718eeIOPcpDHQx1BxJZ+EwwgztGQyiJpNqlCsTuavE+zNymDs6guZNnKMTDhUg2wh
HsGtzyKJgTSyD74QQRg6/NDWZU9i23RXocWgymhS3PuuRpLeVlR2gAELgCFTBtM94KSmz9J5or31
w5S9psYVzkhuXxVjQsuyewH3u1vf9qXt0mAbdr87EPRE26d1Ea/vez3SC1oKWd18NlN1Gttmx+O9
eBtZwu4lYMd/jOSp9lp2saor206FmC+jF+hEJt3Jcu0pgdoAUNLGviB3/aipfjmN93i0vSXr84eZ
Mg2MN6ImGgRzqw5kNe0aZ969wJ9IJNbmivccOYqhxzVLeRr2y25uOsmWewNjMLD26VH7r4r/SRqF
2lHoZZZloyuuZT2x53ImsAcPsnDhth+VBQ0s5ABBiZj7HznxwiuJTFGQS1+QnOsHon3wXAL5pdxi
0d109pVnIXB9PvLhEcTprk4QSPIK7CN32EYuVBY6lZASTP4De4npm0669tN9M5nncIOktOSicLV3
JbaJknQKSHPlKtnUD+Rb/zb6D80WWd+GBbFuX53ISCV0wFIwaVT9LOBzGqN0WmXZEjLrl0aOpSqL
NVP2kGpn6pCucrmfbOUEfptKTyxmamrFWXVuKlIds9Dn53GdyzIHW2F/4JfgA8oifXIWQBsgEdlI
3CToSbKi01xTWStpYaWari45nQ0PQrTsSdz9fa6nFNQbjKqcT03jAWPycowJfks4xFhfPcGIYFMP
ufnHV80mtb95/nETnH5lq0SpfQPpoDzwXW+Zw9hqaNu7ev3km3wqjERUGmfTnIe7QYhh5U2ZpFV2
4pDVPvbWwZsaC2Ar1PlL96Oq+eDS84NCOpdFE40HHYs+gcchFjwEaIVazzYEpCcVZh3PwXSgQFM7
SlWomEYAw/MiCkqTZwbtkTZyUx6yv4ZvAOXwoK//10WFEw+6fStZalfsc8vwK3zUfA4D2it7YhrR
r/JUbXkyvFIAuBWmwydfTXy8E+BCM3xaWNWzWb4TWh1dth0VbOOioEn42hneztOUTvW9jy1s2/St
Ep0BlUu1WKbaRnTIHfekTFXGG/iWo7HwVn27HdB/NQ9/+1oeX3I9NqBk63UshSXr6Qr4NyjekUih
nUdRT1Li7HdZCyDA7HQbzFjhVRsVklom//mBQE9BYTmJYtDc8Il01QcznMQVV2sQ2os87IT9CL4k
WyIJ7kxeEgBLVOMZAcka6goOvWQiGvw1wPO7SeEX7Dn/SsLhf5gkP42ixw/gLq+pf96OJoykxJoV
QqB7qnVQAYWKW2ylkizewI+ywWvVra2/kIax6uZPt2sCckrbKSHS7ee/YgMgAo/teS35EHBLKk1x
S4dK5dsfHqYtO4FdhbLguwhQGuZFvdHjLGtsOtLC0aUK8fOW+iP86zBQ2T1B1ghhS35pZMQtfw2y
E+Zcmm02ST8rceTslZWBKxvlpjrnjC6yUyvS00DBhLDGiQ65WcaWpZUEFchFx1mrfpFdr97IsO7d
sEnCsiee3BleILHeQYS3UeUwR6pkPHzeVc+OqUOOWJflbyqeBzTQ+eWjtfgr7KHk903Y2FGYHZDk
4yis3rnf+ggiiekP3QpK8DNe3kLKSBa24JGVmDBd7EhFYjP/W3wy/ls5vlvHrJ2VZkNUvPVPXVCZ
hESDFAApcqmBcNIgWdvEgMcyZjWyDLUzTxZx3hyQ7x1zsiTzXPIvyw/LX/ZU8nSeCOhFQeju5xWI
z4AbtU3h68X7+xfbFgn3cWGj4TXC+XnRaFq9N9qttFWGaag2hMwiFB5GWI9Kn1lFmLBMlMnWGdqZ
5VRl+Uw8vJGeU15/++PcH51ZSoK6VvTSRaGH7rJW77AEJyYXHTBVW5rbKD9rLvuOsLFZlz8/ti0W
vstTTRzcB8RliT9s/by8y+fkHbTvyedO3C3Pb15Lt+P4VzamY2YImKyBY/a12ie+NxK9TEdNzL1K
6pzNHug+IVxRk8Qhks24nbeSaqFxgyxCYyTjVNwrkFuUUDWS+JI3Pk915qyfvjk0oxyyEnumM2sH
YiTqJpY9ZNpZsy0uVdwFI52sgnB18SAPvbz+LFYbroaoDZ8nJDoPxYZ4vW2O5T5Oh4oWMB/MHQk/
EYk5isdoma/MdVRuKwq1AgmDjtkYvrL6SGSiykppLgNi3B2If6w0QUjAAc+PkKX6lEpVcPHtHyZ5
HWNAKAmrpDOeGJQLD6r0G6lr/YOjBSYysgQxAX+a6WkCQV5B4CPIBwUZobwf8kidjaEPko49Wp6O
a3a98vWr4WTOCfpfIDwozQiOOL4Tjq47WInjOPPtjdz0F5+coLtHqrN8jVxT4IWWgW5aDsgIXP/N
PkwrFRJcpfbmyWtFzEG71eMZxb3FtewNOvV1LV6FVEO0QOFzTe4YR9Colr7lXJhQqYCVi4q2kdtE
sRHWyI8oGiPf1pBWgU//JrwkOqzCDl6Q40oy4XddSkOh7c1XlXGYKUJTEcYqpAtEzwExB03ACT0f
o9rnRueJX4PyqvW2V8TUk/alZc4y+NKze0+toNlJnhFZCeY+PcDK0O7MT6l3Dd9FGi2uMOA0Rj+a
ni6xM8I45gGmmuZthHVcHm+KoN74pS/NH6PKbc8XbhFbmPgMkrSzL4wdyujfmOhQWiOtYJ1TVfat
KtFj53XTmv2nC2rCXegkqlIb4YGnZUxp0U7W2AqIwbZ2oQqFTgLIJa3WyhMgGI6FTc/xNK8HY2/G
7M1KwnVLIpzPPPCVQwA0/C5kUk9DTHO0wqbnOdGqvzISXu7KhL+3dYLXu7bW6TVQwsYD8k170mS0
HcBWB+SCC/Z2vlQqWHiyBGfzKXkCW6hrb2MrzqB0x8NHV9baGbYVOEACX+L6rAbofaDPdFXGhhKg
sXKTvgmM0WoFIHIx3jOUzBjQ2Qs1PT/e55H1UVNJcddMeUb+4UADQ47nnLlZLPsqeoqRE+PfrBfV
TFLgN9JAE66xEr3DiOxqVMNlfLWRZcS5WKFjrNumC5XaYVC/gGWlA7ahKR8LZRjNyp/fC74qMlcV
yIRve3KLQf9A/graYxLRj6zexL56bCxMVHkmGkk2H+2YTSuQDU38f/ybo34SMpO0pCOfwI27uSkS
iaCdC0eSCC55u8AjhdXOnmk7IsUtSSn3+TU4sg0KQml5UOhQHoMKvNLP3U4GqPp1+9/RqsiaGuYw
57KV0iVGfU/d5OP54bkhYNQwXltU4vtNbPs4Sy50kQ6kOrYilhXolnBBlz106uH2BZmViXJ1gGXv
JjpiQHxHEteGFNuGXq/hawYKkqkHOZFieRZ30sebYIIIf5KccI0crZEFumDUwlh2h4Mfr21Uw/hv
tldvcYILHpO+I2+mBjKQ09bYqwvvwNNR0BJ4HC9Vim51ffM5eatDlj2iFJ6nUobeVZF1juqrZfHp
O1af8Wfp+GVKsD/kEBjkCw00YfqHAIhizF8Iugjh912+B7M/Yrna4YQ6RqP3IKeRnKTYYpyHP0H9
cVlzAFB+QoSr6jyCMukMIyDUhJ30Scsf2f0V+uVu7iclF4tvg3SG1t2xs3J+w7pYcctInPiAIBZw
RZV5QeZEcYVD3CT96P8nML9S9X8cV+DvPdYkeEskVGsYMDSV7MOnZ2bCHDRqiI8r/M6oaGBgrCwl
e7CGYoulzWwyKHXcb7fBUPpXNSjgKxr/sB9L7OadtBBg4sTifxHzJtHEfEOq4+zSkf8QhjigkNZg
F1+XGzWJbRv863s38X9fvRarnqq/lfymAZ3xUOKT5tVXhWp0Zpy3MfunLwCeGl1ErvWpUcud8MmR
9JF3tGjD+k+UXHvBEKfkXV8GBIT5fau/x0KQ13QOEAr50z4xj9b80C78nd0tF9Depa8KcH13T0e7
oP5pT8cI6t+uy7dMHCqPmM0uFE2HJB7fY0rhZO27cGK8qL7equJegZm55IOe5i86ZV+af4wK69E8
sDFtuq3O+fD4+aV50daKpChplv9Z15hhFzWtfTNLdOoSKMm8L+Ltv5vVa0I3QqjDoHCI9BmhEKke
RYi6ptEBABvb8CijNdHNej2v/fdRaUsGTLM554N2i5iullEicYA+9ZhnKbvJ40vdejClBaVIvlKk
iIvtWz2B3UwXC1kUr7+zyxXWp5jf7Nlz8zFQfMLnuPjhvSW/7uGOICQ6oCKCCneBI0JY5Sh4n/aA
wSPh0wSib5/rxDnDdW8kjMzOPONmsJEBAvkQD96E2XMppT8zov0L4l1HEEYq4JBtz2Xo2EOUTlQz
Y1MlQ2aQjA8CWhdYSiUqa/u6ozMTGdX+0ux06LQWtV72v8UM6LGJHQGxfcTA7+8tFWVh1HqzQuhp
Irq+Eg7p69s+x0wDqMiU7I/Y8CNKycRgomWTlSGu7CTtecq2kHhPHmT8egCnWI4duocHJ5T0lf+0
MLhvZkZ5owq+ffQLJ54P3L3uirTJChlCUTaPnyf17JEfsCVfIArOQe9DPZjGAZc9JqjC5FuixXmJ
ZyFRVRRxGaFdjOYVPgsvAIiDWkWVAEJOfNrd0+v0Xtw0ncxkUu0i57pITxvksawivgRNe6Exn8oJ
i9oPnztnKWipxgYFITUazIf+1iKJeSJ+jIn7PFUz0CXR0hDd2g3nlGZ2pdkcxVcCxXKL2sQ95gHg
0ydhGiEDPL2z4iKVmsmY9ERzWLDOSl+5ZUgyxwuhF+s5UM7gI8Pq6nRTsKTjX9kgK0K3ebGtzArY
1GS1j8F/CI7E4FvtB3zFabSHjvJxeRB2BUtVNq+tD6PO0ZconUUIdGgbsQq4ZQGURtC3mYqkMR15
y6XykF1k68JlQlFrOZFOr58L+iYN8RJw4RdwKbAESM9nX2OFlqnsx3RAoYue4Dk3K6sXS5/p9tz9
qS6WcIzrVdY4R8hQmGIC5AKp89o59CN1m81jxurH5AcFP5FiQK40wLrUfDIik6rzVlVTzzyZc2fq
eXLafxBodcMfHUeSMpuF49QVy+vvi4H40MdSYjGdmKcft5ipeW+bOlePcNOlE5nTgB4yLb9qDYBe
TPnZfRCoTjZSJ1d4BmRaUKo/RN54cTpFPgkaz90UJUoVDHnoSgeTEtzwPuwkahX/b8obRHbx8Uk8
8rTFtvYQeD9krKtXuLfkDT9oAZ+aDhyphbPeDUqgftB54fUVUJT5ThDG+c77V0ZCEFI5hfa9DAs5
y2Re+fCJsQ0GnnLphiKEl/MvwU51riifdjIb2T8WXshHs6uG3AOGnPIZksvbsLBaphBXuYDVxFz6
K0XV+yNc68J59L+eXDIe2Man8SQ7+KCuH2Kzv9R76xWUCpFjQJ+/KmtGj2FNnSy59+s1DSko3EzG
tiKf8nWXDjE3b0p77z6OvwuGLZ1JbquaYrPYUlsowAwx3GXRxqKFIFH3KaJO/K+6ZmPScP2HMKM3
JHzpwHQsfV9hTxwLRxjuNTjdl+68/Qdp9Q6lONree0T536GY76jAqji9Pw3IJePRsoI+TIVjff7N
ZCSFRsJF5hFj3qjD6y6meTMk26U8QL3n0CF+bvVH3W4z5sDTQjqrVAIuGTCMB3yaRQCQD4PO1XTC
WjuuP7XqTRVgM9GsDhZzqLPRns8fpK/c8qtj7m1vTU9fGdSj2s8WWfXWzuymy33nHgXIPTNoNhqQ
zjR5DgoBoKtcz5Z6TX59EC7G0CKvCwFl7ZuKpC88UbkoaiwYU6ByiAL+bVcA59bvYv5srAVqfbzT
0ofLJkWLdUsMnEfZYt/mXt0JJuL2u3vAxvOsRTxcEcuiA+2uTCdofKtYmOiuVa9cHOlDnEDWtiyi
dl5Pc1J3phtaCc07yR8PexWwfZwlToaXauTll+MzI43iDv7h4pFBSGv5Ex50Z2Nt1AL3D/JhZyVq
csLTxdyIOg4yhb9Jbu4O8zJEO02YZcCiWIxCZMMa3icVeWEYkQuCERVBERM0UHHs3TMkU7HQMQfb
dywyFE6rPvKbhEkreWDxGk1AU3fi7T/RUtXXXMS8xvS+LBIkAb2dc0o4EQjV16IdfdVN4o2plSJ+
lEM1kvc9iEJKYFJACuSI5oQwyLH9gU3qUs1RVHmuPrJ8hANTf1UUoJ+rMF9tJ+d2/u49bYwVODP1
WhZcNfaFHy1h+0Y9YuU/jAxb7Q2KC+siV6IgYKj4mkorS5ANN7Rwkew5SgoTU1Q6MFnuguWtQDOU
akvoDu3UQN7iEMYBvZpSn4/ba264/Nw0uFWqOCXzc+siXfWDl6RBvNLA8L7/1lb4Pxtp/AAwxAbJ
qUR4t6ZWpUZpHxoekljpf98EVxoJswfa6ZK8Rqitidx96LCkFRY7buXLqTG0ZufNogA5IjHGSzqB
bcAbk3eFkwpIhL5iVthjKD+mP8h7HxoALoCv8+7QYNpixGwxHYnwhJDOHyGPM8nXEQncANrXh/Di
i/P7rhwwARcI4KIs4RRCjJDgwNIOccFbhklHEWbYcWBR7npolCUu9/DRCFShegOsMnDB/BWXH8x7
jcIEkScuan/KRGVV0U0Ag7eK7XFC/OpepEoaCu82JpMxijyRVqa8xfA0zYYd3TFVj6dEPFSBO3db
Li3IwIQuX/+6qSNJPEtQ20CD2Tes7gpeEhoHIHKqG2YxdqggBA6Gg2CNoLvs5kJof3vm3z0vv5bA
FIU5G6jIXVcc+dG+Pfn1wRwbbpGPjXyi7K1FdbXb9GeGsxtXHvIurq6T/lRTa4/MNQqYFY2d50/y
rqLIOUNzqIJ0/iE1kEUTWm496BH4SSni8IHvVFsacxXTWPNWHZ18+3VnvxZH8EC+4XmE/PbjBaVP
o516OcV1LEMI9iwHdegPIqk2ih+Y9P22NBNxQXKKUO2fOwnPboCJvdMgGyOrut9zAtJEpdQwmhNc
YSDv0mtsmWL1tJP7/5/0wcqLYPogq5+TNlQk4NMduGBHhH7mZeACSi5zA5XHn76cgVdDoTp7lw+d
9lz41SGjjAvi3bMbqqk2NpFaslLYj6CXdaCrVAUZXZvflM6A0Wq2G3W6C1+I47SUXdtAF1BJbpWH
KNz7f93PeeYbtqLUGvUJibac98H1qtVhHis+vlbYe6YF1qnwC3XPwRFaIjZJ3nZ9CjFWc4NDqXHE
Jy5vlJ8XaKk5NEyXmpoCjNnlmi85TpNdnvcLkyAPMdr8gRZ16pozSq675hIyZoxudKU/o1qxCbkZ
MnR6Pqxgcu9Lk1i46jk/0LtlZg+61pJ720qR8dmmn4k1TiIj0EoafYW53EQCKuzF9teAeJr+NeKy
feK889hVtoPjfK2ikuELYFTtCHTNDO1EDOpjRbCwaS9iw8qF86btMyLtIPNBM9ki1KQYtM6ZzoDF
0+0U0rzIFjv7X9/3QZTQ+Vwurht53+qXiySrUyVHNAWCuiaPI44aJsL0i56wJCgvaUXRBxKM7b9y
U4NK64ZfWEBkX6j1ct+RWfI3+MgPtpsdR30EJrF0UobS9mw6YkXO6mYUn6tS3bmexmyBra6tXSa5
bpYaeJrrI5AAb14J/+kib/Dz2T4yprIKPxPv1VMOe55nx1gC5lSQzbvZ4GvdUKpSDZnaOpT66WBj
00akDvP1g0yoeW6+5It4xx1jzVYS8pQOS/GdSLpMuffFwQCy94IptJELO1AVUsCONlksm8hLeJym
QebVm1hxPZB2OTxUbriP5hBGQQftCWyZNBq1Do1wNRslmq9qabHp17GWo2GQwj7fXAiX9fvKH/m8
cewk1cshFE/9OcHYYtGnIx2Rs6hbBQws57MVVr4Tz/t8awp9zpq2AoepqZ/HmT+1zunkuZ8gbTKE
ioF0MIHk8EJmeDnJvatbQaau87DItq+2S1klWJdyKNOuM+VICO21n8ObCejsmAKa182wSLHmBGXy
ztybvPHs4yNOYHB6foWCoP1PwBQTEuKGlz6a88C/XJmI5xMZsBLb87jycSWAtXjYe/GT9hnmc5RX
cBK9AATVw1vgCSbiBTn3XSp+ZcCm/DXaLd7dmvHBuSkCkDNYlnGKLpw+xc6oahe3e5ZJS5bWT8jK
sdu4U+LycaFjuquz9Yf1J5bd9bHJBpAhA7NAkUjiGLdK8+1mUnbYG7dNm4hsEbcO4buJwcMyzeT6
4LhcBIa4m5emmqjbO+nFhrJN/QUeQt9VDFpRAgb05hPlw8H+QDgOzQuKpUdYu78doY6vpyT3CTXu
fVWgS7yx/rkjIfv6/zzCzm6ioT9n/Qwru95uGdPb+/ufujZjiIJSWYjaKW1Rf66UFKpp07DlFCez
yl6pkX3ifdets85+iubGf7Y2Dr5wH4drS8OrRRq+okJYlQl0JLLVI/mP7DIKXtzATUimZCzC/xIo
ItUjIjiUN8pQKWdQ7jIPLp+cJc6O6YLrpNUbZ+PSgK7kuOi6lNlT1/UxtwUIsM9+Cb9PoxCj3V9e
qGaOGDjgdvjXcs50i5IWxtsjDCbvfjAA8dAjZoT4WkwBwURUatN5UbsjMjE3KPz6565EviR5y0fH
sJlQcFkPOhjH8bjj8HXTDE7FW5ormjLxkOwtsVEJKS8RO7n2Q4LUoXzggESsGMF6zCPNIUpUXh0W
/dij2QLNvZAFdd/SuwDgpCFdsnJeQcvA9h5VsLCV2rwlOzwIcBBCt/ksGa5yJH5OiF7G0SeOClVG
RLXbXakan2zJCpbgmIXudJr+Rplm1yQKSj72B/zmns0XaVfGRZhGQJ8sev1JmmEVfagnWuQegWfS
jxKq77/tNOjrvNY8oeT9lSwauXR6ulj/1pOyTBlTj8K+oGEdKR1h0um/tcMFNTCuMHItsrWC4Wbo
u4Zcmh5v9M5rGdMq4krXt5emccSjpTT+nx8H+kwVQPbdLOGsWkyoPMm4Tj5Z9wZSzwRRxfdfwdaZ
T44z40soMsX+Ji7/Nnt1kq8YT3A6zbSlPuhD27hbFWOtGTzi3BGgGMzbw9A1FsVFhJFgko5+U5ke
14I3ZGds+Z44qsp9wjKCauXW7KIlVjP5jYPHpQ15lD37Uz1nhBg/ZEQjvZrfUkt7BFqYmqMpmydg
jJYe/kuN9KWJkz8RwNcF/hLBRffjsgKYV4N7cJW2EiWot9XMFzh9KuJgbi3O/T5dh+4MMc/DA95o
ylIJhXBK5ZS/0rMPxl63KYMqs0Mnqp9vqs5wG+Vo0IF3AQ2Q4CVfMacbh1M0IM5ZOPSy4V54Gmv1
VZq2Xx34cxG9Rao8WpwiKFILiqivhJV9CEsRxLmyW27XqBMZJdA6uXElSLZn8d9CpwS3pc+vB+Mx
koZ/3pXFk9GVAVkE7+TcW5EBYM+Ont2zoO01y7OjiaAUuQ4HykC9uecVjz2t/8yo+Dlsv5rvlDwY
fu0ZbTOZvfJTzbcIATK1HgIiUUI8/YxzCayjzYp5tmVqxngNrkK9fNsV79j/OyQL6UJ/oIX7hZnr
aTzunHZu4tpBWyjZYlXNNgXPwWXidSPV1qgW9uPkthQxA0ZWBeV5LN/5gC5mFU0TQsozNwnHZF8s
vSxbOyJnAFB+KRrtAV+3NIyipEAk9P9+4AzeAUVS/He4IRGCvc4CbEuaGDAq2zl7gRGbxi4YBE9w
z02ZTt75tAomV01OA9LOAXMzUZsrDvgKJp3RDkv+mJIsUu3/SkKXZakxsGZl0ge6ynipI8LjjTZH
kUyEBe7LT06ShWT7pyOlNGUEglDStD8ul/Bsb/YEyp+g9Hyw6/3oiJzoXJsxULTra7lgZtEtqIUv
+56rdUzl3+Zxcim8DxbdH2C6582pqQfSQOV4iQuQTWoxIeGbD2lWbFTKViUb5dLUeCIvkXphbiGg
CDsPLWkIXeUWfz1vNdqPWAqGGVip1/b+oTrrDKuS/Iik/k5RA9UuyhKgoUMnDgKkYtftVQlAMF76
zIcfDS7a0e6LnRdyOPggS4kTFKqe8nT6ihA+uQunGk5OkR8XyHrAtpF+Sdmadu9fUi72xLkIfT6j
gpZLAx3thijf4vAGg6UWl/+ijQFMNxFMATw4No/NCmhJkoBpLa1v0gDM4pWda3Zo4R7/YdLqIP43
adn5UOL8ka/JjS0VRnhR4lCoOh7Mo1NATO+k6fAs7AsSh+Nq1voFKZ61YEW4NbExpsCwmwKsQn/V
coOcv/lCFzwtjE6CHmu9OL44jOmTFgT+kiqrx/aEkP8tnPZOv677oS0C7Ra+i4B0yg9AL6E5ir0i
9oreqhh/hMXbTgXbwy/t1wrzOSl5obN1J2mbxB+HyzJpn7/FbH2aBXDi5lD9ox/suRjdwaTUOE7j
g5DMoo06zKKXtc1Kp7PjHa/tP4tZvavQpHlZWYHwi3D259m++4IdG/+ha6tYPLdDj+dEMT2kLmqr
lXxDAUOoGZ4bGvVKRaAliT6f48uac6iMZp7bj70mZSWgX81ml5M1R4QKoA9qrF+VPaJI68PtkUoR
QgaPn1y/vEr5hvHCYM02kl70wcIiAwoUGe1eZHF1+3GuwprcPFsD7UTHjAfOlwL7V1GKeYWsstC4
Rx0Lx0MM/8YG+TBAgjkItv3tQZt8D3bRlVgbKWI+BrxETqTeL6xCIKr+9lUkGcsJaL95XtIzCUAn
RK7IdupK02yQod2fzHNdUhmiz8G6OHzNCipQyeg1PvWrRSlgZQptHAaWu8qFQ5fCL+MrECc8Mt0H
HSeMv+JkDL2vWt6e6IziYD6UAZ8mKjwlbX6UP0Im/RBJfDZtdesxJwT7on7B6B5JA9m3dUcW+EW4
bTK9FEWHKLGBZWxLfPvlq1fihy1vUEO/pJedgouc7Z3Pih+smidK+FG0xIbFidxVi1FuYQKPUX74
febsraIqhuvaz4C23GqnICn0S7ZusQ4hEEeVQ+qrg74AOluWKYYRZeN4VpQ2Fpy/nj7wpuz30Ul5
EzwiqZFJrlVWPCVChM5ol8nn8GTo0n/De/iIthgkO8uIjbDhmvYpi/AOZEkuR1zhi36vmlTIzXEw
z7cwTY5Ie1Dt5q54P6MdCbjoVm13tdgrkRVmM30ibNasgBSLD/vwPhP01YfTUu8ZO3MXZ9IguivX
t1xGHwxKCjDKNsOOB2XCTRBh0vKPRUh0XatPmXj3zhlAHHtjyBdNekKBsZs6L7wdYrXj8qC2PeCI
E+F8a2HH0ae2hridFGfec1N6wqOMlFE9uQA2NWggsMqTy7EP/HksXTCHFJj61XI9skB25pkxKnCf
qVwbBLQZ7iOVm74kPrs1IQnHATJRCb3fxYcGw+jtSs1Vbxx4mc8FSRfAUCO+0VD4meY+f8GQq5ZZ
qYiy7vk1nuxcCo87/30J4WEXvPQei6KbTnUrNGUR8kx4DtT3MH+7kmaxBi9UMWRCkH0mDk/WVsy0
AwHpSSglddupy/f192kZltcGsJnLYJYwjILGCQ/YYY8wXwrDbDUupwJu02TWAuxQmqSje7KX/fx2
2oSRibF5777f6pnWBK4r5dxoJw5jhYYzASyMFOYdGw0++BQW/JjNGkzH38dbHOfUVTi1+/On6Kya
JZZEiFm7zGuUD5JSZXLvq6neKCLH611Tk5FoYJv9JiQOLSvGqViP7CQ2u0Tz6J1JSHNNuFS7WR9G
7huvcbw4kQySr8nun8Gs+ch6LD8peQ/tR1blZoKslDxiKO+LPDi5hwNIwp08n1565TP76dm/D8ax
KX4QMASdr7++NSPdVxgXq7ap0hX9auSkxSecWNTFt3s+z4jZ6w3gP/BSmbz7iXqSsJV3SvhYY/iP
ZsQLMMgFEiQaep43+1mZDC6e1jryFie1UnyqgqvhgaICYmDrZ7qFvaWFEeXKYhuMERJUm/O/P2TO
19w1rezTgeGsFY2tvWxQw9tffmI6aAXE3oXG4hApnpDHbZj5Ivj3y4VA0rO1ExN5NqzZ9Hy+pBJP
a/57bhfTMnbAkGJ8S3I7G8CEbm8oqF45WH2u2Oqus81GzuwNaMuW/65PLWOOxAVeMg3f4XVicAza
NAbdyvJbS1WDkvIOXrJVY7zU9VhHVsglMjD7aeT/MUQSxKQPZOmBQxfFo+vKMwozt9QhzQqsXu0b
selu8O8rJshxn4mZcLf/y3AX1JKN6ADL2hro+otF8uZs+vG56DfqCoH6wQszewwToRdwcQ61Aqtq
gafrrSrw69wJGQ+Bq0sQ5HVyEIa8J9lnepYmkFQjTCtMEVFSpHg+KdZcopRoCzhUm8yxW8o/MZLB
lWuMStpvvCm0d95XMhMvFSuDgjlFpeYQrAk7Bn900yEOIiQKImr7beyR6ROIhAWF2910Rjaj3B9g
JUkOrX9Xbe3W7aFGwM93NjowELVYviRXVcsqF0Z8nKfCT7YB0RUM7mHcFnaDMQJyM5wBWSGeUo0Z
HloNW1VjpHaUTHMUNWiOy/NOoPgJ7SoCrFa6xShQyUAdVeq6PMVpIh1+G1mPBhQI3mLnZduCWhOU
Y0DIVL9OsirqB61HZxOW8kZaXF4yhmpy2i3fM8+p6vQbcerEDAyUIRPiQWbkHIvfXlp9RFfYHIrw
SIzYvrzqjzKRgATQ7zHp5L9yDBAthttO03GIhantS5uGnA6FbmqCQgWGxbbluAlAeZS6Qnyt92aF
89hXaCSZ8ruRNxFwT5nDRS/XOsNwTCR5KuwGCtIsW29ta3sihKY/lzppr4fE6aHgL/PltJs12UWY
Sug8wVMQilQm4kEfWm2Pi3jk9CD+ARyAEv8qaeNsnD+XqH2OtzXyXJdKL5GW9KfICgKhzWEuCCea
L3ixI2qXg+FZiDtVmVEtT7VVP2v/JjNDgw5BHBAcTojcHn5OC168YotQNNUZWmZq1dDVyox4FRoi
mliTOK6b7LnXnDCiPo9LR1mmfk7J/kRw8i9IuMM4PL9ffjRlenVrI7xbGztAGeb0OWqRque+KnFM
qXbwdfycePqGHlgb5ExG+2YLpywOi2hhj+mK5PmG+MoM8S3hDuhZZYfmo2p3EcSrV42bPdSiuPDF
sy4IP0qTyrOX1DeyrKMXaUEUK8MQW9haS7LmuMJ4tXq8xi/ZWI3jJXIW5jp/r20RL/lHrb0MshhV
6/YTkQKiyBYEfQ5RfyzjpC/buBe47Lu5RCNgSdYwkYXHEmfAixgbWpEc6cV2wV9iVdB3vRDdN61Z
7cUF4TqirmavAYGR4z9F4vRzWiDC8H45VtEjqThbmWF+M0L38f/iolKg4HoejCxstIYw0c4EvxqT
uRWxjMWvRbHKP1bkoGnx0qRMs/QeU2t2p18qA0UyVrCGWE7rLZBSzHCz04ViTl5kDb7BL7mcNVJB
fOFvM8mtVi2k0TTODpWxz2Iv6EfXba82GunNzQuBngjVcrQOWlPsEcs8ReRJwYxEqD1qMd/tRqFq
IZ/vXJpJM8poLAYw4/9K2x4vMG6ghDQ/N5eOBDcQU0hF7tRcM6Qv8vfata7xM+6ARiqvxITceZlK
QGLtsX6mj1QO2IuYS89uFtlwMBe2o44oZV9jbgONQ415fvInqebS6PgLI1Pn2hDPrvqcD8WsfKdp
IN+UnskvBWKLzaQIX5U7nN43OVje9OBz4EfGP3WddHv4DE2pr2WDxzW70qX/yViF9JderPjvJgUL
6JCmCY4ppZ1NpWc4cOJEA+SD+acuSwG1ia02PbEkIlOvXjBotyZIAylKRnVSaZqP9F1ClVkO/cMA
kx69BH8INIwSLIdgHah78KlKgoGvipccEaWwuBm9WC3d0TjeFr5I0CbhpDHvg0fCyvMfyUCIL6Hz
zvOtkOD6sR14pLZnRRKagEdemlLvSmgmpYd6meqHifEZEqmB+XveKA/Z/DarUIdtXfy9oWTyDiYW
8S0D+ZeMVYpgu9RFBG0RX5aEO+c3aV26kJLjcMtuAdED5VW3jCRBqizm2hdMZvAMUZkfPNd2cSx1
TS9R/Nz8KRDMNWjJ/7bw78nJqDKOcQ88ooR4gqeyrjF+Rdn20RrKmnQ9iUZq9tulLgcXqzT/O1Dw
QZdmB6V8Q+LobdAaybF5gWlZGFvsn8YzKs0Es3I2he+hGmVN3C5xk8k17ziKfzCuyjUr9wOOiZNH
hyAImx8foAlAqLSkeKPFdWHerufoYTHaL9QrJ/znXjOOH0hLUTJC3DCRgA9frAptlrEygMrlIdwJ
cCj/4nSm9/1Gv5Yqa9QDCg4AKAaxM5KDiMD1NEZOpE23KVTPUcPEMbrCr3mk+ODneqdc1+jPsiQF
4lRMr4lRQPMuf+zzSnmnnOhLu1wa/rj/4dO7zZHJat1UIGlXcL3bo88ne6iOtcQF9OAFcqwwWIM8
+EwKwSbHzEzho+0rqRlrrWZjLUTCHawIPDbad8dX8M3vA/u08fjPCQXUSXI3JvMb6TTOgon72+mn
yRnjE5xE4ufAyKaxYOfg40QEnQyAoPDPrZOry06sV6UB0vS+C1Ggd5CQsaCJOwaaDKhNumDDI6zB
vkTJ2TWh+4S92qa6uI94CC5RbXdt0TWm8slUusEHNbbvy19LWV1YW6a7zaqcaigpcj4sFJMGdmnH
Meejgbi+wbeH4aJ1Eyqjfz+ieK2c0fglH7mqikPCsPSPqlOB++rNtFp/hVGAtv8Rp4XoH1g0Y+fE
k1SAH3ialU/G1ToFkIsu6f8nLmceNTZrYkt0Vir/OK3yRLZUW39D9kXKQS/aEqbj1WYFjMP6OiSV
gUClRIBHr4XMXWOWrL4TR2zMJeIjgJ+VgKSV4ZvH5+EfA4zqFnff3alhZLx5AQkJBfd9H5l4IrgA
5VTPp49Zq+Y6FezkcPnqus84wHEskiZu92zZ6XsLESrv1wiwg6DD5DwHnfKNVFydQcN41W2A1aOf
LU/yEj+TQTpg1HaVjD6Wb/I74dowU01luN1iyio3F4X1gg+/8CzbU/iHO3fVhzW3Bq7bng6CYBZ6
mohWU4A0umbp7x04wJBqCsh0vb91BiGvPyt0Icys/8Tfg/Ce353zcvYEO4tGvcS7lknkcsvEh3Yh
A2P/yObfK40ukX4xN9XK3QymWSQhbjC2Z0On0mY0CNSA4KaexIm+PicjyDoMn5OFu9WJuAWV+5ZY
qMS1BRLX+1+8SvfOJCOzigE40SfFMsuKO5YBNc2gAhkjN3GataeKAPkXjUB8Sz81fZdCR3gu4138
rTK6DVrvFzaxgmxN6bOvp1GVrA2Tc27gztY0FLAAcXVyDrLniO8HiPAhUrDB+jJJbi5gK/xiT+Sw
hzkB2bF3izovRbf93g9tbdiAqfGJfIvDXDW+fTkwseTHsGLefPSK9Qv57tzF1js1+w6nljL9ts+l
n3vJq/WbIeAZYsfwAeZ08qv7sRvrcWP7EckrHo9tx7cQc9bD4MXGQ+0GtlobqEN7aE/dcEzlazh0
of0Y4XhKEj8ZGaKu8N8kIe5J2i+G7QvoJWh0yv1Xz14LaA5y3GhOFy6VZW+qJLZvjVfik54pUV9u
pgwQ8o95fK2atucjQ95fThNXDAEe9QAAwdcfvelHzF5Q4tKqmf+hBcY8R1sYqLs3SC7ozn83azso
Q+4ImEaRHQnJFSdD1FYrRSiefeZuIsxdGv0OIpRLDwBjaP0tfG5cajBSNMfCqnRTHQtXQ3K/xrAb
Pf5a8SNUSn/JXfJxmflfSvW4wbGL30s757nf3qxt2OrJj2SmNyFxD0Vq5oCZf5uozrS5+zAqIKli
RfOvuD6eg6KhWNqHQa3IlKrSxSK5xpgTbJE8IcVmFkMtEyQt0DzGhl/dlq1svTjY2SaTpIv6RRga
L5jxeru2ygC62OYkYS//A85anYRKtcvaT4YM/vnEygUw+LcNRk8wNg8pfP4z4n26GGQsr8aZjMvy
23UQQr5GI1QBEm/Rr0DcvFxdQJWFovFWa423w8Us625oC1XyXMk8bVUH11eUOAkwetEF+m7OVHlh
4yBMklLIhW+uO/QexOWKBJdEmN1ndhmMn/4FLE4vUqlHSulYCjvjya1OHiyo90oAyT8tizCUjP2W
7G1rS7rUSf0EsuxeQ17EK9vyYsFVlprw7uRgA0uPrd0zSksg1Wry1+sxUCTVCIZ+Ypxu2iz0EXn1
UKVcx2lnT9UtXeEpkeH/OL62sdqBYXB7S4Id3DdmCjZi9jPP6/HCVePPWoCOZXGpJ4Kh60pkfUOG
ftHuNimBeG7re53IXlUHDoYc0DnLEPaYqiNP8gJt5H3bnXVX62mq9970rzZ1MxuVTWaLvN+bqIcp
Q8l13S/3fyoGnBbUb5HMtOUXAJ0MbKlV4Q5m4elpdX8dXPzdq+FQhTI+Nqw5pL2lxXfs+Z/NBnq1
LTSi905EJ/61xovk27o92hTdMpIArrFBBpFSfUqVj8dv41OJoenPM9pDCfnU/7sf/zAjJavRNdR0
83yNeVJsZETfh0/VqaKSxoDL1un1gb7gEreJVBK4qLfvxMesz0XGkNM7UwSiboUvYZQ2FaGg/U3k
IWT0cdfePQfz6bcQycOy7rTCr/Ud+IgcK4gjuaUj5qWNZdMTWywvtcSHzd0U1jVCXgIFyIanEpHf
Ojxwxc/4pdBxro/0kUudXaETCbxY5eMzwJqeCAmUjAvRMVYFSe3K6LmmUrlmZvZ9+h+Cg+i8EtDP
qeJgwbLfPKCBT8XHHWtXuScPyUqg64yb9/FpjdcHkBaXdSXT/AyUtRSFI7LLG2F+pgFdmenJrdRa
c8Kkh831qjhNxRPTRniMFJar035U1jUyfabsPK9WhFma2VK1lx7CGrF9ui/G10Bf5Z68eOqsRjA6
DCQacJUVyhUvhHXBf//IJ8f8IsUcYAt67w87HJMyXXyw7qy/QZetXVH5z4EKmLanxrpr8DZVMeHS
dhx90B/TwSeHuof4kVBHzgqEN8PRfsNlGY5I3w0HHeJvPUoGKuifuvIwZF0MBv98dYepxHSXmmQP
rnKRqzZDBJk3HGRJVpzKR4bog4CZJ3VGwaTRsp+MV760vKtackx2FP455iTgknUEouGsPyTeC6s3
o8C4vM9mSbnyRDbPZXxmqr5qU1UQ6u7ipwFND5yl2wHMFWh5CuyCH2dg0aIXuQpU1zOoUxQK9gUA
hQ4/hgdXs9R4nPB7lJnHsa9VYwEVxjzoAVEbOYbCO29C0lsbKU1rBPZdR+a4Iakuq1H/l7HcdpLd
jQOznnAYiSRl9aGjC0cQPP4AIG/0y7yAPuQSIF+dzM/QVTDwyrU4knzmxwRFMQ0UT3hWzPf2B1tw
pjazAsjIafAveLU0WyqPRYVBBwj/W0nHPrDOFd+Gno3GbGkGP3cWd4VHa1Jymtt0qr0sogmP8J4P
noNpMUADiPSnyeYqbWW8yEOrWL85Jw2a164JVnDmx9qB06FMc5s7VPBmFM/v2k31EwYNprywcwvo
tj2uI40kc6AY8eXu+3X88HXrG4OG4LM6VZpUj+8zkv4C7M0S5KGiRJB7G7K9YyB9vRQbT196l7YT
1g5d2YcKN84wXDp4wlFNLg7vZujQ3yJheiTYkMFHbdlJr+IaJ7J1J93ZAnKh13p0C3MHzeGUmHN4
iv0L87/HwxKLFp3hBKcUbyVVSiTq3yP6vJxIlsOwlSawzKlMNUJIrZ7raJiWpBuIEz/X+KsQfcTR
5i8DdktDIlNX4sw13ttE9ABxsindfoLStYYNKD/Dm06SjAU1bax7vKlISc00mMHwNput+h1V3lYI
zVNGbOo87IxnbsmDXkHG7jqP1iHmSmnrWKkmMpboeLSyxBZaul6NyiSt734N9DUHgXFfUwQbx//m
umHdm+EKfKeyXX8FLCfTzPCd7EfLqTfoKP467M7EW59+MXjs0n7IeLbCufLltzFPsp+4DstBUyGY
h5cI/RkLWbroiKs0q0Yh4Zif73bdLA3CSRXWBTmLfgwYXGaiEZgVwhEoyMpTGyfDmJgBSNoONWBd
Rh6wM6m84aN8Dhqr7fEaPdB5+eoKurS/s0UcrTTPu7DhzSeotFfSrJ2ahrTFG3/yeyLK3+r7Hsfy
SejgzTCgtPpZI8XgE8MoxPw4KB4PP0bv9+dRSkO23o+BPQ/BAZJUeEBZl5ugp97ZqSE3dL9dnGwv
L7gO+uIh8RsAA07xoCdj62e9y/cCYGC8Hr5kuF9DyR02l1dUdpwAMmlx0fzRjNkyXgZepFCuQVc8
mt0lzyEX+7ljTqSs5u6HywTRKjWEQvp5lFMsDB7GpV0XIZ5ANv430z450+ijdQJ3Ec0HGk6vdt3n
XFCsoSv9E6sqmLVPcClbFQnyIf2U8wme2gRwoJhUPxCnSfA9cI72z2YoXE5qvzzGxj+MKWnn4Vdz
Z96UP64W51fqop5BWuaE3WJHj2dvxDeOnca/aL+JPcw2Tkv7FSTeO1HRQqjhH22nHaPA4RWR3Nlu
dbkaZXAvJv4itEBbUlK5PiVoiD5PmR/tHN1EiaoVgQd28iYebxZcZc0fStuCql8sV6h6Jkv5BqZQ
5xhvB2jkQkLkLMhQI66yVIaeBMbsSbC58oq1s6K9WPdkNO9dbdXvef29nSJ0n9LGk1vOPb7uVh3E
b7Nt9HZAez/9MDWr7XBGK34r1pI8g8x3VdgYx+csg8EbUb8lEe+KLEQOlhCLw3SUs9amCzOqZgJx
1Awed8WabRuAoUSOh4x0XOOwZWESO9XTte5S9FJbN6UDw0Q7rH7IAmfk+UYvdXf8uz4pyElgSiq0
iiL/UsozioLDw/zGqgFFX0WeinswZaH/mRgy7d3GxZ7Ijm8xXT95dZBOHiiPsTwAHDIuLEX67nDV
9md2yKscJNz+4UhWiivff5E6U0XhEHSfugamHpJKydR6BJUTeSkNKRXvZWR85sRQAR7ejTkxXdeV
29UyEHTI87ux51GT9PcxuK7K4/pH4Q56t9uu3QQ4OgmC9eO52GIVRULpVFZFd5t7372eiRK48Bul
AFwA9lE68LkF4P7NnvP69LE4+saelGuOdvLkFL6i+OE+RCiw66PTA2XjmParRbANM1oci87Z5Z3G
WY8mGyEm2j1eJeaHPCH5TqYAoCpzCZf39MNzrlciW7NvP+r/n2Nzpdy8CdL2oZqiMJYv2ZnJdf0h
WwEs8ZAElaQGGj+KuoVeBFkevprlNGmOl2XIyMT+FdvG0RaZ7jTdmVkF5FWoBfqiePQFEmYi8Ujb
V1QSXhIsZqH/ZjSyl9hHFGXrvo+7LKtcDW+4DZsTnMlKV62b2XWb1D4mgMS4hUSyZw9cp3Hsr5lp
AlkCR2pBLsYSiJ+6PMmlOxmI486s8Ubjaef39XcB3ynGDEE8S6ympjbmvVgdGOph+ePWr1tmLMa5
0OD4vh22qitMZ2qBIRIq2aIQv3d4rO99oDOwop7pzquZ78Hrbgc+RggOksP2Gd4+5GbI4/QEvBb8
ADdIJ76QQ/2SjrLvMout1qsH+UGhGMyB2IAhN+x7EzE9255hJUfMwHOgxm2fMYTO7aPyL8Ce+hX0
FcthZYgtiSLSDFuhb/geMmbiG9jo2X2sSluIFCA0duZA4Je33n/dDobKchEaVBmufHmuSUJBvtJS
03I0KRAhngjD4qKSje9AdbSA+kXjsM75l/D0MJ4zyTAC6PlfbXq9FsSFCVyWhNyfr5GuH6S02qPe
1WrE0FuCHfDgOEIa/gfVVyHDQkgeuIdpHt3kuKi3WZjUxBsRC/uDcwURG5t47Z3L/xisPdpeJrTy
qKOmyIR+wz08MtLW4bRm3Fuc1b7jaUWgLf4U4XvshS6YJyhKHiE29/b7mvU5SmXP07ZQfJlsz/JB
ADih/gLfxhzQ6MGLWAZULsbHRXO01cMR0EyvnHsBuN2ZRsiUoS/fU5d3FmfiUlDsToWOjCT+HT1H
4o97b3va6w7ROhurjSv0B2plV8AzSG6bfoUYNFMYghT6ma2yMGneu7ltifoyIiYHZBGEFUMHICOK
R9KBPNwCTYvS/sBJSFa88gWDajmqDcYr4JedObsMkRKKq7UMMt6E9I7cMAKZORsajd1SQB0TuT5I
pJdLYYh94rEIhljf2+teuVf9CYTlID7OHyqVkO3BW1i5wPZk8vVfMfvIjNul6cJwlgU7YfCsoQIm
pE4lUm3Jurl86YiSX5uP1j4I6Ebzg8cBUtbqjgwUQe2JCfU2x7ebPVeuH89c5Ej+myqsxW5S8zeB
wN1lGAeeQ6xUJsq60PPJxztBX1lapyoDI0WBaVIMhuoXInPMWVOHQIrj4/3UWeTaqqclVSBPj3iJ
GJVZsiJqNiNHOVf0K/LiIHLzgBFWE2hT1+mEpV4AiUeYRKSZ70i8gGOuhI5be0bAzeZNCtOVPXbC
tEzh32KPf1j1DtKo7rKyS81CJK5CBq1Tnhb5Cw6IzhhNtNeMH/R2rjqusv4jtq841PuD8v9QgCT9
ihengOkRyC7UZbj3VTnECAH3zbb+Cvlxla+eMTe/W4QqlYMQmDhVZgM3i9bi2ygy1tNSi4FKDpfz
Z9G10sgDJqAiSCzy/deK9eVBCsPclcIN6Nowdzgd6iL0y+2B6wVIP6vSOCjRvQHAbppV+JD90UP1
xQn6yHQLh680VohDCcP2Sa4fhUyTnkKCseuy/2n5I6B+VKmkQtBnk/zf71gz38G4mJzlH36ojsyh
c0WJvfkGjI52OMaHqAeLk8lnpDkZPRkvvxULxS2abofs1Vn/jtAPJyT7PQdi4wk9MnmlOBC+kEIx
+GELEsEIJdHue3PMjkAxvJGWXGW2aaV4B93EtKbc1TCx0i+qCqJv+7YiqOycRHh9Dfiil1CZzIyC
tzxFmPnAoMvwQcqvZ83gYzbzhDW5UKN/TzApW1e347mij4FnDzBRiwP4Su/XPKaSVbl7yQx5IARN
KDPI/qtBUJN0mrZwyipxBpBZkdlN+kw3ZxFlpji5kDy8MBwIzVqb0xl7moj2usNklnbivWAANKo0
Ch3YS4bWcbhC4Gr8ilfwdpp0zIdAo60JnOeHTEGoAeVd/+Ca9kp0x7fapgyxT1neDB8NyP1LB/rL
SEk+JSXtAooo5WfrjPt/TLkgpZQ8tnUCLSa+mSgbfAd12G4NRWMdsEb+fNtX/DA0vMPmhCJ736s/
zbTr2tmqScTjot2IFOmEIjDRxcBsf4dQv4XGqCIe708rYU08nFU8GSuBmhyueT2nWZ/1x+XeULbx
LBRInM0+A67yocuko38AkzcIdWBEmxnOodqoeptsrE6g1pRHmiZfCjpadtdhZOc0pZqVlQqjMeL1
40GT1PbFv1weJ+YrKIVtlQ4sEduu1NkYAjXMw677bOBBBNSJ15e76Aj0w3q77jLk5ZwfrDkaVqAy
49+ajIZ5qe666U4zs/kYHJNqQZB785um8uKASez/ujs8fHgwHPtL/uGMg2V3C7Esg98O21z1UZXR
Si1JHRXdlBg5R4RT6qtMfAs5RO2FvaAySg2DpT+86CA893VaMtOcVPIp+HN0ZYXVLkutnGxMof4G
G+85Jmuj16khV3+j53aAtrtHHO5NfVTw+Z0CJ4W6iyt2Vykew0Qzdj7FQ1qRbnHqTvrgv5gGDmaQ
lE2x/vlqAqrin5FbiN4dLytJatz9LieXeVTbJ/KNRpw4aK7Tzcvjg58LByLAMdQ+qkLVM3BIoNWQ
CuOF+9nHAyBX4YHvD4psqAk3jxqichXkb+tJt/Re+PaGN/4k4cqB+YBYWBuZCGmDcPG/UIoFFtzN
l8cHswt+//i1UgDNMtH5CJzUTlDPKwkgMP6YS7X/0A20Yqt5Q+M0cmNdY19+90deYqQeCnPfE7BH
598HUUtmfqc3zBnH+yA1Iq4nC+jJDtuIL78GZOJ1+EXHHi45iCqoVHUUUBU4CLwMrXHnEDI0KqZm
Set9KexHoTqLVewtVfmNV3RkXraWFEm9b9RtmzEu3zcCsxHzj+BxQSS0jxpl3bRs67r5+40oxJ4M
AdCOiMFn7gd5xUzIblqD5cId1A880XlycJB0Mb08nxwOHqyP4W3hEZjNc0YnMIZ3wdmPZfs0aPqe
wAmf23a0jdWxW8bk4CRkkfR/QzoOQmQL+RVL593Hl//7iveKxx+EIPBfz65B2YdlLpn/mLt/+g1E
bPKGFGT+XxBNeRUmK4E8voY+IRLWMlmHUsKNEzqG8Q0TmRk1Bu3xqNmM+gSprlvZgaR9nTQjlp36
uLNEzRYonA2aFfmoH366qngkeFlJ+y/huKC1OZhSGEhD//mwxZpCjx+KxKUhdwqkoxZvavhtGWaW
3OusxBWRvE/JVwufTUry9+7avRqaVgEOk55tiISUcSwH7u0q6ELI8YKdePlMHmHfUM49ne/xx2V/
9I6AFxZoX3Qq+LwE4JqxHjFmzRsNvsGDicq+mPiIBeKJn54OouCDgX4wf4n75ETiNx5ZUcdWzTcA
EfUF9zVANmpz2R6PiI8VwHg3bplGKQ6IWiv/xchUk96KnWc0DQkF1E3sjR4mNaMT7Dv8VZZdU+gt
REkUt6hEU376iYpjcyk+O4gnuptUGpUZF45uGjbdk/EUwALLwF47NzWI/0W8uQbFg+x/5EZvGdBS
mT2t+wb4VnZl8zEGT+0OVduAtqL6mrGOr7LBgoTxDPM7tY3FcWMnU+UPWmuM1Ub8MauqG5V0O2is
2XFrueb2pmIVYlzZN6RPFD+E23zyX93rV+y5aSfFNM/KwS0/z1hkW685licKCCis/OpfJtgkcxnh
84d3nyD7SSA9qQmebZXPKyaO3/JotLOrELRkhreYieewpvApWvpunPuO4MudBrzuPjkGLkLhnF18
pE47hKbbG5ePAmrlK1TpQMSdnusrBgvAGH+TS1iPzZQswyy+dXJWCR+u/klhDHuIU8ghxSU5dI/4
gDCt2IkeUeZKiZbP9W4FeI70/nMgXPVdWvRzCbp6JPpqESfCb91HX/sWvHizOSu6VgOl5jjDS8Q6
+sauFASBoIaGDL0xoy/xN9L2Pfii6K4sDieIYXjS7YY/gn7+UUYamvsDx6EgIumbfQcLs2L2pKUK
wxqLqmUi6cwaoomixT9Kv5FgC1nSQ2JWFp0GOHhYsaUv6/JQzluYMm4cPluLZPUw/OxiLK1TGf69
EDr9bGLWlU+197g3/xviG0Qq4GRLfrqRtYXRTjspQ2oWKgMCbemi5VFphAIEP7KrLNlZWcu/pTRa
O2pazL4BPIa2epfNRoYlF+WMUr9UCDiDSq+dztTYIFqH2a7ICacbOVE7loln3/ox3fM3ShWlk+xK
rEIOijqC6lcC0fhYXUvBEPMBIjs2jW1L1WUnct6CT+nX3PbBeImvtVIaGBNEHQyOIV9L4UmEXr8Q
atUlanpEdMr9mD+FhPEzZU1uIPb8xpVwCjJrRxTLko5xvBnn9csduI0diUc8ZI23z1Llx5LhfaGC
w6+Nw5N0WZQI6mpRicGd+YukewldeGS4JwfzUefywKatQ5OimCi1+sE4nEXCUzP9tH4hCuif0B2A
Xb9kaWnd1A8Mnk75dTvrqOS8C3T6ro6x/Qe2XbHpfbixJY148WzCpjOOR1Y/xwPtOpwKEGupj5L+
DFPDHRVREn8Xjvj8uzQkhgo3x4OKskVWY5OuGyF/dMKV5ILb6KzquqN8TTr1hCOBU2XqwpBUYj+J
ISpSDudVswm14+Y9W65om6F75CmgvivrhTP+YH5dSURU0s2Ne8ZzKHzSuaEOkQCXclWkh6yInsu2
8TtXTMjcXNZo2QNAaYpD0Bx+Ycb6laEUspo9VkbIbCNGqJIFlq17IBs2g+DX0d8kSfGGXeT8eccD
+E7PPQhxqoYqy7maCy62dVS/gbUhPYI4U6uu4LN4Mt4BeRTGGStb97n23y9JCLRfXQ3tp7c0SErc
uwwwAeC/X2DnQQjRqLpQzxsKQ/b8B95kJ8fDgDr6F11w1ePsPfzH86CJeCnSQboL55UkNJLvV7QQ
3YDKY3V4ji0t9Fk0mydjI/buZXkw7EnSrt76VUcfs5ZDrMK5ooA4+agpzFA5QFU7vLZmNcn5IGkn
XGnPRvNuNH+kOxd2XO7KOrGzqmsV4ZLo3JTfT1JUZvLe5RAWWlYyNtBwjZSx2TXUdiRo7c7zlBwl
d30Hu0T6Xo5OWjDMKL2Uy6yCXh5E4WOmrzVMgWGE6mW/k/lZTjkVF/edkhSFuHSdCThOojbQ+7K4
OTPMiyn0KAQfl6TZLd2QV1TKtRM8S3nKpd5j9XwwPvHn5CBM26h5kbQfD3Lg6iOEGkkfMVaK60kU
QEdcmy3GogEvVtvZ9iookm4rlz5/2TjdvTF9yVY+Sb9ZaH1cL7VWnuJw2cI0GhzkhHP9D4g/L1Vd
xvRgZQFbMcVVcMTjFPx7We1yJhELT9tEvbEoljEfJ5uHdA9hhtWVdovB+2XsOucy3SN7hW1PEk1U
tBPYj8Z5Jj/oQJg3+sLVK8w8gvADapYIHQVATA/yYuvdmhtDhjdsEVDbHFSdMRzwci2M3p3E4q0P
SB6dEXOS8EcGhTYvPE/LAleCUOHhQ0WvYM4Uxw1jItQed4kqB5UCssInV3r2bljKinBxcYrNq8wE
Fh5UygK2wqgQfIMYPkm7C07dLfxwvC9dds0cwtl0lKqAlemaZHTSICMtAyF/FcvMcOSN1ufTDhhg
hgMd5Bcnw4Z/geYVrIQQpoxsN94q7Pv5QpcRKFDrZn/y7PJf5qYya3wAQe4ssRr0EUmvKSepZR4A
w5NaS5tLGXRYLYnIsnxR8Xz9GOJvM2SKHCYu9T4HrepsQoBQ7KmErSuHtGZxpZwHs/bIRwnKSbNi
/7UTPdZDFd6iiUGrIL4gin5nRstNkUMcyzDdpXYzgB4M+obl4GhyBvjI58R33GvMVJht4+QFDKs1
lQcAh4skyM1RyeQJcAmmY3Yn052AowHFMfG9HcEtWcGxsEl/QtuZNcJA76UCscV6yDINmvbunhL1
Sg081HGxiVh6s7tfX4KqmL3VMZZsuu+hhZbPUQ+Lxk3tTe+3+w/FL4pJT3INvqsKx4hoGqKwNyHI
pSTsGJXzh+vqSW6zMwDtCcrUxsMyXRQ/et9LdULmxuH6tRvoVa22vy3+JLvk0QI5qTHAgGx61I0V
cBuC4Ezn6ZVqHhvmSctkzQCfWFb/3DmUpsdexT6Wyc5fG7tcMCGQ2su8YUI/nvvQvMVyhJYc0hhT
KASbS1jSGYtoKaShWmsAnlZbhj+CzFVJFO6aS15anAbV+HJjJYRbU2ZkZ0E3/duxHXwag7pG6BUc
GoqGVtrn9uBJbrWwroBq2Sl0Tlc1/e5r/hvrs0+tUnT8VYSIQBC6fLv4UQnfRKtszD9tz2z+RQwR
/Lys5Dgf4HwORkBN3fGn41cBBBBsQ3BP0EVrjD/IHoVq27lVonuxxgafLeD+b0T5aJAu1nF8vHqF
wfg53mO+RH1qGCMzSzuf4Uv1fhQTPDJ72vkS8jMDziZ+J8W/oH6VhI2Addi4y07bP2HggbUpnRkA
UHxZiTK7uMMgERzH2CQCd+KPKkx/pNEp4xd3rdDnNtPm0eRmPQ6vQzSnBxm10i2w03LTUPoMN/8t
KaBH3oX8AgiGN3ib7Y6efCjQ59dXbeBNCaNW1ewVx95ZCfT6xn2SpOH4C/smEKeYvkrQ/NXOegAf
wyP/Y7S34HVVEc7q3NA9569b0lVKVd8AvDAAIDHwWp+695pH80hGwDp+mbK3kbaM40f2h27csIvP
XfURBMSCyr6DFDag/Lh+N4Bf/6y0GvfyAmj7OqrkgmUEsIiaXlUFrKdLHNMzGA9IpWUwfqN3AdBX
BNBqifbc0fSRFb8tX2oTR3Thi429fjaJGH1zWT3484T55cSPDLTs16fY+doWJEegLBdFlkDqVoO+
jyINlIWFt+7iE7Y5qPfwz5ClVBlLVZ1DQ8JX+bIk8TQEjYRVcUtRBqrwmorn5nmHqm2kF1EdB0v5
sOzQCXYwZ9kufbMWZGnevaHlG/6HVg9KWV+YL6FqY3UukXHXt6OcGSRqtEiizCmjPL4PDQYsZCwY
yo6OKfTiVU/mqG5E9RyWQEyy2749u3lwuJkFVC6YP0l5f2cqAUNraXdJad2piyKudv1MQlgPo1sl
b1IV43I4fZtM5GChVi9LSHD15GlY+EJex8Zpgw7wdlBKsUS9dEJMhAhZEemMniCcZYsq2cctKZeZ
tVNIgnRF1XtxN6lf5CE5y8QPIRCOf6TVwq6BH/FDSbc27jrXR44ZFX+Gy4r0V3GF4DTeNKk6NZwk
4tRPyPjwb6c7swvqkvXH0ogExK1FLi6brmVChwKdAoY+8+ExR1+zNhRkulNFps4UW5pxRweXXb3v
pPZP0SfVSHTfkaQm7kSFf8HQeHfEeCXu6gSwwq5aCqgDPRQqq67RFvnFeazriUe14JtjLqbYz+Yt
AoVKN2taLJE57E2HykfxTyynCMD+ZGNSEavyvH2m4/JU7v2m43927poGvWBRdzrY/xUhMGckGEGz
YW1S5SoiTuJvINGNU0zWRQQCti4/tSow9vjeEBiZp4oIST0KMlZuhvAcYwVCvf7Qychm3rYz7Lyr
ODconJbj3Z3UVQGCZtLt0FVZKBQ9y1yRVM8S5tS4jANKil4aovGChk8kFwCHqLraBO1ho0CyOYIy
oA3L53xihiTKAHtDU8CrRGi97gWQkF0rEpYgaCrFTx510FZONIhKD9a46+RGvcOjMVu5AXxLLjhX
LTKxTrWsebRO2b7Jb6DsmkF9uGjjJdGeSBc+zOx/I/5lmmpCllYNnA0xjkiDwuVHktvC4+1zLwR9
paU2aiGf4fCrx7zWz1qX5KSbPNiqbjuMdoe5mP3rlKkMqeTzWOl98qtd4uSkMBPUP5+G5SO+SHqA
L0oKTOdOequq/ntcnsM2lmu9wnpcq3CfUt1LH6D4Vi7zklnORZI92TydXXiPCCYD/LkknPF1UhSR
59FCXyCaOgm5DuRSm6CaxXrxcKeiEkWnFW4AFEhdgMDGM33R/MbTjXBhOjwxD2Qb3GzOW8po9pEi
LrNDmW1ltHdSczoy1uY1l94ln1+yDKSxxc8TZyHvmKhfCo7TpftMpzQf8C+CEhKVi1RXdAtE+PFH
kh2IsfzC2aV7ITo2WM1Oek8xLPh/H7Zn6wDDDSNDB+uMs8fKKC9OXdRqE/hnj2nzxXljZwLu+dSK
zaaN6cyCM0NsW2ZfkE7+CQZetAXOTNBHOI5/nCVN3T5/Cwbqy0sT6+OVTz0nmfqi/g3VecE+f4YK
w3mAe6zi9BFsGkCDY5/x0sFPFl10DiUfrO4fzEqTbFca34jKypmBwQeAA8b/o5hIwJVjMmrI04r/
nGpKmypf+slYAws8Ovff5CQGyiNjuk5/oAYOQAJXSIvLJkGIgERwN2+gBVIh8dxvq94ATdQICqEh
CDEXccvg/vHNCx/t/f9xsqQugWfiz+wtTjsdIkoxtk5LuMtMjXBAvSdwO+RWhGPI8fTEMsnbCxPH
5UGH0ji5SgtNB30befPH9gDA3Iw7hWEaaGSjgyyp1ZNtIaIrqdYZh58eLWKAkZAZAaKMut0hTewL
I5JKRNBCeAejo8M2Qf2TKSewxmC9VpYowgFXVQr24RC0cZxAYi9rBTZaZgd9/qI0Ju4e1Ipv+VEq
W1zattS0E6UJ/uiC5QXm32dYy8rW6lMzhG0QEzBfi+HypVqTnUFj3V1NfKlDPDyTYNLkYJNJ9Y++
ZpGuA+hCc53nYXh08JQ7Ui74z5bQHOHD2iCbBu656gLqtm2/zTfeO8BEqos0Uup+x88XvM4OKTSC
h9QigfE2vnhgxvaBm+Ue1j2gm/t36846/F1zlBF8FxQmgcEvwkX/3Ok17oDfIzi0GDaZXvNn9Nq/
HE452JcKw4WH3QGxWoQnKxvlErp85dD6dAXks+9O9xUQjaof9Dvj1YSupJO43R4xcEvbdUn3TuoK
EdcL5yBLTp2hSKpbtd2v5KeyrJfyNHmKfZvn1AOfOCc3nWi81Xrezk0/B4LL/rSbtVWpZmIoHojd
FnzTbdxQa9lgAsJo2ggi4YtD5gaW31TufZ/El3Bc7V5Q7I469Vzamq/Y6ps+3xkGBtUkjo0XdBrc
hF5wXySoFkdZ9SBfmi0s8/JLTXDv9R1oKXH6Hj5RUcPO3ZJs+ju3lpNnXMM3ZpWHgrgVHcjHdwBv
OXXqU11l2KwUXLDUwHSo13sFjCtXwexfWt/cu9Btf//F/Z5BcyEJ7hXL1klIUGW+29rTWiByrjJw
UZTgJCSNxZq+k66C7tpu1fQnI3ODuxRN6kekIsXOZV4mpnjT36h7tTD/NwOrbhK/uLv44OASYKKp
AMurpeLN8p/bawieWCTJPmLub9IjiBaXXdDmdcacVSv9kM1WVRUv0Xv69FqErJ2fjj8NJZDnG4ei
ZbUTC1q3HYdPLgp8Z/BsJAR745FJOBR9nGv+Vi/fYtVdpaqh5aayxbk8soso7FwT4ih41N4ClGwm
fFBAAXEzPBq8fYGGklgYrLb27m7UcDZkW/wEnEZzO4cVPajMHdClTEX5CTfyUsBGYMv7ttqWI+NU
A8L8MHkyjAe0BhsrAgqePg1UwxwTHRwv4wCGyLd4meizXwwfwZFrNV5SsgoaILf0YjSDgADhStjQ
GerH6tT7w57WQKNOwhQ4ZCPPSU9w7eGRMEIc4K5bZ5yVXoCowlRgK556yXQR6UDal/HEpbhUnhBt
aUlJrKRqXJEyEEgfh6QVF5egLRZCpY4qorVl6ky1kyuQ2Dq1zMJzHbfybUXOY23kTkQmQSL8YBDs
xe5Gud2Sr8Y3xeb+tLt/21vJB4vanUKzVnFQpbPti6RpCkNWU/dg8L+t+hNfkENfaTEGJA9myroT
IXP2hUOnEWNfOCgzQbZDfMdULymxBnnnwEc5Vv+3Vtz/ttqp42kkT4vi6Kqdv1c8/53D//npslB7
ol34TedutusNyldfcxPmvuvUw6WfKgqTB4GSaacr4M3ghcf4Wy/SymdugsVtjgsxKtB8loIuej6r
4oHE+NazzImaEnOuDIatWyBxxEXkNf0wE1i1lBJBCUIbQ5+4ucm9nJmsKCULzfPrJ+TFqHnU5rPe
qzJgo0p/iaWs3PiP3GuYe9eUa4/Jdg7vQXz7yGW0aA6vFaP8HGk/9tlIWsFUSYc1hxG/UkESLT+A
W6YAbIK7wEjCmHfu7TViNQR/DCp73rdeJmHUBU6+NRXOP+qyaIvJ2srSnFbGgv7YQJ52pCj9DbW3
wE6wg38fvZGWrEw67oghIasZmp3ud+GtB8o5AVd8VoHDFqbhPIb9GVxOcNlt4TYerKYF1YvQPVrG
INjwdtoaprSUJuAYW+ZQxCUZJ1HYq2YMJwLLzef7BWWSbeavWWWB+PVezYlQ8n7SJHU6FkxEeWE/
tnBCENISQDhcFIldX7ZhAxJH0RbABQrxaHmbtpQL+KpaZgTeRMFo6//TPbY4bCUsm178625wTzty
uhIrjPeKwh+gGugKy/Vx6fuaxL+vzZUBWtuL7LW5LPK7Ia8Sb9/jfO/8vbu4uHnwC/stOvImKiwg
+Ob7LoxtpoVvomKho2Auj9Mhwa8Y/rbqm+aegpp2hM4fFZL13OOJH5CYgLltSXMilTmaOLrI5pwu
2WzvDhSSmybCyTb7Ful54YZZ+WAOY/3ZK1TF54BhZnKiBbPuTx4qK3lrdKbGDJ/m9iTba99Z30ph
RkXMfK54QV/j+fUSuwiqcNs00l8+8L+AHWdha+/jeUP8NtogGWGTgOp9ws/yTYotdEpW3XxqWRr7
TwClftylTr2f4gWCYc9VmvLLeDbtTXfd+qI1Y/U4wGjrrmZKyxC5zESZdnwOZCvkiQ6DwqWFWqiJ
slGctKjIIk0wtetBu38kiz7mNeb9PbHxw5cP23VPn54jrTmelivceDul6TKmZ8vziXgXDqOG2m3H
qEadxTzM6yjSxEo2evkMXUIgoDWqKNaQvV0E059C80DjeZsQVfeWDi7kjhGaJvJEiwxaEPfXRjLb
L6kFvXDX5HZmtjyTu4+6zsQD1Ln0GNDJ3dBZSZxhWHneUMj4zkFHRLGvi3xC4mjP41c2CQDQmGjP
r5tn4ZYdVM4Ep2q5bIRqYyUjfdO01DBn3E2TODPAHyVk5o1adsOYzBABlVhBdx6gFHQmU685QhDr
YwEx2pBPr3EOXe7aWMQKITAMkIl6uS7dj2PObJWcaIlvaBDVoFmSpyERnqEU4eo+wgN8KT23fpjC
xIeIMJ7PP5UHWF/0ZpnOL9170V3mIrZgaV9OxYC62u9V+9kboMasjXAqdEp8bEshQF9RboHsQGGD
fxc8/Jr+GtKU5rFHkJhsW7afzORm1eozBRxXEpYEYPBX52dKrhf9VZgwy+t8roWzRoerHYG4lKHJ
A/8cHmXUWgMmjnhxCF4eBZMxFN7H/5wbiL0yaLtcp5FXy0iIj44DVkfj+vucG9bZe1ZtwzLiXckv
a8t7WzR6P0VrFBDKquzqpFOXMEIYWDrxMVyeZerG4oC8/wzx81cuV/KKtGZZDQzTxdjLtyvUQKgd
XCx+xO552WspWjUdOtCq3zDPs57ecGI68dvoGpOOJa24B02yQuayT0yggX1tAPfU0jvTaRLLAKYO
hJAOc1zLyy+5kQE6jm62Hl+lUma05Nalbj1dGXpCeKkDAlrNt7uHc8rm9+uNHgTUCotuS4CTgBEC
QlF3jsZb9DYO8y+MzOpY12rm0iIUwf8IFQdmJQNrleB2wrwzCjkmd8KVzG6C0OR1ZcN9S5MBU/o1
h4mRhG1JeTC021II1BtxwkOi+AHT4KoaQTqFDGCOKgxV8nn1bJkk+RJ3RZ3rEEBnnRtd4qQVoVSy
BGhPT+xDNaPTevZhT4II0Zl6mELsGCYrKyZYPgb2CDrV+YJZ54eeXYog2WuFIb0xMRBL5FliCtbB
rJ56zsrnwUqn1Hhrtm6FY+h1R8epYsElxnOM8ykzO0q6JNTIr3HC0OPN7810WMZl33MvQ1mGAOj0
F/ymaCZmteb5duzpLywKbLX54U6W2ZvTOEk3XMg8ju+oVIDHUABCEdP0PSS2OLYEoA9d0HTK1LhP
LLm3CzWPol7oA2laACClRYoVpsoSapydjqn7UtJQkYQoHFB3VBLFJbrGaP8XwK+9MEwKjySf/WjG
TVjaJEQkR6l1U+jxJTQ2/OBPkDqrnMpjx9tG+I24LIbKxSdrqBD5jDf1EEyS9pgmReaQmtP5b1lx
3MAKRMmvtanmrrU/Ot5WiG1Mnta1CjNzMzPbU/iFsgNkC0/MgT30LMkqWnIolDNimEsJpm8EXY4E
jKqtXM7GfiDfhslTCkb79wLRiUWuHTpbVq89ohufSk76/ETYcxJEIsVVJJFEQZ+2ZG+rnhC1OZUk
TRSRTeuXWT+KmmDcpCECZJKddYTj3N4OW8vmNwrrgKHy5JzJvdHfsYdvGLp0u6KLOBSKc1nRc88E
ckPCkDoOwf9H9Q9O6nfCgF17d0mE+VmgPQnJ1qsu/0/Bw6mGk5TNrDqhxO/TZLxkiuwHqtfmJLG2
C5LuraLsWsN81ZfrwU7/OU+oWUvSI/obJVZL55XgGe8QHfIrRO50ZyWLW3eui8n0sooAbBQuk/EH
3Sx7VAorG0DxJpF2dBHna9y7yEdBeuysCFUH1uoKHAbeCRu8N4loVy5BnxVrGwW0cFzaRxJ/WZA6
qJIrFU2ki6NyvuJ52uSawqfvqf8WFFnNWLvhC0CkYn8GZgv/0Eh2YQ/uozJ5EgQOKkT/UQPvynh8
sarfUnXDAg810SwdnuxUld0Ea+wo2KWHO5AYcgGYEN4WSSFV7wHmFbcv7oVwyIDLXFMtRUs7GJVz
A8dLmPZ/868L2EZKc20aT1OUPJ8MjrVln0mt2osNhTweE/DyhF2JG5BezTToOBkKCg1v6xTFVQ7l
a8awM07WzPu6bji4xtRlnSnQQ0A6A/JlkLUo3sNgPlRQHuStg4IgHr9nDLlqFQtZaukIg83CDxcl
KnfJsqJymA1bsTv5QevtSpBGmR7M4KCAsbPg8yeCQledW4iG3C41At8m9t23YS8HC2nuKAjR8TpL
nuQ2xJcNy2bH7/7vqyAFYLRzav9ZshztQ8aOWGZwfwdr7c97dvvNkIncm37+nzS5++93BddFIujP
ywaQB1iwbcmzCb+KFy3hTP9JiqT5xLbYkOiFAiAR79lx+uUCww5ED4ISGpEQJ05XyKVm5swrlwKA
3eUuN8uc/6nXezCkgZs5yfMFo6zmxOCWES64tbhpmOTV14wRvXGS/y0cbeTiIG88j943I6ExBwV8
7dD/uRPZ6XIhdvD8WvdDvDIb4m3WyiivmxN+qUnoWJGkaY4GbTe/X3Lvgd5ZB3GKTiY31K350Ny8
vs1pJqAJZua96DSJCT4S6O6UOjmVs/1/egHUGBKwlEWPsPoSZHqKpoNLRxZy327JkE8D7AN04HwB
dzRV/LzXf/7lKNaPnZYULgx13ilJIcS5IdJ++WJjjZmsx4fn/z8lSmG2u8lE+fgzaMch8S0gnc2O
MJkVZMSZ15yDBzlqBVMDT139htNhxQ+kSD8Hy6iStMpr3OrYbDTMpWfTww08kwGS7KMbfM4/R4FA
RC47tnSlvmRm2gBSkiCnjwyFPryalEj6XANzfX0VuAmnGxu6WOZmE5cdhbhpF1Hz+0yHX9/KZL2n
NYpHA7QpPGVMkr5wKqg6iYVNpAsOKBk9+IrGknxLZlE2ud2qndniQr6JBY0c+emXVrRPXEXoIm20
cXSHAWzJm0LwKm1qZkwLGNFLH5JcErFyYvEqLC5W5wr+iiaNQOnLvCVbgyGSUIn0BfUAN1seqKn4
bSKRsMJ5y9L9mEv9ZwkxpF3O9MuH20C6CIWp7dVMcZnK1A5iw9ExvCZ7U2VyR4Cz2M1aW8yL12Cr
1MZ2hkJR7uf1wqSjl74oKCrYXEvZCm0BBNHiLpsYRdpG1ZnuuIxkl0m5+w/wQlml0QRWQMo//5pD
yFuCw7tSWHKjJXeyZmBqlxNO6KS/qyp7iyxuFvnMC2UhBxMbmAo0DMPF/iBnId//RfVjPmJ2EurZ
NBc8UjHZk7lCXO7fViEVDShXR1u//h5kh1S0VttAltTIp+23QO+kTau/uVSgoyVo+cyUAThbDYzp
2vKCifW2uKiV3834/Ph+Ne2iS0DnpNgYTNUXtY7gCbtpl6TVGFR1EUmTbilj8xbebq4CGeq7/Ei/
ySFF2yHvnlT3q3xVlLfxPSDxEmOba3S3ZK9SolSzrItdEAnWmXJRaMVlke9rBaH6TsBIA7Grly+n
KcXO00ZmOqUCmqNdVims0rNDGhF/5ldZXH1bi9TeWtaQRbh0zLWnWn58SIXuwAzVCjffIGLcws3K
l2Mst6oZHOHN/Me9UKDB1CWJV55x6pe2E7fqikvEMjpY1PXS7CLlbvNMiObVfNeITdgE04BA31Rp
DGJinDjDUduE9PdyE0RCAPk4TT1puR8ZTY9+AgNk7tot6nYjB8tqMQLh6JpmMow17aBm4usNArhx
rWP0JjDSGLpZtwky5WQIOVmTY+BijZRW0d5NuId9drbCTi386M+o21d+MsqHX2nIGWBviubTbuNf
xij+W6IFIVj9xoXUXOteyNF0vG6caBkRz7qjuiCkzoKvY93TRKd5blQ8PPvyKPwyzI+YBBwHzpwa
ZKCtl7rljHKluol+k+XihBvL8wA1SavP9LXcEmhdeqJfhhE8Ob2ZZ7PxUN5811/rnxbVnuu2Fhwj
XJjUE6LKTZe7TMSKChjbp080RKjAZqw2t0IWHw2tvovMWF7IxC0mcabgQfhaEb9lXw2jVo53w65O
6vuO3oklmyPrG2dMdao3PQiEPrWLmXDA19cyiPdl6Bhe39ffHtM+5NDKgXrpHOu7n7ewMIX4Kqdi
LAlAVxSbTXPfqP65KMeg0smy6nIxyEu0In0Zv26UxXcVC34CA+57OUIzuum6629lFmn48qR3JGAj
7L8X0j2x0Y9ThEJaxnAQ8SLIJSR+QETWcKhTKEMyVp19B1tro04Z8LgU9r+GSJqqhVCyWgiDH8fb
lSaBoxsLjBv6hf6hlDvKz12QkLN1mxsa+PFBOv/7d+ACBu/TAwMHt+PwdwXq6vJYA+GM3g33P2Gb
FTCeP9gsqtP5wuBE4WCWreLicTFTh9i+hOR56ctrBnVYgE7PayPCTdyMlN/wrlUEYrtd3Zxb0kIf
m9FMqtzVRcRdHLJLpIEJxirdoPGh+Se4VzX4deTefaHHs8r8Ore4QQ8BB1bfcLgNspw8Jv2cXJSB
1SK/cVL8jWlVjACU4Yu8DCqm+QNWvA7V3o0Qt905HYHm6ZxzsymjNaaHGxf4yW9kjtGe0m9056DI
qd79yZ8IXwvS2jXk90UdRmSu8ZCR86WojYTfOuW9PEnSzYbB1v7GmUIfiZhgOIYWctKIz4KGy/Ww
swq2b3ZU+Tp7x7H+DkytTGK2f8J3hp1H4AmnzPcckOnIVE0hLMsk+O0LyImhm3j+JQBqegEyLka3
0g+FqibDzMz5YjeO/sdLB5+L3j1UHCYOBNOJ5yzPcUI0KbZ46hOsh6UdJvxIS8Sbk+qyycg9Kh12
Efbf1rnwklT+TNGs8BzVL1VOtcJziXh/151ONj80PFXuqhzDBdQhBaiH7Jd+2Zq9mzImfajDWf3c
4OhwbAEeNQT5gw1rNhN1ab9E0kDv8WX/w5bgkmMq0ZJcIZ6f7PHaPGK0gLvU+/qUldeiafRtjTYq
YNLR8FZUiFa+oaCuNQ+k2BPXKeQ41lXS10xI4gUT5Lpamlcit8BwHrip2mLbZHO1PkP8ia35qdKG
b0swFPB1U14orjVQYwRue8Ih0tab/hijqrmPPgLgQf+EX+4b56RrPFGGmWYbekFLGkved1ZqfOEV
X4dMYyTBWZImWoTQTgUxCdedC2IUnvOCQamZJiwGNeLpFtiQ0Uq5b++766F7Xg2RweotXcON/vB5
KsxJ1EAkaXrl8HZixhCEY74+43gbNB15r/Dvzcs4x/mtJyKVf0ek03WuN2rOW6Z7AkHrqPWRAlvo
DED1IxPEM0w2gbG6IFnoaVUhz8PF0Upa5KTCQ3U+ql98UA/2Dl+cMIMaK7e6jLCvDd5pgMUwOy7Q
tDANHCwpuIbMzDrbXKMYBi9tryGnzReEYjeVW92qSMNsOT3txATrrphcHtmqk4bA/rUy4Ja8XVS5
nButMJDiO94qiYBM46nT39Tx4QYYloGTg4w4lYUDr07C7kpqAZTnhkWy28xxe45I1RlYCmcBi9Y9
Ue48RqU+RYVU8xV0KSf8lhXB1Xqn1tKx5Ju3h651RnXQ1O5BjOZ314menl97J5OmS57ciitpQ7XW
jzZX3B27FVjYtCT2F/Psd5AZWmmlHBF/e5tvl40cvY9nm3ppJ+Fo5FtosfDA1kPVTfDjqilOIylg
NVX9fRL47Paqn6kZmTrVb2234TVo1bqiEFEzkUmR93X7V0gCS4KpancIRklknhXPNBBXirz1yOuo
LbrkM7aAeJEUsQGZJpn6ElKktG5SZj51DOBePXg+KlDaxEHPcK41gZtKs+2eV9tkQUKjuru/+wj+
Hpi4bPZqmaX9lFlEJM2/k0zFO4bVQGBIlFlcVthro9RwAhSfM7kNaV8oUl3PxcHg13ChsfUOwpPp
Uq0K5/mZB85oXtgGEXuXJyaAJBdj60itsipGDSqInoZrNIDw6SLpsYZj+sdJEcEluSoLw+1Mf4X1
ju6JgKeaQtBuYbObKVuSlD9+rmD3N1FI4P/FiidKeGKyCgBJHlEB1sbKU7PThu7oZwcK80T2Zpa5
G6ydf504PdcuBm6lWKJkoL7VcPMyKepzYVsm8dqXGL5y6EcqFfIc+a8+R/w9I8WU7tZ5itsIb+1L
TO6+rnuMdEhOFivK/ZxDI7jhFD1AS7IK89UVZ4JtroWX3Be5vYJ4O6I+cVFJr/5EUV7+3bQ3oQwR
CXVGr+qD4YygxLtj/++A5Wazi3qiiEPkxKAUuei6p30oDJrAFupo8EJRptYWPl/CirZFK2gtB2rs
zNjDuPCrunp6g54JjWRIR2Xgge24FGQiJhQoMxrtSfHlmnqdJAdxH50vBtuF5TGBhc1DEexlD94g
StnH7iB9D3hFEMwAaqyS4JU1XvuRPSxIc/eJmVatTRaErnN5/skmG5Ekq00YId1gBBVhHTZ7t48J
cjYg+fxAuj/UP/H1Nd35/kHjajsVvFw5V975byfSWC22/FDNYXmNPc27ifQ5wc+Ugth1fitu6brn
1BqlbHyLxWlHzeYYLEp3yNS60nC3MOZRlQFgQBzza55BLgqbKIBAIG4lLAiraAg4aitlJ86RO2TF
kc6+VM/zgsjMJyweQVc4rn0fItjbAzoF6SqAcUnRNNnyJ79enz4zesCr10Jk8q9Bzj7JLhHZT9pJ
POAddw7RCn35tN1IPRIQ8GpXk6QgSML+Snkd3V+NqSiCMz17743mBwgmjOhYO4PFVdQuP/OJndkv
6WGjsEXq9IJ9a5znXjWKtMXUgDXHOlQDef8uTXKtWVW+ElqQw016QmA6O80ucY2iNr7tFLge7J+D
wUU9Yhs5LlzMs9sPPjDg4vYMzPeH19AmBV8J3f/bO/E7c1C05rGBu9utQLHZS4v/p6SDqSBRJKLi
0O2aFH3ugh+3jiMLMSZF8NDFbssM6Lr2MjbQ94kzE8ccD+3v5Vsr1FdeMRK9cjG2OBy5cs/Hm12N
StwqBlo9vsrQm1lXI07gZR/MDG1r3tePJR75x41m6oVtCa+0WdqkfLejrTaiJAYGYl91MJ94CkOY
ERqtDmwJ8Sa+/rfUDcA7zumNloQ7AdTwT7eopJpUcovLZK0HhYrQtDFq1v/a8r9kqy7jCWIGQiOs
8jZIhNH8mrfK1xL2M9SoRNzaBIUHMi5OajpqElg0NVjalGFUvnIkww+x7xMDB8Mr/hhv5fj+YdBZ
VfQX83DwsbnB9vuTy71kcO9XZGXZU69L1qfbzqug0QOh+yKrRI+RrO8ZbJNNB2tBo2bYEBbbUYaO
6kKeYx4k3ROoZkOZwqkjziEStv/JSFnVaXl9xSJezSDXIqk/uHgltR2Zz3tMsS73aotHXsi+7oxT
EgqPDDAj9/i8Act/+8h1VyQ2W+LXRtRXrW6NyJzbw3zcVjY+58k4YrSyuuJ7TlxZatXXfY5xf/U2
nQjFD05k5BazTjvYAXIsfwrP6FjtbJwZ08oBOR65Vif2mIhTer0GzeRfrvqM5aWfQu/8O4mHAU5k
HNrjBUgDCq5kD9jpZmqRHP82hTNiWwJGSGf4F2Zu1ohxMslBZyCqwXmbUJMuMDbHRNnmNpu6MK1u
oXg8lGF8ZzrR+2XdZIxltJqwF+e6qBe3C2L0sQcl+wL6U1pSJRU0z3n+9zTjte+4RLuenp0Ks8jX
wfFNSBiGVGcDy0H0sfSLGmpv9YAqoMgfUYEjiyAPLBmB9vtYj+hntW3hpDG0EDQ425CkbKk4VRcR
+QXTjLgLdaqeDlF125v7FKkwIradPOOpIc5LZX5iH7FfEIE5YFZxXwCLFG+zNQjFg27kuDWE7BPL
boKneDxyYn/grzFFuV/Z2NdoRDuC1VW2+i8lEU9jjn8+tL2Etcnr/AbrXfi4rVjXZXV6jZX4kRg4
60QR5dn3oTK71WeNZvrBcUnwMGHEakj2mtfRBZ4HSbLsHTbHq4Xz4j45RMRlaYS9RNLuBgdTVZbo
pIz6EA+1EUAksTnwsF8I/sdFEQ2oUk5wp5fLABIF6FApb8tIxFP2afT07sjPRxdH7zUZvLKgBCji
acpoQ29XzdKFN0kgt1VbF1GZgymkGAv9Cy7uvIGAQIeVsCk9u9uU+Ro5nWml2J6uhsb7xq5k0zqZ
F/cqTinGCpYbPJtpMWbiqGPqmM9CfFlGDN4UfPAnDoxabS6BG7NknFH4N9E8IDRpyw2vd77NDlpa
pAOUSctxGw8MyP67Rb1ALSxT45Q5xmv0zy6lMC6ZC3eBbswU6+BZ7Vh/dEzC42seESKlf4uguq6g
8wBFwDoj4Vn4iqj1pAYe0+dUxIoz5vVOr/jLpNxQ4sMQahZA6jKyk0mM3SGwXxMRnEkpIHU82pU6
pk88dg78CajHjdtbV4o6TrgWimlpfj4ib1Uy2XxwJ0qwsl05aAuZeF/tX2GugIeDyKiVahuQXivb
3NTe60Wy3l5vOS2Lsjt0lyXNtc73RnbRk/hshfrj9sr6gVjqXM9cbqnPXarGE1Ge2wWsH42g5PQ6
wdMEC7/4X3yworAQiIfkCFiOrjyv70yh+IDm1RwwiW7QGKmI2nByAGatHkV1ZT2JEVK0FPC+E0mN
A3qKJW+rFFnXZvI+jeQiP8/tmmse8aFX68HsowJ6gtuhClGd2M5QglgwawJ4LkRlBuTw2YrJqPDg
rffb875R0qZHt+06dQ049uOb0A3Sn0+AkL05S8OYP365Ei8O8+rQTkN1fwa0gDoqhe7WV6oVIPWw
/mfr+2+toloItSm9yrfh/1VGgSJftXIiOUqUO/CulwKdXY8/260R/iBB610XVDyEcU26wrIjnlmF
zmBD7xKX176hFC34OqTd+RTFbgIHGjGfHfJQs1TTt7OcUZGjXFoS1cRLmF5sQIMNxvCoi/xEuNRm
0qrgsgN93xGihf357ggd82eh4wxn9VS0DnWWrvhAeb7lxSUsXt9wrnu39kNrFvfoAaNaKB7q5EW9
fTxFzBxVR2i1o+o9knzuWUMnoT4icBnGR/M0v8BEhUc7qkmUclcjeVKp8K1goauJCDOA+ta4SKi+
90QIWpx1BI9p4oxA3STNOnmehiEhaZCFLo97LL9UFgqua8t1l6tXV4NT3ddQ3mMf0I62LaM79ogL
qBfSlRLv7AtrKlEuX/L2XDUIRUVJLEHEyybLTGuUbuptMtBwquLmJ+3qAbvMegajMTFY8mzfMXfs
t2nXG3smfY9Vj4llda4AGiYvb/mb02l7kgc67ou3zYG8TZn3B86V1fgfp7V5nKQ07uSaeXzzL/V7
dwIVIf7bHLSfsrwFAQjzCMVhwYqk3WGHO14HnBtjRyhB1/Hoe7nqQUyT43EPnVgG5QLnCCRQLMxX
nZvmJ/lr2OLLkDFUOort9On1wNzRL/hZEmagFhG8dFKcprDJ4B4an/e+13isH9mMlw02auO/GdiP
mCqIA2H/+S80HE4wcE9yGfUo+OjI6yJvBBk/m3cWJYt/J2dA2epkDpOOlq97JZjnJBUn0l+vsGp0
Lt27yia/eL837omEobB/geKGs8IOjs9zDjFtyXFfAbF+Kqk0OrZ3MUluxLiQe3Tgw16aba1jF2Pc
skToI8O+4NZCKEqArFd6rjXxgf70fwqhROdkN4ES1/FjdPx78OCg5a5pHSXat1asMKMewEBvMfXv
vpS2gsapHVhN+0CWUKx2RBuxC/xE3ZrO0moVNwMVkAFDAJlPqV/4+WxOlYmsqJ/p9u/QrAkGSfxW
nJeZo6poB3SYUNmq+rPPu5cOpcHVJFRtuGhEomZEj4dW+K5ojHfF6nK9OaUhmDarKPjTrc+UkkMQ
r17ye817GYoEgbWXnUHKW0rITOXpC5QQE/JRNv7Dq4oSK06vqw8zWR0SFJWdccE2vDQCWw/SZ0GL
pZexfp6OAJfveBSD55EvNHPTtAlDKTIlKJtWQ0RmkCNxc4fneGnkMP+7BWS6tgV4HTkjZsVFzY68
Fvmx68pzoO9ZSFx9KckcyVRLbc1AYga5/5lYknrZ7Up9lpp45vFpY7Y+yhKm6r161P1/WS0PKgSF
tnuzo+Ul4zt11IHFvd0o3SROOSNdn5V0Tog08Jb1icgFA8n4WkvSpo0xjGqvLItZ3AK4MV5pAG3w
setBKpVWmHhZlaDb+KKzgu/3ppoInzZxPTUB8upqy6rXl5b4UHMStECwX4bElMuIuYNaSOG8MWWc
8U+SWCu4sRoUL9jqqqEYZ8yCBDWUajiH7+yS5laNv55sImfODxhS3SCJ/OMTRaiLj06jOA7kZ2RB
BhwHFvZXcAFRRL1uxIkZgxq2L95uB9FgAX2FQ6fVWaOsSL82yvGEdeUgtm0mbtSFGfBjpCTA+jsc
Dr5E/nWbXhZwxGR52Auix/RH9bNoFhQ7HuaIVgKUFxHe0OKFrZT/519BBBGg2cRGXRuFJCgNP3gU
15Jk6eNDSKqGVWYRBB8mVDEyzoQiv2MJIiQj2IpWHLAWJ063w9q0efg6hysqcjg0zaRdTXXG/wCe
7DbGOyo+Ok8E3b8f6Gs6I+WUxasZkIQzHkyK3aBbpqSsf7Lh94wCQMsw5Yf5vp4udrLORp+hUhOb
K6YPXbu6tl2OF+jN+0QZVIzjNtXE61qjNpYugJ0P9/oRvps20BdwBEIgPLHaTLIw278ixBiEoSj8
xhHpOVLY4tQMCQO27ijM0Fa03kWI77JSiHkIKOBxpQcNfIoAr3ZkYzXiBjRxqlQ7hi1c60HV5jeL
bGW7pZEl05xcSNZT4WxziY5AW+v1AGRZqXaL+DPnc1PE6ooH4nxrhJTtgTW5xitgUyYV6LiFv2Pn
oL79VWciOWErNz482NoZBnyUnWkMBUIjycdhawuP+SXxulFin376uAwRuMg3tlcMwK14fixFX5tg
JpMaBubBjD7XvChTaeL3yEc6aTBb6rTfd2Jq+/2pooj9lOqsBBmE6IH4QnMAUC5vKCMmspcbQQd1
gkQ+30psPG+RaZX/etaC8gw2zw4hQQkDud/CY3qkpOwr4wXdM5pcjv13MaNfTLCxQX/eRdkWpe8+
vj8wqX+1KTkOlqFODaCd/FdwucEsmcWlO8Yxy3xcNt4Xa4h2ipHJ5xbj5rzIlQQ+8qwe7H5w/8st
hELQEt4jzXSM4/XnvGnfF3Zh1gCf1yKa5hSC+rkzYaS3gDXn6oOHVjp01I4IOn5dWAxMRuAc6+MM
FDYuHPSVmxWUufhwnOKXeSUAxoQQ6GaRB4U3zO8JC6Xh6a1J4sFnBrGBKw6YDTDpIg8HZwAme1nh
EJyuSW/8zRMCvjnwHfJm9WbAxKmjZgfWpXFYzHtWbtrL2SJTqNSvH8y2DP2iglDysR+1XIvt6Vth
OwPlOIJO153/PkwwV5aGWhRTBe4zGob4FEMQD2ENTTcvob5zt1k5GRIbIGDZJqlMIDyTBljldMMt
o8ghD1bHdPnVIxHLkeT+ZKRttugCk9Deux942/wneCPdZOoi/hCmCG7XCe2UbrJlsmkcFBGz2KNn
5xFukKcf/+jERQxNicUZFKN9lWIK7wwi8q+7IDnMY5aSBgaqAH72Gl7M6f/kNXfd+RdF8Gy/HY3P
VQPFYwa1rafCwHRfUuLyO6laKP89a13vo8QbAzIsSa5dCkTOK3kuKqos3X90UOKCbd/UemxB/m+R
KgBHuBhTMM08u0gHqimCTTX/Xmjoz0QjOcp4HXdvfUpnNJgf2/s0EbLG20bzFqOvrw9dxQ9Dylf6
F+53aJT+//S/xMjDEqt5zCh/crqJN1foMWJtK244bW2I8rbdP0k9/2Edt2GJJ+wwe6hqqFMw/Nsh
ZQWUnUHmj9Z4ygLINyP9M682nhHITMHCbCGnkJrhw1m8BxfjBTBaMqCSHbyYxhOks8ninf9Rp0aa
w/lT+sUoxHCcvAjXYJb+Sx8QATy7H1S3CVdPWa7U1ZzYm/baLZBmKSBz1EyKyROseL8b6/ton70K
YCVHjQAVobeK3CnFhNryVt5tIzTFRWfYuoFoN4nyEVwtkEadwXnR4GVE4TflZYAgnkfQj9M6/moX
089jzevfSWx9VCGa6ylR40OUxQBQjohbMF7gJOgSgGEXdq/yDISfsnKflNWBm+CgFO745G5lBJu+
llNDewJNgXojEboi5MnVNBYB/hDFkn06HKWFC6QfDFieqqSnLcU7G6ZdkRGO5S8zqAYS7fa7svKW
S8f+6VhE4OIAP2OrF0YbmSJ7c0169e2eutOcThGDNruG6+OU2573/fNz68SSoUcjFqQMHhEdjvUd
9NLu5Ij+6AW4wQBX4vqTXWZJr4FwCZnKNMywweBSfMdPW7USvZ2/6WZ6sqn8FCiR4pT232O6/Z3r
KT4F0Kmaq3tuXm2swgnqVKCfuVVzNvU4IJZWHM0zC5slBJ2xe3qTAknjjc5Boh/WIttI9yPAFxss
UbY2Ghd9mYixG/FUt6IOIEOJvkZnJQvvCrOY9QoNnsHv7S4QGZjBY1XAl5S4biPf9GVKLmfflyC+
hC4Lsg6nj0L7V9gIcWsFeKvUHnlEl3o2/y/Vy4TFwvA+jwx3zoNW1KT5VKxeJnG0h7SDt4aWIdsf
hrWWBQKrmRXMewa32FhYZo7+J2Qhh+5zbfd9qyAofiiadaSgV+DBMf9W6lMAyqGaK5xSXFx+ke9q
czl83x+pix+l1Q/AyaGdHTs894UxLGAvKRVxOZ7ZOOXn5zIDsZ1+pPa/u0x12I6DqpKp2SG1Qxt0
/6bGapoyUh7wCavPjm+NzjR+W0xBpVE3Z5b00T/ULbMF15+qalwcBC67ZjokLCg7WP1r1EDJYW/W
P4GzfQrRuVA+fpbp0ow5rz32OTxJNNun6uJE7lJiblFjYzO99sMnYxXJwjnwa3naVSqix/pfBWvh
/zN1gdjZ71PIVURKgQo4V8wptwczb2VcVW4fATDTScQeYcKUPc2BMw+BS0bEI0WcVuaUS+dJVO2v
I/s2q1vKV+6ZM9S24ndgbNaUuW0dHPn18NI1gTFZKNfZjwfffGG+WkEsq+V9UDksKeswA6j8lUyu
YbOiptr0vvYAMRVDubr2KW2zt0mACp71NZ7DigER5kbtCe1D3kQulm3MPGEJrQitFeNPaFHII3zL
KeOkPRMZAyuf6AhJTyPU8YRfRJQuEL/mLH+pnnuYCZVv0sQT/2i8jA2qpuDyHjPZazdWuKfoxScB
dXHBCjbjVJQnNmQ9Y1vLqTf1aikAHYBqhuNXZGSSegZGTOQGizqnYgbO5w0csup+cs+dQBalYeih
xrkTwZqnRwzwJ4wZ/IlULlgjMY2ijQBV3LqeLYnbZbc+Re6WDRMHOqzuGnWkSDml6THXa1ueg3ip
GfxImZDMa189q53q4gg4pVovHrJ6XaLLZqWYjJDrXyba89nE6epWAn9LJ0dHbBX4byZfna+eTzjw
Ibiwnv+JoX11oz5tfpGLcJ+kOA2hGwrfA/CJG4eByvSztcsUyANS4jI+G3hhUo2NZ1X+iM8R0QUe
1ZqOZjAJEWNx20ej/Qo7ULDB6lnoK92LZZ4SHvO9gflQjyeZcByuywNhQ7cqLHAoK6I7c3iYJkQR
SvzKF2jwRRVi8Ji1Ly0iMgyiKSrZE96cDLW+EPE59MGBtQ6CIPxeCQDGIkXlY3kAgBbeP3doaG/e
KYQSAE7AO83mNi2bB3Nq+9Clyik3I+DPXngTpDtDYODpEoddQgvw/LV+eEUeD992QvHnWR3tXKPA
bG6k6M3jXiSgmffFcbtlQtP1LoTmyKNvgBPzx2abqf6zWl+ozRnFylEk0M58m0i/hGvpDxuPY1B0
n8bK3UfoVaPi2Y4/ZjOG54Z65kuZqEvHz3tPTp6LMeW/aQFzoPXRB9wlZceHCjwD2HlcLJCGHez6
SqwGLk0sAmd5dQKnJSM4RztyOZdElqi1rgON0yqIFS8ruua1PjZk9RvqJ83CuruP549kSQsTWoGt
KQyvGrS27OpEJcXQTbx/7Jbxq70cEUabr7WZYyH8PdavX+Ps7fVhwzleAR+/mu5wp1yUWfAoBjBi
JG/xogDD1XgPt7AH4WTd6oo0B6uNNG3s2DJEOAsmzzoqux6eYGQvqIIHWkyZhWynxrlCmb8ieg1z
ivsKoVx+oxFdBYfVMw/yPTD/Is2xsTu0PRz6NigLZdZbzom2i389qjK0q/k7DcQsSj9p0JvLUxv/
dv1lQBTOTuLpGjt9A2scRexbP3fJxF43MPIJSCa2jdEPk4K2QgmL/ITWT3ctN2fwyOc1VjLsOMzx
EJG0DGYJuYEXzR9c+MMSdTHHXWqUXnrgHDpfW0vgxm8xR105RMiwOlDjvSepT/kYGDNhsEXzqdKt
CghbL8kZ95jgCx3lnzjq1G4sTKbAeQK5QxcqEf+UBnRssBdJaaaT9qaqKPJgHztg0wN5lWjL9ZNS
0NPYDEtJWxEOVCxiYB/zwl02Aw8TelP+eoPAu3tmZoIWYae7vUaLcbD9s6hnyT3HyF/rxxGR32od
DBLhcVGVCN0STeERA8/wLDr5kJgTdqFLOnlXS7dH327TjCBkfoqF89cnlQimIncBifwSwDhpf+JY
UVUrdOrxxyZnIC4COlYVrMNDFyeJBWQJvlx2bvqRsu2lKrk2vD3ShSrennjK9KD1NIs///MVmUjR
U9aSTqWHEIwrlUbAU7D7yeReSIbWp1xSjjoGTJVbg21q78XppyK/OmJwvCQ81QMEoO8ynm49+4sm
071Uz/MxE+jG2o4y5lfwpDquUMOL/i6b57XiJcOXstJrfkFsugNtIP9sKb+9bdgpWvQ++ISHLNLt
Fy3QuLNEPnqMILKe0c56HhnpVaSbYtizpm1POUETTLH//tOyGNbOlQnne6i6ld3qRcmVSeJ+05pf
uISqQRJgbOqVVTPfENow/E8wBfyLMLbuIyO6g71R3q/+QAhDxHkL1reDQD/cr1qr4cWDBdafqFAS
ONIr4PmP99lghfCyxItMN6hl6mBoOGOdVTDTQjonhQdjAPNNXJYasdLrGx5kM6BRhzzGC9XEL/j3
dxLP9EORXVFavq+Q8cCwZEj/kY+CS48f9Eyj5c9/Vc4NvZo65AsPMb85IaTgaj81KZhCsRAZeCkN
f5yMo2Rc8hKS6nlE+uvT6DtE7b7vee11Jz35yXAJ/bAckMmp70bMuBdW/uv9m9wENqtP6sa/cpd1
k/5VVo7zRigJYK76zDbuVEAkcEoZ4wCMZaizO/SKtzC57ENkJBGQ3BdzUtwB2N5m3fiAb7uyBpT4
GG2EsHrzqf80J3tnJZC9UaAzyN+UOMPTenZTpr4fHtyHkVxqywqwr5pMapaMUSUnEj2TJmXKkB4X
TpOCJe+9I3jnvhKi5kou/+YODxbBD4BpRJk0loyu9JXAkjrKtKkpbkuz5WspN8a038rva/cpPk6s
MD9fNBjJVYEgr0naalVZq6qhsky4+ZwQCep2yZ2wRERSHtobxEWf1I4fAR0wIjZCs2Ch3jQtQt4c
VlKfLIlRt6LCN65YazmAk6OcjMABJYywRbAOA0FcYpmvNnRUvAriPkRMKRkq7RtGfR5bjggckUdV
q2EDju6G8L2WnrEJpBDj+ZO7nE2wQN3h+tSHC579YBsWp9xn7jt4yVjEfIqlH5tQmjvG6xIAA/cD
yH8ktTVv5+45iG5umAzkf/Ar5qTZW86xKCVcewMhipPf5bopKq8v7FHsrcx0xUUw3U5AWPHdqyFN
SShdfNwUX0Ru9EsBUcq4KJE82NZZXzBmLrA7CBHC4plhsCjAMYpSOd4DBc6+/IjX2wEj+j/sdpMO
sQuMF0qpasEe+phzQ+KOyv2lZob4B3wwvbqzwKFOTp2A2SUi2MmK6UoKcgBP+L+HYbr47HResw9L
cfXEI6DTzDJ6RqykCPQXBOleS9upYpSgmWSMSWiPqRwysbzaCLGH2IrLGWLXoTTtV1rWPHtgzopX
N4j6lZ/T33o8JA/S45a+ElMJxn0V6pMSfkhIK++uJ+pgRClKtwrUAZHLxReWFXKaFC+fgDVAMCb/
03SEpYUWMW0nwxFxC0PtmatIqHRK8HXiGasBdBy2ipESuOxVbF8vYC4sz5s/WsouHDrAFewbsLWX
d2Ed3TH7BfbIFLIuJ2jj6qKOwc7o6P7FNXek23WQNJW5ezKjufmd53y078QKjlBAnnItZoOhJj4/
S1STVenNDJwhYpy1zCo3s1tm3DcTp4O32Dz4+4LrJYApJpn2y8psggWd36grFJhcvSOGsNoISBGk
Tb5zms0QH0Z/RelR4qs54lmOgWZKrHi0o/BSK6LSSb9A+i2vEsphkmzVhwNUyF8UpuK5DrAD5lPO
5zjWeA2jeW+I0wyOto654pi0/WOI2iVuzypuBNV5zqWe8W5h7KVvA+6+F0YTc8b0rQfMvqCAwB8e
q4bmotIS7xwELAI23/J0WbFosnIr08Guwg3+E2MYezMncLEuorpT6RGLEzFScAaU/aJ8RdDx0RGD
gFLZYOOau/PEUR+GP3K49qf4rkjPxgffznEi/Wt+07ml8FV0n5oGICxVkh1tPesO6JkDHvroIm0P
Ec3sfCZI3mtr8BIdT8yHGWCuawi1O3hEA5fguTZyxpshdDQpaEdKOJ1/ZxiOOIFETVGmjdF2nelU
N//5o3QggF1TJL0v+26Xj0y+yI4RiPALMReWCVjMim6MpLLAlp4oZkBOHG9v/Yko8Xdr6PVn1sBO
mQ40a5xAQ9d3WIkSx77QU83rozkM+u0t++T+pVAg9s+eGo+rojM2QsvtE/IBMz8jl+jy6WRu1aEo
VXroYYW+SlYcpzl39tUJUgm1um+mdF5tJ37Z0IwYHhKbsrSfrviBSwq9d4QqN8WYBRIcPpDvooYw
Fivx7mCczgaoiJHujv2clY6Uakf52hBqjjM4m00R1fBSwBPkk5Thyea6wYtB+cpE5zpcWBSC9JU+
J5rJFlPYo0EQ079tn/mmFwKQI0Qxkmsf8rsW3IvrD/vX3mDu3qBRECMxrvntJZw1PxgMhDvqRiXt
5NNuitOaH0Wglt2TA+ioVsc9WBdA9NYzDaNv6ATrMmeYzUNDMMM9alaK74rZ+HKzMVNUW+Ra1M5E
YxvYbBFfwoHEhwH8b+ymYjKb23/tIkz+/qc8Q/63e7s/+kG+sKnQUGDxsxQMhmdkek86nr3mMzqu
pEixDvDBn1RJWI30slKp3L93/qbm05SGztrz4dczFPX9PZ1zj8yhwfyq4cR5TrUuA1ONXz2jUUce
+a7LZW5+SLYBgUlieSmLmGF8SnNaTMo8RQ8qUxlyGxu+13CaWlUpRBIvc702PbuY8ioRe+2+khyw
Q/xVBD26aMhits8CbD0mnyEA0d04IU0VJY4PyF/+CGHgdgupzABQXSEvbI2G1fritjWT012fFy4g
NN6fp/VRj6iVOJBNRdJo+vF+YIiiiDPHjNHcObpbYTf14A1IGa9TatngUM+GxFV/XZ2y00BRewI3
Bkp4G3BnERhtGEhSacbdWT8l7lhHZ9mf+QNfyINjadh0khEpj/dV+KbgVAUx/dIXHjntkBxdJQP2
44NFVlOrw3wPpCWlsQcMRVnhlvDdzprEFpLu6lnkyAZQwPheP8sLdCeZOFuQSsGZehWL20q4jcb8
BGsHv+ytSJA2/QIE4LTyXIU3zWz9UZpgnuV34Kx/OSGHTiirCJq5gSWnKy6FDj1JGJTqCu9AH4pv
6IvmzzE1mQ0nFAOmZnT1zgWfcf1SQxYuH8BgkS9vYwuTkpsPz11ObIpDeyJA4kqq4/eDLzHlIjG2
CbANNB5WT8wpx5s1fwEQr7cjwIGYPAB0iMKWaoUUCw6mZrvbfZqNTgzk9cGGPkuvSjTOxdNyGgWY
ynigHKQpQi8D4hikqriwOHZYJy4uaAoMI+/UybBOgLiFntGKiJYbOL9h7S9WKHpEhsVjnR9kmJ/5
tQ8+mqq7QaG/YXmUlW87UXFBEe5B0OHx4oLuwVAbEvCEJSl9MzbclENvpXs/KZZ7vXrcWhc7Rl4Y
dHw64hBGtFs/wFx6ccv2e08WytZVEDt7T8ckMod4BB24P61zApbVRaR3xqhl76gSxu2eSDVoZEkd
EgQA1WWTfCpkXHvG31TQWeK0xTGUJhfDJScCffZv9NZ0KHeCyZEHW8RrahZSGWT+AGC4NTfuo6aS
D9ahygegKG1ziwKpjfHy5jjNKF8cY67RungEmNLO/4pAYj6+hSyB7nx1ojKtJTeAhgWyI5VQWlDG
G9vqNZZro5N/APclenL46G+xDXqPh0skU8p3BArxMj6Ui0zRLdhh0HWNfDYgdHfWhiAiJl39g881
P7Ohrn0k1L2XFWD/mf1qjCEFz/9hNSPPFCBL2ePlJPKiKBX/7q9QopuqaOGPtqrGvW+6oe1cMMGr
CRdnY0eGGh0oThwsK2fuZtOcmlwDpUpQHga5n0p0CfXUqrqisehnsFoW8Mq61lE3JUiMhhbn9BHP
YAx6YUYCRQCt+gBG6CLVlyCXjyP+7U6J1Cy2bviZcSGbrXS4ymdg+K7IRUTrS12IeJO+Sa76OcSS
gU6+CkiYv6sNM0KurJ/7epJfYKRh3Ox1XaqCb5sbw7wlPR5OxtUtpYyHPKXMnqk1jGWC7wDYd4gu
IZeJtHXk8V0RafkAw2DhrOtX/kByTNYXSbPTkcJBhLhj33XiWTiWuLbW43g/8a8MPFDguPTp9Q8T
BuIrYrW3yBf4E/+AmABQlm51zBhp0/MZ6QDky+7B8VnbzHNBRt113/HQVQftCRxNwo3xZ3CrInd+
rI8iGDW/Z3nuDJlrluTholLq/mhVOw1C6VfK+DvV5asAFZVp8aV9uYmO98iEJMVwe/zzrdiim1dh
plwC0I9H7+L5TLX849f3BS7ZMEQzSlzJgrbIrDUBbfgaQyHI7253MJ3yRCQDI7djroxAfN8khxPP
KBWC/7Pjn0dG00K4+blFfdtEaPB5eUjUxM7Iax19xJeuI+3PG+XiwUpsVP+bSrZ2P6PV5QzRYJem
ehuIfbjFiEA31CqP1xZHVqZB9f0xppWu8oGs5kuJG+bRPHpL6u+KZWDmRN4NkeCtbYNyv31xYRA3
OrLgGPGU4ydSubrJoHv9anIeh+GH4iE6SgwySu6QwQgwORo0JQi4sAOyTvnZeqBVIKD7S4CBvrO9
Vk07bKkqzozpzu4me/jikZne2YnYcHDkOlsnszmR2AaHZu3lKqh7QkydG68Bh5sQGjzRl4wrlQ0n
IWspwzjSyjMbrTafbNts4QI73hqZvmaQVfghn2bqPtKbWh472+5JUBWYPGchAC3zl1IaDPJQWprL
zEqZCYK+/ScIod9yAybluT349EJiX5UTLyschvXDX7XZR9d07OqY/GWM2+FgfWueXIxLFCFsPVr1
UadrW0xaXv2SgaHXbHDCJ2iPOVLOT9VExzVYXaGpYuM+4UvKSkt3PmbVWLGb6Fh4J6D91/rt8Zqt
MG77OVdsXCu1mw1Ha6x1n22yKZSuoiugsu7GbPPIOzrfFTwDuuwIfkJXc0aLTFNY75v3UZjo63BE
MSQNaUjcBfhpGYtVGyh3Gj5nBN9kjRBV2H7iCEGWf8kmXyNPRFrkT+PDBrh9JNNL2GmXsd80Qb4H
ceww8H4FYe8w1TFMeGz5GWLGfrLLvUNFaMUL/8wy9gbA/+z7AQ5TrhGLuxr5FMTjVc6CsK8yE9zw
GdAvNae59v1SLKeuyoPf0OzbVKisQLS1IQVYoK7CV7nxdQ96dBJj+231lOR3VHafTm1jXpTwNz8d
5b9vxFSWWO9jdWgmGqq5HprmYHGBuCeU5CHCe5f+pWGmCeLbIp87EvmRC3Kn+pyPDG+q+TP+HsjX
SH1caskbXNOyYIerQ7oL82u+xA6A2HCRGotyvIYfxHJ99/F7TW/knj3ZlBl49WcQGtOX6a114byI
c9X3VAygwLDVT7+8Lfy93gCZHnjlIJeDfv4Om7FFQsu73lzSAEXfvqudanIsj2ckDWexr7lT2Ihh
M9m3zkEPPYkofw7Eeo8m7zCqx0CfDppbcUCFaC3Q/O1kKujIItpzBxnlTn73ku/HVVGJAWXK7/qB
f3fCouDoF/7AQhhUEeGi+Jf2T05AT0Egm11ImL8uJOi5mQlS4hl+XC4V7eyZhwUBzcc8dbbVwp1Y
Z1VnRusOiqixspBxu9b2DW2CFIwcGPzKZLKzijDSLOxpOb6GZJR0J+K36AxqgPV3SOYmKjxm6VL0
9xIW693Ll5/TT9rH9UOyj3poXFgwXmUSsPgRO4esrZUz6cxDAQMv1VbbGVnIgnBiLs/D1PVb8LOW
c8BZVk1FWRaHHPFQcF4hnoLqEJKYA1JNL2FkBHWzeBIOXq2YCZJ6B2waFyfA8jFCJOFN2qY35wXc
StlSGQJO6vpikTZQAUBs3p5UX1Usm9RbwUN1Kh7CO1txBUcLLwMAFpO95h5/5hnzsXNy0oKPLDMA
uKo+F59OLnEq6md++NRtwAtXIcpFqD483OURRw0R9G0q6nrfk/ByjODiM1GnHp+FYtitQQ97LUC9
trIC1EbRrejHwvDJqGuRTn/NFoUH5teGkCPRPql9Rz8Fx1PWrz12MhcdKNz4kfQXBWBARg7JLMP6
Goq5pmpZe+GJHLc8MJXjAmJw+Qco2rjW6X4IIKmfxFP1j37mNVEUquujRLOBdc2E7PsU50ou2EIF
/HJsDkFcD+YptllewuntuDjuJRQJa1uYii78icUYrT4mSzVL3hx/oLO8w355ei3kA+EMfa/EabQ5
CM/cOGpmIpr9mI+VaGp59bJVhb8TjE+OF8ug5wz4iZcui11Xg+eewoABrmrbAdSKSzZfVtvplsGF
u27BgWSx7yGMf1Xj2oVD2c3jS7bAHZh6x06moDsoayT0o3/WisDxvYsGLRSB55C5OvQwLgDrkixE
TlC/Pu08rx+bFjhMQQaHH2S5njmbTfmX3fcfapz3216qzxZ/JJ2M5bFgXOvSm/TgSZ5T4m1gJWZl
gw4SLGLkzmZEVFxIMx+Eh+jP+DFvlH1CSifm2rJ/3l+27bwRu6UsIngpmT86Lm6ywIQicvf6kUzL
gZIJEXrJRFDnUcGf4lA3lvsCftsY3nwoWnRyrX3hF5QVeZgqso7mv1CaMutbA5F4dvf8bCSllO/Q
GAkK/w66PrdHgJF5FhmvEi+qShFKtiOJoTXwD5NplwXSsbimQbMUYWWArtYVMRM1gp7j7dyUQDB6
SnAiGfZO7VhffoXy5RAoqSsPEXejcFAMqDPg7d2WiDCSOB/LEiQvNMYTemcEYmOilj5CEw8VwJNN
Wk5uFyewxnlJ1Mo+vgNdVQnH+nS/Q26oNYAkenkz8XZ9ihJKNjazk74sVVklBQhnzNDLbWlqNJL/
KO2CqL9y/Bze06GtYKxzbqvwWUC3mHFsQRUBNbnsv+1fasi1gGhfb07PSCEJatfw/bvbwpS42A5h
qRRIhpXwgoa0M709/j7hjWAJfOHhi/joFGdqPgmQmJbckHxnFoHlq/bZSrmPW0m75aDJ3XkzTLlm
2r0Gp7EsnclsYKnOc/o9pEEWEpW/TTD+k7n6oNYgKBbMrBSvgNIO0QRQyb3XsalZ2BHtK2OoYS16
+S/pH5GxfrmgjZTCbYsFeosDjUmRRr9PxsoTsHxF1yEOhTZzC2p2RH4oYSv1A6KYhbhkjP0AyVt6
/xkmsA369obLoz3oxWn7V8MkeNG7ETdSK9Axn4BuL/wjY9oUpFDIJGML4Mzwa0eX/gXSb3QobEZ0
uIwNeu6uAk0c376ml27khGeGck4hbdpXWI+HJasez4srFlHqLnWtXH6Ern7G4A3spigQwls6LrC6
vJwwWdRB0jIshS7MbDhBTtPq6R24BK5Ngr/iJa95FE3FzwAMsi/M6vzf8NsMVJil2r6e2EgHSOYE
7LFqw/VBQIMDf4fYbVW5YXHWR+cZXyczTAEAWHZhdNcPDwcyTLgC64AMogblu73vOcmNCIxlNx0d
MaP6IVYyL4eQbUB4zl0gNaMG2PjEU+cIWft/vkmCP8bkIIwMHNsqXQo1oh7169qfsOz6BtHTOD8X
H+K3zfomsY5jMJ8sC5B7Z0ZuvNA4q0Bbk6fjwGjKVeqD7R+RfK9uqCaM/0LzcsQeR0K73aWjT6gY
AnQNqGHg06BERHnIV8U3bk4ZTc7EQVrfa2Nv0TPbFDol9gNUKaKrv7f+df1ZXOVbID2tUnb8xU67
JFpnt8CLbf836qgyS2xiLUXjSG1O/wEuu42D8bkydthSs9uP47bIV0BSGZbM5CdFudGM7ORF1xYv
RivSxljlEBYRFQXAWxJh7OeRwbGiKExjG0F0Tq+OCsjkHghoG9D3Oyu5bqqOgE5eZOvZFepHSGVl
bujShHVcu5xKIABqeuya4CCF470vcIlSzASS8O8LCFUf7grqzSHbPme+Ty+bswxKKPlOV6j+/OnQ
fix3y9YfxUG0wHDiiE749W1TYbtvslTZcnlXaWQ+cWur39R/js7IJjYndC9k0E+iot+nIwLunxft
ii+TTWiwvvI/YYf7eNK5YRvAaAoExKYDSt4O2VrepOE5PSuliXPafvFGpaSM4kflXvkZ5BsN6Dk7
m8rKO+qE1AMlECnz9Cq1P+R5tkKFPw/SJxF1Spdb4j5sbZX7lqHup9B8qJzl1Kdk0iIwKSupBGe0
sKgEVecLoGXW9RlIHpuGH7ADC6y9weexYTJlOtMiTtGaFW7nZN6KLe/G2hRexulIkUtfX0a46DKT
I6r2pE5nCXvGWRi3EcW8ESiU/6GadVsVnLDDDUPz0JCK59QFRGivWlz9W37YXNRWkXropO3uQSIu
d+CfNP/kYyKtESOWZfSzp6iu0yOGHdLRwpDpiOGtjzEAiZXM7bp860uowa2cseyILbrSpkUGVF0Q
dxIYMYvPm9j3ehZczs19/lj7NUJW/Iw22XDiS86SEhxP9O0FzSxTE/K3GGDxhTc92T9NuTMXrlij
zPmwf9qfaLCmsJE5nsdpQgJzG89Yg16sI40JlO7gekF0fbpKk0jMDlJZfohOt/8bHV/Frte+wXnL
oiUXmnEN3jtxlhX+r8+qvPGB3QzFwpWdVSg3qviWE/3pZbY0BHziEqTlKqdaNBfXGkxjrtw7YmPz
q7lQLj1eoCg60a3ryS/tzIrF8DvdIIwvBbn51CRWPFc77toOBbQG9dtuOHCdQpQ/JF1u8BO9nCkl
pJ+w5PdhWnlUj5z+ty9y7l03iwpK7NDJz0DJth53yqHojT6UPeF0+SUxDHRgAIEzQ8G5NlOFDtPA
U0JnXmGZ9cqE/+ccBztn6OfsKu6gujitkS6Lel/yMqZyEemUv636LVt/xzZ79Q7HWf22ChHidx2x
LrWQMnAKNpdirKhQlKr0TyE1rdmUhuJ7AgXIpUr5AnfnhKcnXb8k5jqO2ss/WjXQET20otzn+MTS
ZpUGFRnoap830986k9EDxThish6+JrmanOST2iWZb/Zq0VtcbDHO/GR5qW++VaUfq7xN7f+ckP7w
sXj3rrs/a9DzXw1sN+TVnBPEbv5qBzkMC2c5RjyBhhoBnkmX2pkNl0waJcav/BDRI9FDBnJ2bIEY
h2NjliqepjdLDkXyXnVsgq4IZ1Md9FpFuyVlp8RqqfTxt6ov4NGabr2Hwny8L1vlnTVNaC6nRYGk
vVFeX2HyAnpF+qNpPHqkZEOgIYL9tPimUZAEdJFreMlHdJTz2JDh6T3i0uLIxt0yxXk6IBDROWLs
eqoXaMkKkAflUxwL8btwiCgqRP+tg2ZH0dCRMCzqN+PEBzLJe7tie/fPsfaLnKGNbVxi5YpuORH2
HHKSK7GvA9oPEB/d3MNbqXvgzVszYzjgWOUTTUGPvYZs01X8aqsKfONwYGx0ARWGOZz4Fwom7C8e
qUqwqRq1cTfJ6t5U+8HIkNmUJt4PTFRz6t2XJtmjf0e67wCBf7LC5WIUvmO9KHHLkFe57BRjlzp0
y/9z3lPOMECPoEL+BPfPz5uhIJKtnbwjWHjsls2QUphJra++c0i+AjXhEmfrebVKplKl+MAlxjIu
hzqegBgzpJA+92vZwA7injrhZwf61/iF5ROjN2qEXESgXS/Wpm+6O+jZ85nOhFeOExvVqaRz09wb
IVRR+VtRtUmQ2NEyh+l67dSdqBpGHTrHq7qqbSylcDsjE/jXmSeOr9RUMk5vE/kDzEcJjcawA8NF
030xAbGtMYeZP5x4Xn8NsRc3exOWVS8/naCFcYHUeE4q6WoNyj/oVWsMjDorPANPwP3lIHxaNIXL
BQL4m3C8gNe9noKy+39uRINuMUs1Xgfm/2Ri55u4CTxwlbUrJj23vpVkZyp62mm06htJl+ZNpvag
jKQn6cHArsWCtjc9NeIW51uGHzhs0sOEfHvjVOpOQxZiKGE8TEKBg9DRrsgQMyZquB7efE8psoE4
f6H8jiGE/gTXKhTY6BXPZeqynYAaN4/pv3XUhqSID0Uodxt5tehqh4XlvadI/H/FFdKykQKZn8uj
1fqyCluVnT3P4ZY/ZY8AXTUVYTcEDP5CoOt4r4QmYhfdd7qUjATTX+agnN1aiZyViM3aiwbIKTKx
dhRiQysrg7V2WchchQcht9IVYvaA5mS1WSf/F6XxfWgRuH1gAYjPK+hJ/seY2qpS3S+phFApC6vM
b3gIl6ir2rfs8UamQ6PPaqi3pktpOWbwYb7VkNL8FwKKqDyC68zD1RdRLi9xbDElS6zMzLP2po30
963skGMI+rmNAyVy0m7p4OIOtgdr/6g4FVEZv2tFY3aLhP3zeUfA5+xlix6k4L/2YK5v7EVH9gok
UKkHmVumrXzT85CP27/sKyGzQRKcwtFnYnqAFdxpXcUidBZbACa3Xv2GPifxHcaJsCLq7+NSXn+r
SOTHBQQlizy0t33lgWUIvvaiLCTvV4DuSh3EgOjzgmVnzt6LITmkrL45SwbSU1V/WUMkJH0mFUP7
L9y6N9CTv/sMICZhpusPZdZk+8E9usZUbnXcJZf0D2n+ekyg1YrcYSTPbQ86MmEToR+V61g4ah0P
TstW293XwZ4pbV2le7RSMydO7Bew3aX8TkMBWp3zCLiVTUds2nd9c88XON3rWUSsophUj9rHUykj
Llx+GlGO+pVVSFO+RMxlP+gpIJSc0JlHGpB14P+tRnThbVQV3Bqnn3z8t5zK5Fark0yaCjBl4Lvr
DT84pd9qKMX8W2azHyh9Qg/0yUpunEv+FqCb9tjzqwsUjdPQjqZbvn0EmkVTxV+DsAtRo3Y2wIUI
jEozWo6Dy+/F4LRO2l7ZBRdDtzlCUfiSDyEpJ83nu+TxJptsavcuFndLyCExptAyRLwmURuws3NQ
lzHZNOttQnTr6J21WGETHe9vX52XI0pK0GYPyFERW/YJAiIzoCPr0G8rX4xYhaLDQKah5ACwKiiO
XDaHPPHQBySWyi8Lzru391qYHeje2F+ztcq5uLUx5Qm7oJazOJEiZxGh0Rx5pe+l5e9TPHXFjT1X
RLyWkwUzymde9OqPx5cer+Gdfw0dMnGYuf46V3eKQ/2NK3FMpOM9LNliRlDd0S8sagWYH8GCQxtf
3NclNAPo9vqPpj/+9tQn/5LObDRsc2KCFhyHh8Bsb6d3/g0z7s+Tl3BYYbkFiR47ocSy9rodilth
BEcHHB+ETuL7Kav+2NBTp+BPaL6J4N7YhTi0X8J2HXwNdpqsKfE/4DckbPa/YKIxdVQJNDBsXWUq
F2SI+Kf16auCchAGdZ/vHgAzgFxumq5xwOi/O8Cn1U+Ea80vQUfhXUZgqBW6sD45WNF40VVOCT65
5nLm/FZeq1xkYDRchMXWA70fAtmtA+04P9KVUDIE7a3LUCtyrmeTJetHpxUd9kCMxlUTKeM1Nk0z
69IsgPNqNcu0kvJGNBsRyEjCTVyOfpJgJrqxZb/+0iwfQA0vQgmBRbRbcPAqr947Obt6/hia0H7Q
eNOmga5az8wccQluIQwDGcJN9Yz1H3WRcLOXXU9y7Lx1OYYONi6EBODO8CK7ZNgLgCiishUEP3t3
zZyV/2i3QrId1Px/BufuFpJzmQuSa9Zen5S3DS8gf5AD9YFhSR3WjB4QoduB3Bh1QUgS0d4Ms+qH
al3uxgAIrjp9oB3Fiw6qnE6uOePPrKr9q2BadrpL4nfGtpINjhe2wcu8CODgauh1NJ3+2NbxeBc9
QEELA6GD0hzvmyv/KgXGntUbf4rK1dJIkN2ukjXhspSoqbFp10vVZxewEWXn0yCsP88EKYv+ocNZ
9c/XP7zjXqnrntemGkv8Nv7ozQaA4Hg7fIjdP4PY/7uz9UA0fFT9V/l4vO37oZkYBZVVWT4uMUVM
5spXoGv05JUjMhRP5G8deysjrwCjLVqrMowIENOAiosx/fT6hnF3/s1WpnlwYKu/jsABzoQ3YO0z
O/7MrNEXogKF/Ma7pKnIKvakV8I5n3etzmswrQEUeurDis36rbSpMGsu+XEr6kIjscHAe+bfoO4s
HIGQvyq6sSUlIBpJvbxdu+7n5sHYTH7h0Iig6H/Jgqh/l33VIbMqTlQvduwjC9v90JZKAhwWmrJL
6Al8kToZYCag5tvtREEnSZn4oGSbsI0XbxYOO25Y1/5kLxn3dXTDUUTKeBh+sHbuy9U0Elxy0US8
3We03l7SzIE576p2RWS0Sym0KDG4KB8JNC4WmCTMsC+PKg50auevIKvfN51hd5dWJ8w4lPGNJWNN
HPRiIepwGPAOniTK2g1evs49n/u2VHl3CH9W04uotogLctw9LNjKIeCykWx7G5TwNhEATis7g/oU
4zI3f1jWyx7ivtp66i79ydhCDX1EmGw40BD7I9ewvoTGA9ht0v5M/QBa0ZhMRwpp5f8wWINWA8X5
ncQb0WkIQQ4i7st+TH+iQ5xD584v/0rvCuSVukT4tPAxOTHBPl6re4G38rOwOlHwS7Yw76vomIQv
1KUSBoZ5Vi7s5D0F0V7nC7dz/gQUoDk5PjkQYzbwtp60yffzAJ4dyZ2v2u0h+gsyKTN6ijmYCr8V
CoRBkDDfk7/vnIZhRhz6JTVww2SR/pG2/0WFiBo34Mf3vQC9IlEEnk7+2IplfuIewkCczdmYr8Pj
spodnhreFNXl8DQRsUAfafJNgmB7gNHbqpJN2gmT7m2xub9Lb2qcfY/kKsOf86+dfhEUUU74L2+P
gf5DUH8x8FjISVLNsNPzHJr5qkDS4TGxjNC+z2dER9vs2xnyvzlOTqXyKyOqoesLVurHOu+iFOEW
HNXTyq10Hhf79Ep4pOB1IGS4kOWCR9DZ6bm4k+goEDv8fqPqYwDJw25J9RfhL91mSp7guAfIqmEd
5qQQ3kEXy2iuZYH3E4gBMX5r9OSL1cliOmELUb+WfEQYyjn4/eBnYOoEOG3npsxQ9c8JOsgjb65Z
dYWIal886aP8LPWLYstm0l4rkEWWSaKaIjG+4h4tkemleVEtnu6VHq5OV7PmzrJtkvJT/DGS6g1s
+u1F5HwiElpHatdcTDEu6LHliiRi1dPZXYBuasWEU/GarMKSPfgENR9a0ZlZabfaePfu6HnNjDDl
zjsbqTXhU83lBWOz8t9ZJxYalKCYI/C9OcEh9K2yUXkU6FVQ5ebpJFSFfqT3i6hzabgq4Ez31TQz
o34Yugb0qt0Ey1C6qsJlk16fu2Z/1UzG+62RBncKQmNRx35F/YqNoHr5WBOUcAaLERfNtWzUUj+6
uJaBW2nKDrVb7hYF0uQveM+2/C2EDxf1fDlI56SwpIVvCfX27rtgHf79wRxnCBMbJIfKrFsTHJbK
EYw0TNkL1OC0UFK4D4yn7uosVc551soITYL6HQBrjiGXY5qt2lVexzRoFDDq6vqCXcyze/qDp1vL
P33JFKPH4QAaEcYkvTRUIyRZPvutzAY2k9pUtS0l9mJbx+KQh8hxy/beTXeVYS5G4YXUrGKsFalQ
lbmYXjnUGSpJHFmoaRo/NOIregrNbHBRk58kksy2nycw4MBrf+RXN0iOY/2Kn/iR85aOays+uYw2
qtogd3NzVzhf0uNPe/XUfcYgIqFi9Ln8ZCCW7qSJzIWWKZMXhiP/QK4SeO59NdRbJsIHdH+SJuRP
Sl2un/GJlh+d4/U9ckNyhUjXW2C4kRgOv+ZCVJZE8Y14cYc/oFIUbtATth1lclHbIVf/6RLayCNA
EHlCMOJOMLx++hkVYk8bMZNtxPwFOHpHhQMgH+l0OA0ZiTli5/foiFOyoJ3oI79ItPF4Jqi/LInT
ihNHzZOf88Jaz6mWiFuenYqJfQecG/6ApgDG5MELsMcWTuVhprmMYq9sV8tiqTLqa2Ru0sCm34Me
H+4PREOzo/lA4fSswRC3SLBPCCgM7Gh6e/2qtd8/rkcXd777WfrhU2Pzbmt9Fc5rLqdKIwZtm6X3
FXkhWg2DBjNi0j/g24AUSXt5OgbmI9a8651UxyfApKhHLv4zq8NcxoQT7pSmOlCsJuAvYlGS6i6X
BrIlaAoqvLEP2TR+38xWWQd6hAV60p/Ct1siZhHhUj9MlfTMHi6e4D9zEUWExCbuOpShfvygcCxC
QOZ5nsBtrFpI6kXUPw+CwiZfOGqG+5K6rlyIvgmz1yjCyhh0z33HAozrkKxClzXcQp15e2o/Dbb4
9RubzePyjkVYhxdUm780BiRMus46US2yXngZKPrm0FhmFzYkBPAqhbkLod0xHN//OVVKVflp5ySC
6NL5CdvatI2kGTKJRrKo7qHlCsWiSFWbapo9O7BlIdpf6NpJjSf+Q0YUeIg7MRBVhNNspbtXAfyQ
ash3Mpf7HboyrCyZTnQ98kPfa3td8clHlpG4R0K+pBOjOhgzTJd9bXzjZBjszHh6H1Nx9MUlx3yd
n939nkdgwyMW/vSDygU+1J1Bayd3cPaIy8oCBTKmhuZAy9EaWo/OUq/bDG2NvJzJ4TpqurwmF2H9
h9DPSa4RQmnMoBOOcGK6NzFMpcx5UCKsCvcpw5EVjkpN940KOE5mm3hnvYBBXFGkTlp/YLacZ6wy
4o2bRvxF2/VeSpZrNLB8f/39BqfSOV3sLVrZxHKhvZdY8oR2ZpYEDNz6hoCEgBR+j7v3Aqg9W+Ht
GMBQXZFiSYDIkOJMNuM/fCTx2GDGbMkOmfbvvOs3p+xUBwnkna2NLCquRg3mi2Sc6kEzboqilS9L
l5vf4iLRBF3k/ULAFzE9BCt3KvybJJ+O4JsP4dq7XN0RUvHlsvtKI1tcHU8Rc4biFvAwZgnsfZN+
xKnl/ILcfPp8Nu0UChY0LDWY5i06bUYegoMnSFQ6UGIhmCW0/obyC5riL1t0rouK3EAMVpx33CzC
S4FPqSMGSCnXB3VDluGGczokCVqstdtoMqjDNrCJiZrq3L/BGSZ6t7qo2qwa5z90IpCIVZvcvc3t
DTqicuU1D2snamxFPg0x8sNNUw58RP+gBDY2qI+Ms8YoM4iyx/FxsevrIh4fOh3hMrItt9w2rGPu
wFF38SptKG8LoVVOqRrlJfmGUZodM3QklQYkGohZJce0k7daaagfbvuVgC4upys+XKHIi8XWPi4W
jpKqfY6Ip2iZtx5lS3brINYiX6odI4jTlHuVAOOgiOC8wvubMj+Rdq8MHvSugRIsey0eN2ArvJSm
CunKFPYC0xpNNq3o5/UwfHcnmTpCtpnW+12STPmKoYOXIViuHCVrjG0K3M7cTIHIZJZMdyiR+f7T
xYYB91gbwGoWM00vK8NXwFkTp6ZHHfa2KAQFIhuRJa4qnrGDYITEorODp6OUqF+VFcX4Ab8JTBqe
6KVPiSee5ejt5n+hH2JuYwp6HTUwLfh+Gzh4MZwth4O1UiFmXcY7BT3PHu7q6NZdCVkwrb3qrfZu
6I/ADpOghIuNJAwPQevMbef5gGLHqvmHe0f9RjVBdPMhiQCkKeu644bhg7XphQExAUQz5zJKyhkc
Bzev/dUhYCnz3oEdAdH12+MMG4ZynVoq+OJfj0qssgw5ZNpeNc+lHoYGj1u4SydxayBjNbBntkcL
UxRAMYhufgJ/kziAjAtW9TYw+CxWcX40ZnPTjl2N7jBxWyEOARzqXjW+BIwSOsdqB7CmnIKuGamp
FGhbl4LOzisahoUAS6z6dPdaaE1TYXiSIfs/mVkXstBFIOtiDOfv1pghplWlgJfilipg9Pa6jC7A
auB3To1KZThfdQUezd++73LHIeHYeOilrm3VVLcbaBgeT3ooZTSURObKEPDe2Nh8pfTkrrZbsreR
YgF3jQSMhQKzvx5/hGby07lToJgbXIpl/qrUI1c0mFSQjpKJ9qZWDJwckUWh7t20R/RifE+D/A62
32EbgCMgWWMSN9gVkOoG2y5XdJvtfQ1fE3wBNOSEgbIxvtyJD3JfMJe9vI10kxHhekd5fONuTyyB
laOCcgNylZJTch00WT9vQOp2k22g5t8cqlFPXXj/XwpYoxi5OUpketXf6aTREec+mQHT6K1jnECw
i9lfACV6LyOAehd3Shs1XfVxOfoDvfFWTjs7nTonxo03r4k1XqBY5WV0imJIs3i61o9FhZ+z8XEL
7Wjt9mge3adwPUJCPbiRTMSw+KgKputpuR/TwAiSBBdtHC8UAcb5st89TYHCWxpUwj15Y2c5TeAc
F6zmMzlbO851RIv/YB3hlYwnUcLsnfN3btP1m+BHkcJ5gUTARfJk1lbc+fpH22xfiguN0LCnF7El
Do6GRHprdRQTaIjZR8z/ksy1CLNDAhIFZt778D3DKqiRrU3AzZuvZwwDy/UEx0J+LJSI3FxxAbph
iwcAtHDb1ZRqP1IgToYMDoomkBhrKHpO55n716BDA8ORYWwoEVjeRs47E3H6iDOfvbBb3rIzVjww
zcihgcouyiBHoaHzM7c9K/YjEEyAKfRL5iPY4ZXaJutu8KNqL6J0hikkZ62U5bWP9P0J3JS7i2Cy
N4V0k9wxXwB6DADJJqxR/2PWC2zv7ECWnJE10SDhgyXg4Hq79vMV3CxyytgvXtI3JimlNY91nLHc
Q/feE6k/NHYCG+FE/GeTurfreR2/OiKbwXXv2m9xmgbEHFbHD9i9f2e1vlwIUmUjuoVejingAqSe
8c74R0jDsFd02K3GsUdeviMU9f68Dde/UqWJnHfyqcuHY7DabzPa/He+epiABKdqqV5K0FWoONY4
GllTTpq7g5vb/IKS+Rtk5L7oWPp0VfIH4fcozOOamN/cXpYJEciXGChRWHWqvHpum1fl5EoMzDw7
nZEOTENAWlW0tdZ0/JVXPJBBNZ4kPXsrPdEUqfOMtbpxXaH3pni0OzdM07k0Nm6LZ5/5BNDxF7Nj
WXdMhJhop+TsmYHOf+JMWhlGOfpYl3DfNZ/NXWThblrtZ37MC9EwSe8bybLEHkKsVpiYuLOTReiN
+YOj7SYQD27Jz4MNkKs2WQDR1V3FUiQUCbZH525PiexGtTC3+CiaMzVaMM+A5TSVcUw+iWAz7T//
HCznmsuDl+tRYHvpicHjJAWpsounJlMpY9MTbb5Be7zQ/LJkKkA/qBSgv3k4pgGTHehkUTigxhmc
NObc3pEN3VFh2Ho2B+sfaSh+MbrxJsd2MYXnKEZpWLohYthunR7bgmHd/33hWAHnKTJllTdm/trD
k66FeqtcEgevFi9ooGvbzsBq5KuQik7p28sn4tOGt1sPLjeH+4DNqcG4NMDAexztsPABIkOMTW9L
/1rQtkgwcrZ7bks/aLKv52A+vXKjuwlYIpPa9lMLxhz3pjRyZ+0XLbd9p74oGySc7R9uSUZv1KKP
Rp/vo7bcYBcROGi2as6sGFPcyho58Q7DuCUhS2e1XZ75Tq4mqJ3aJPrF4TbWNFKrS9qj5gZooPEg
UIrMth1zzlvDJYu9Ddn015lMTDF3YGcXcScY4dlVAJZwCPOy8wBbd+tZglGidjAoDxeLytt/zyOW
b9E9yaJSCuJzfAuBseq34aE+HhHgGhWrQelEbaDwz6+xgCLMuq/mi9Cr3QZK1l4Tf/IyoOHEoHRs
nCS+se4aAM6HttNZHwEBmq8Zd4OfoQDSldJcS3/3UDXs2V/8aPf1u6Oy7TgHgzbtislwowOJWit1
zLQqPFqLhECXV4S2zJPQ0LK3IveUNVOYregNwzETI+fAt/IG1xBN3O1eZ+wrXNczq8XE93U0/R4t
Y41momnlFEQTslnhvFvWZfdYQh36T5Cn++X30ttrDL+cWxVVyT4CSfc4xWhU2oT0dumT3RQJG9IT
ciA/G4H7vKDSBdaVp5O59I9wOVazyRfhMAgCRn+PDGSQLG93SHgv4Vh4eAF/8slMay7j2CpkYK3j
30lIMEjPCvuc/4yRBztulqex6uWo1SzvJUgh5y1jTY4nsq6HFm9mf9t28tCjhijOp7kdX2aN/+yg
1fGpqELQgcS3yiP5Gj5RpCSlFEuznBe2tmYtQmQaSQNvfz6NS7q+48ZU1hCXxmEZPVgX5fNg9KO/
CkS90/JVU0Wq7jTCzCqWA//gdoFTX6c3GZlR8OC6V6dwlsPfWihFs5oS1fOvN8KtUCRFfSXw4g41
BG8Lvx2HTi3RzWef3OFAsy6VaQT/ZcHOaXK4OUvzX7C6WqGaR8kHkr+bgstSYBGeDXHa4m3h+eK6
3p74I7ubJKxFwYHqooVY/Nb8iZ1mmnEP/rDacTPLGqBV9Dya7BXHxDj/IZ4PrZUwN5ad5CoXDPAJ
HZcXiwY6XsiN6UXWBogL8e8T2mNU9TWBVpPnI7FsLF5a6lhRIrn1D17ojTeGzyw3Z9hREpovWyAx
Qj9UxgdF+3yeonUlFxoCTr9CcZPZR9StkHUaddXEPy89TuSClDDKAp8ipEC//inxGHvH/wF1PdLh
Wl5XGP8yeybxMaQmrjdynL9Yi4XMbNTaDisLh++WHrCH6LhFFiTpiie1sLgbf96926vOW3cH+FpO
s1wcG+H3yfHCdttI1ffWZ/koks13Xxh3zedvGrNkyF7gkZgoTwRrODzq6KXBQ67vVhb6RAAMeTrj
7QFhZVwJYTMt9uCJtK3nLanpLFv3JHftkzTh5xa7t0bB4qXDgOvi9n1Ph3mMb8i7ImCH16MDWWKI
f11uQeEFwbFVfARSdK3b/4Fr5Uo4jQijbUIVQKmfF/I2QjtiJa3GMAZSmOF2GiPZwnQl/hM7EHrd
7m+24/Elf/f6CHL0/LgxTVvJAW5ahJ2wl5jkD3+/so7+LpVeHoklY71tmRQGm2Lh3vMSCiZgC6cQ
Mi00RXFfAHLU/mfx68c9efJB9OJOtDQKe1lVQ07U1mASeqgy8KLhQAsLvrvda3guVyrfyJBQQI7G
frEX1O7VilH0Lw5spBvOweXoZdZ0OomF/uUC4WYKafpw+kvLXPgW7XGxV9ffFkbiV8p2ctujhvWf
ufewzFCR3uLqdAQ3Z8rw7E0NjSD+/JeDVPkrP25gUo0Hp44gBjlcC7LuK1JA1xbP4AXyajMMJt17
72wikLO7/gNCsJnAWDZWDQkvyb8n7HvNpy7w6+1Sjxe7QH3K126M8HE0ZEPnxOAKRDSAq3KBoJdo
RMy6thZoNKLA5nVPSBf3zXmg1eH2aaGiEMaOH1YVI3RA+sVgCYIK0V/BrYfjNdHG4aV8TG2uarVz
/4l6PXvXJL2Hl7W+wAAaTA2tfnxNyuvPa65QqmGDXkbqdU/+XorK+qgqSna4tJZWh+nCv6yXykrP
DibpGrRkK8QWKBpaCGKVpuCogYyfh6z/gpuTtHijErsRcS3nvK/GlYSk9wSKuA3cH2z2dvn/kWfe
QCRhqmB4zZ5zUOFnKD/MiCda+mefT1WCzY+drGAp7/nXWzETZGHFQCnmSqxTwlgoSdFeLQufiC01
i6reDrEpW6RakMr+9xBUfKy+JSixFSg9zKqKJ7KDyJk6ANyhoYskTgfI8hVwAZ6IDX/tPqpwklnX
KFc/tRdDlyLjCIK45QTzwxEveLNSRmRM6fdzdJ7IGE+SIcyj2Ig1hdANri1IKhJ+USK7r4aYJ+Np
e/e7OIFqHqQsBxE+6hn/TvMznPThokj3NUluXkxHcMb0MQny85TSxKfrH7Op6nXVL9lks8EjG26u
6OQ36ukQ0rDx/r/MVaU7tOmm/Cjj/F3aqVi+2Cyalc2xgg9zfxsIRrYTcRNmAwe9ZcEW+HStCzIy
/wghLvCBdlb+cwfa/xJFjDinAVZ1Nu1l2UhBbcUwOJDkxqwTntFeg5Mz9Pxolqm58DnQsL/Va0mM
UssCAvk8TruFdSW12m0xC6RApMkZqo7pD9NjccbORpi/2Q+s+DP6JGGUzwzJls9asrdbrLxjl8zC
W/DtGPZF1k8+hXj7JFWoLCW/yH49Z7d5izXOPnKFezGqetoIJCAeZGLU2f2qXDPyLHS40CjhYdFt
4KS+O0+MmrDtsaxw2KTQEOFUty68ss0CVl7v+fIGsnDKYA5HtfGKGnas1V5HKqb4m0RXTCasUaXP
nLOkD4ocZ2rxfF49ePPGI7ThQ0qC+9nCqsAGbCKpXR6LAZMYGiKpkEhLs8ZKS/R+7Yl0qBRKRsLB
vGODsCWXp0YpnPlSZ6LySSTemKDTZpenvzHjF9ujpWKSd2+p6Mlf1GhpK9sFExl8NoEBo7paC6C+
/cdHQGpo/ashHk4VfAA7imozt3xX+zVUu1UioAqp4juunXeV77mxNLotDr1c9fapyb+SttT7Gkr6
C0RI2WBMjK3X8HkRfa4GNJNP03LFiyL9r2wUayVy8XRTGb8RkHlrkKyN3ZqUD2z/bCTMA8HzUIDc
OQ5amoYuw9E2bxrdqY3h0jZxehxiJrdVPgd46cIOQF1z2CJ7+tdCsH39MzAen5qk1zaHf+FTcrug
Nv7GaSG2x9XgV7df76dwQ+J+QIEQT0NSpWz5vmU6xzQgcYe8iPQuKk95UFB2FYPGwUTrQawliyG/
wKTDFkvAoqujDNqjbE4XwrIFNUuBhSrUHkt5dbWK3PUZjIiZAWI6t5axArlY1T1IbGzVMGZ9W9uJ
XzTdf2RfIXbuWBFNVUbn9VH/KGu2kI/I7LfXnS4fBcWGbBz5teJQ5IZBLTptdMs3ojOsM77g2o7L
vcfTsd0KiM6gJZmzH7vsHAsRQn8+/SOrVLO93SIfVokK7U2r2bkYBPBBBNQ7fFi9ckvgNRdoxNhf
tcXUmVpCH2tc9ULNAnAwlmEYaq4dt5ua7uJUOs5gQsHHjtWYC1BWSRvzqtOCr3aXBfDG1Iwp4bCK
uHdg0U4KycSJo4xlABPWNSHuDpGq2g5qxuGgeIBKe4kCMiImsTHLM4HmBqwN/mjHdF1cms0+KLKx
2d2Lv/1Flq3ehrOiRC+dUuxcwZUaknigPTllgyLGZHOWGAIuUCu5+OmQDyoMZF+vdkN1vLtkCaD5
ycNSSP8o41G0pPxs1uffZ71RSJhsra7LO6+Fsf9rKFjnaEn+KSEUzMwK044rNeC3omPC5YJW3mlj
LF9GEicTITb/7f+z8Ch9ETw8026YkT/mB+xElfKviweMSwn/VoAykIB/I/5CUW6sLZE/WbYQ8SnW
m7s1jfeOdxB7f7G9Lk3kLYGainI06iaLLMmQCdFoHISD2HIPNfJ4wF7y7I9aUMveAy85uXABuBAp
ShL05TCv6HYllv0SRR553zAFWxBOKOqrvoZCdRVJpFVmWahzC+eJoVqr0KH0ebyOfswf95CrGqqZ
mYSJC9q6uHea3UVVf67AZbUVxkAYsTnaUuR89Ux4FgHitM2zBrSurn6yPK7hWTrL4WOeC2mDhWpU
WB897NC4Tk6yOVybLePq4qJPKZVgyRsf8DUgyTEYp0CxQfVO3ky8v5HfaFJjXU7S9H/9wO7sOw28
0sHZS2JAIcwera7Dim2rSnbyCSqNh83Ok6uqibUkbBudVCGbjneC/6I+FTIya0VqGBjP7UanCQVs
Bzq2SNmulpmYnyaOVCy+7vpDkvo+Ymd+SVEN+ahUDmmGYWpRjRUwZmMWe9ga36kTQlXf40J9dCpb
KtknDMyFE4C3Vmoz1xv8Yxsk2kUlCZwthwoV4EEbEYfNs4r/kLJVcKI/KcjRXJ5/tky2GCxcjcv/
1ww7QcuqIcLYrVVeDAHVEWY5rQnRREWn5uScs1v//US/+lKC8SQvZ68nuCcYoDU8q9hoLy+3PRX5
Yy7p6PVJSsf5Ap3CbpieIkpgMYkzgaZc5a2gsmB9d3L4IBtIAOWRNZWSafrPzzsVgOwLNMIN7PJs
7T+7dBm4ho/ynDmri1wdssTtnF0FNKfj3Zctn4ssv3udVypvQRed8blcnWpBpJSxckWz7IE44Cyx
B2l71i/msUxGERchfSZAjGlf6aPTwnN8GNygfEF0Sejfx9Wydyff8q7b/y+hYU1fhrY/dmaRINSS
XfqiNuHdXGRM/rQncRKvNk+7l5Odr7CpQV5VRc5LrMKJq7W0RZ9RRXXVzcG6Zh2aZXiyS4JLEUMI
KcYA1lGiopN8a2wGF7VVBZzwvVY68+MC86aGyT2j8fQmqfu/8aienJBYlnfWjTSARtRZX0RRN0tj
7Ia42iChdrPxqQrpPgZ4rlwD9futcpEzxx+uUPJ+abwlNmFk3inIfTp7BsIfdVS0vvrnGEw5oAfQ
Q0AYIuiJsHBPBeCrld37BEfEpgcz7YYdWQLMzI5+b76JTpD5+ojtOQgWMg3kTVtfbF1ovFmZi3Ny
CowR7p21dt/zCpSNSZzJtMLiZTSlgpbGAtMOKOZpS8LXklH8es+y+FjRjXVXKt5M8rfohrpaxCJj
tkU7u2ut6n4biQRBLSQEpCwJWzsJKfXV+rI5XMcJDnNgDdhKXWxpYrKFdC+eohOkdfMVFP5AaCKu
EF3pYFhMmvt5ufF06mf9O3bvwaMs1UkxP8dDZImLsOdRXzfZ688gi2XIBQBYaS2QX6Lk1xZPFDAy
T//aZyIdxs3Vy4oUrJBB8y+u6BCGzS3EvMwvqE4Bf78zm09GMRmbziWoT3ShUC4nNFlNRpbxkBF+
B+ckThbrMSU4Z/K+gg1rjmojuQh02LDkdSLQYYocU2pgeHweJcDRYtNobvl6avvMDxnmLV40IQC6
d5+xXXEQ/bDXDM10YeTGyqymA9NeTHOw5fDYo8B0Oav7sUEuuZc7mwhgIHFcoqqqd8+AuHFeQGph
l74XBpY9USX58w/jA83+ASW4Zs7v+Aw70b2PMm4qCt37E5PbjFjgom3FmxK2DnSEDviUSOBbtudo
0UNeaq5+0CcxIHxL8pz31HLlLZmHiI7BaVyPMajZK1vw77EjDKJr9vjcPudQ9m1FEJz/Egul+Y0J
Aa++6v/cpew7QPfglc0gybBg0T8zKyZ5yxdq3sIdOFFAMmaiTemK+HfYkxt4N8Aa3dxeK18/A6G/
1oERAN62+9m+gi3Ul+bU0Eq1//l1xzZJwSQmIt/GC7WCNtg6EMkGA1ldCIAw83rvBcNk991xcd9C
6DOY9wl+c/QxiatfpQxJPo0ejGKsgpksBjUC0cG0EpEnx9MOqSi/h0HPj5prPIiepdLwpipYHUJT
HQ9mLd/eoAlqeltDK3XgnNUHZcmEgZFu8smW6L/WsAglL0/lN3ROBf23kYOyz/xlQi4znX3ysLt5
6aB/flH1sk6Vav+0+3ADVMa8WREDP+1SOCfbjaNShKRwr/t7wXf1Y/uc/zsznclzgEMRQdeOAdnm
YcFctQ2NtiQIfKsgSVRI+viqbCJMc1zyxYKIPlCaLdffoWf3adpzPy0tBz/gQ2RI1Oi978VyoKmQ
wBZ7/kvi5hvCABWbnbwSr0gHCfiFCQW07P/WEJaLtkiuPwlGDCEmbdcyBg5s1XtymT2isc7DqhZB
li7pEXXTlCo+xPumzIdh9vvOSRA2UCng95U7Coq2ipFutAQFI1NrRnS+hH5x1NWMk1+6TQLPbLvp
bzZjAbx60muvMjJI2QBdf2jDFa7vWkEILBeDT0xEMUXH7H0Zsdvcp+o3BRU6b2M+NULrCQspJOIo
FVietVGgi94m4uhVkRLAbf1tVx/nRYeeszNlx0opiWF2idKEFXkLJF+QeZUkk5KTBIikBpc1yFMA
Tly+sR219PBauUH+E0m8ig+eIbxY1zcftYoxlzqlq3Rdxf/l+4K0C4OfYmJfFLPs2rkcxozmfSk5
EhL4PP+Mg99uU6bCMEaI5Aa3QKgSEME+E9q8YQP6//JDwNAWuANSsJfJSdsr7wnAm867VgOoO4Dd
PmcBXskLAMiv6Lfb2cwde8EZgcAhQI4cDV2qVgD/I7pym2OhDhqAQzRgFmVt7RJiRA2gOJqqcjLE
0E8RGZxl0LcdT9chsOGSjkjDwZllbjHAKtSWOUKmr2FwpmDIlTLDz2+AmR2jdufZl5meDrlZxQnf
dFknCjuMQXNsbhXPanfiEGZ3d6DdDelWaaGAZRMKpTjIx16tdG41ZVnhQqAF5D36lNyfZFHIMnJ9
iuGFUc1q4HtnQrKQAMfVq0TV0hhodlUvFFfpqH5DQ7V7VZPgE9nG4ZdE0Ww9I/z6pyWCdoCpQoOd
lD2AD9RPwlsIcfV8RXM8cQZmOKgZmGUntMlxgeDwe1spXVtnIqzBgv484PhWD13pjHtaIZ8FpRJm
pjNuR8r7oTDLGMRUjLoU4PEUHEmK+Qa+yywLkrKKW7YUMcTqDBM1lMw948LXGDNlje035jI37ckS
hPFIiYeNC+syXtpw1OADS+u1yKNhgGFT8vNsnimmqqbFWL0CIX8Mifuszu10Qh1tpwTOd79E6tIs
ECAsB+e0d/av1F0Tve5EPAWIQ/yWgb2ciUva+qPSP7hM2DMEUH85ygOTdZDW6+pFz5wKEFVUNfZw
USSZSyM+PJrMbDu8Tsi7W2zfzyxNpPOpacKmsKNjStsfKUMNRCmpY5Yue9Qx2/rRv/Ku2YmQmDHg
75wB0EVIb/Y4awGu/+HJGDFn9qZPbYEbhLzX41bqQA8gM8ui8nH1a4pJvFFo4bMZf7pFR9rZi6Xc
06rZfbE1b0rAs5hByMt78cnTTwk3gW4/WFTvuxFor2ws5SAWl04rYhmAb7mGLQtjrE9erJ6IDEF5
JwrHB+ZYP5nKS7lNJ7TkBf1gm+ChE6RcE138g0iUiXS31RW+2i7x8tMmNgqEC2gQwHSTKIx6c+J2
wBF9JQXcdO44mSv2488uFuDb3fth0SU1b7LnPyy/tuKAGUMvSa99tJ+dekixLBtQg/IhgmvJQ9Fx
fUTsxPh0sPnV/nWYYX+rxVOCg2wr69HXO4q5AvB1jBbH0fYiB1SIoP1XHL+ZIbiwMN6hDYGPnXW+
mQT8RfrlSpzQit9BBsYj/J20wAY6HC/fQoMQcgY/DRlOjlbGWLzOpfJh+/7/Z0x0Fv7AW2hywOGL
2spm9Z9QmWPS3KaDlI2SbSzhqfE3dl7wzPNJSo//87GNcU3NAUmnpSBm6s1UfVLgGPqY0JbWEYrs
E8C621qiGgEqQQ6hgxsyItzFKhUYEn58Xnv0vcoUpXRDJeoB7qJ8rAYsil2xtaLT+IIr1UUXUNIl
oVsIYGcqBDxwYhFbJjbYAmAVWcwHzuIIHLpnTErQ7go6NIuGQy7jK8NCwLzC/e1+eU64nM9dvTN7
lvUuiGZBCERGzUIcTjrfT4NnqFGUgZD9hvYqSbiMIKM0M2L9pUsxLLo/SNhKhBsTThcQrnw7RxfF
il5FrkkxVofsmBEHBB6VatYWCs32X6mZawRI6F88qO5qip7vjIKa0YFThMnUx9H1zJHbrhxFkAz1
TGabaNcnjVlWsMQ9GGkKyQBXPifenRYeHM62vfjwWo5jc4Zx9EChEkitFU7Sj3gQZE2NvZij45sI
qk35IznJVmEaKR2ZZLdsHNgxBL3+4rw4PYg4Y5fkRSh3ptEqZZ5d3T4+wHvrkPYuY6O1aY+kn1Hl
SIOqAcERr0+gZjbv9J18uU7WqWbvW+cG1U+xVerKAOJfOjtU3KD9x0W/SuEJ6E+pPIrGkhHBTUSW
5O/dmqW7q6rUYTVmSqNcXTZ9sXgdpLjQ4QwSxoGjnCbkEfmB9LSFXldI4ecm+S5gdEAdavQ3DZwx
gHpTHTASRUA1tlZuCre/9GQ7niUMORI3qzJO6Wr3w8grpMQDisuKHmQvxdQE2Y1MdYGS7tz4USrR
lVn+okCSFewg3ers0WWbLphEUz+W7hV3j6/z9W20z4k5emwcBk0OR8uVppczuUJE52mLKPMz+a6o
4NDsStmhmfsUQT4l4wkqqx23WqZnnuqQI9fBJ4eRlFzEmyebPMoxpTdbZEibzvaYAPIUe07ZWiWi
PaN/KhgiCPtujycD1ATZCdRDvm5upkVx0ZrVkbb6W/flIbx/v1VJePjOS4BoDEhwkgsFQE/FHD9c
LZkGREKmQWGvRDVi+EHCUSk6Kh2CoyOvSCN1scoD3sC1hTKFPyIqp9DK2Y8A8cQVUMSHs/OQVeyG
ymdMqkUd3IiYpB7o6TEU2BX6qmgHnIVQeMj0RHRS8h/BpmPaJwo5vqtXXY66333LCxCXLqN5aVxt
bud0dZM+tTzJHKglwVnOr/XS5utXC7ogtqA0dbe9600XNAkinXPaCCiKqCUKRcG4YarbHBQDO24F
VG7+ii8a/m8amN9dFODC8uNS47BHX843247Y3Cz2i9k5ti75pu2ijP7WQmvU+dBO7uFWuVGskLJk
4xoexTxzkUCPCUkU8x5hxc+8sgKKVPgUqbHUZAbSYrcIHvX+UiZ59vUzhKB/N5eiCB6HZmQ7qrbm
Nr8uQAc+6oqtj2+waWR2xquSRkF2C5phacrAxpKLhYtgGLbAtyzRn+5nBmuRT6DzTpJwBi8qlHJO
N4kI0VohJbxhtkCyNlrdUwVxF+8O7zO6WTwBqUENRDevXHtOioJpqMBC2N7ARDpwWKbCHHMGKpzk
SDTpK/0GqWCbk5c7bvY0QK53eNIscbt0fBQegKNMjS/35nksQEPzgKQ16x/y0xI+4JeoMZjZWsMP
RXDvfkcK/7S3QHf8GxoSIesovTFHrXlfr3ozWFR0Kvo7UFlDCXUpnWNyYUCuCihkg4mBs4rFXKoH
MNu0WQ8kelfTu/9bYXdRh43owOG8MmX7lGS/hqxvvpRWoMMtMCX6dbMxQwhKs/QAJGz0vuYv0bgX
lj2zJNn7thVBKBwFTLUStlTf45iBzegeeBPUU0zlVa23ua/D5Cg6p4rRQa2wbqbZhh84kanBa22u
kNxYfx5kY/cMSFO5Q6qpnZ7YdbL3qper8SCwPp8qh2/TLaqycoahZV/Nsh3VZ7+DB4UwOVgmxunm
xShYL8bS7fgYRDQXNK6R2NgCMVctCXEnDbhHX84s/2TYjKf8xR/hFfY8KOkNTP/bVuFDN2XM8/6F
v1VjKJex5DHIyhftvJCFKds5pyok77uhmSuTZ8tzqOe4xvQs873lm/69YsVCqgDAfbjwcj5rv0NX
PyInh2vIT54pvrgWxujftEEgugMDQkvt9K1UbuDMIBjU94m2A7wHtfK5mvj+DnFMxAB5doWENcbh
oNt1L5QbhqXlRyp2lMHgVlIJKdWiily0aa0ZX4/+rQrUsU9WpjXZxnAXtoPGtz60LgKflvk6SOjN
AgjTkM/vwos0E3lk/zfq7pejFtzcZHtapQpfbD2yDewAUNXgtbYDwEyQ7IaIeQvix67zB5ldBEiB
qhjObt46nKVP11ShJUFAwjutICHwOz9Gic7niTCT1XCt3TWYt7oEcqcbaKLREosujLMwjPSfuEVW
xlP2GmQ5mQdNECdG1eZgSA5e+n9aCc564DLEM/qA2P2iYsVvKsnbZDWZl9Fo8VntM8pEGVyeAmmO
z7H8SW1AyGGFicGwOe8iBFnr0+uV3Zy8M+8+Zi0MCniCMR0zCTKuYAmLfp7kHjRXOEjbrpm4Qib+
9LKi32VAZ2fd1ZoNYh0960HQO9440b19owsLO/52/dfQeOdFo+a7N4/njfoSkCfyRLdZjnUPtkkf
Os07Rpn4bzpPVf6Xxc090A6Jz02knNvTp/JQFTJ9beH+EfvtnrgSSWoWn3u8JpcUK0yJz302xR1W
SE2Q6zsHt/+2+diLiY4dQzc6eYudFOMcQGuMk7FgvUv79Cw3aWkp1PBXz2DmQtOWQ5mmEkQYocS3
DGSHEXakRzWI2lUNrYzIcJc1Xlg4vNs5aNLDcyrDjtgTrUUS67aKh3cIWEGA1KzpYIgGgbBWM1Zj
U8Bofk1IFXxQF8ytY1WyHKXn/bhbuNBcHUUSdAqEEOCkGGWZoVezpX7A4Oron5pf/+g3aS1slv/f
A1OT4YGMG8fFitKpCh9GsC1QMgxDFk4++jLL2UduivSYT4nVJviYQjpusxlpW4vTcIwYnJdtv06L
ASNI2g4TX6cEyjU04/G2F7o4Kg/JDqPQ2XoLQwotGla529Sx/dD0tr16wy0UF7BGMKbf1juHlDOt
7C430wALAh9b8NMmCy5/EgD4cIGzvSdyX+2EBqqfzJx213RbqentBxEyEkFWe0U0as/h4oWXO/6B
Elm79QNOBG10jcI5BxSMHjuUbc1iD3wobV6osO2GY0d8lgau9qIQyEhDyShHAs+A/ro+V1BzTDbX
/2c/rvHr0A5VloyAymmeOT6hIB9neLXGTG3BBxXePgbCt7pWQIXyzCB5QMauNZzr/dkExnvOe9wV
RbN11+5DAnpRzkBxnEP3dwOwgXpATbPYVgNSfpgmTpVpUNE7DMJUWHM+aansHaz7tXVe+cGxqANk
4vcJTXeVXPapv6RyDUw0m77J5wjQbZvmQudy/Q4xXL1heGV79p0y1G25gjwCoHnRw1id9BTsPSfK
g7PRbzsbhP2Zs1uSMoRv6uI/YopLvYNF+I5qsY0UXNUdHnOCp29bfUssdrtdTpSosFcaTAmbd4bg
jySer3gsr+z/94B/rRMRaUtMRU2Oji0kbKcwssTgfU3nGl46pNxD5KvakWwo/ML8F1LEqV3pMUoa
PhLtthcAm2ImGpmB9vhoSRP0uM0jJpT0J4ST2mnaUe4rbpTfGw2p0bvjAaNu+cVPGw0hDmgOXa/J
GAqX72MRr8CN2mqpokOLD5pPuZ6stkit7ZTs62bJrgPi1YtZrbl87iIhqmIRM9JVa60fLB0eO4bV
PZ7tcH0VcmmpT/BaXYddGTJA3LyuO0BOeKIt0wPTh3lmU32UnDxpeZzvua+6FRmjbgnmBQniW2fO
azYUPqrw4PkN+nPc+cO6S5oM131S1p/7TemoIpzGLWh5WLDBBqPFkwMZovpOqND4512jhxNbrUSO
U1PWGZL9K+qitizL6STKPeWfZrb4/OISe5G09w4msE9FghEm6YolvaKyUwrY7rOFJa9bdw8p0YVc
5nxm0oxiRkwt8gy0/7SVnhOVV7sLHZIhv8dojORZdlY3P7HK9PhXwOpA8gFb6L8YwWNZwmsFdTCJ
tup9QlOH7Zv1KbbFk6y+9mTDldCtALmLjk0RqOmV0kETmRXNpNG6xnfoXq5o243nKxRdgg65ChBm
PkKW/6uVhgIBoWUnh/0hQZCuKkSyMotX0U0I7IBnAdtyOlT/De/HtCIgRlvd292QMgVZC5khSibq
50fOiJu6kOAaB8UE2VZu5BSXWJRFhDomiCumtbu0LJtu+jiVI8e7vTMCIEqIKGGTGQDby6XbjG0/
vcM3jIpEnDYF4FHL8t3hOBzQxEEDY69A26uXRSnz4OJfUio97OFvUvQNNOETQj5T/pP7dBlAJf9a
oOOxQlGJsCgmT5+taKlZejajH6/rAfY3gWxyhwogWrBjBHvPGTtN8N5NmwicSjcYfvRl88OG+Tak
brzB7qVlf5UvDWPPmBLbf8B3te++7frGtJabDv3U9x/HS6DAFD4yhvNHcdYH5g9BkrAEdyHO9oo8
bWwhMD/Gpr+yYk447E8tmJU84Hn5nUlYC8AisHK4tNyc8VbwcQbizEVG6w08flGw3osuo21F3qzA
OfTEOAc2phgj/l6CVSQgzpxzobirlxBq2KlQmERnppLgQYMQcVyS6Iy9SUSfEJ/WJziIFgu0Hp3n
/c3OJiAT0/tkhkhJSCtfgRBIY3cdnIUHYO2RbuZWQBm8nAc3av+/1yUOVikI4CjvKGLnJGVA47e9
5O72Kxicmhqd6MeKUHHsHmoYa/R1r6rgMVI4flUoMBHvjan64AiENYdeoRc3BktoH/gh/hKTms9A
fVZnEoKN+bunVbo1BHDSrl/x7UuVVkATxJ9iWbH36pkJh+/kSe148ApA/pV1nSRSRHQSsx0WLx1U
lahooWOzzww7uH2lpdX8LUrsdB2ONG0jpHhCWZyFS+4cB9Gr6xYd+/qhp5g8WnMEwq0ocp6TxgVL
1jyVFEcy3erq0goU+DU1VyU54m0yezMwCAu+z4h9LR+1DFvG/GnhRGuyKqDjWfCJcWJr/V0CuALk
tgYxHkCuca2heDJjYVIUoOoeRsSyEWBdhScgOB+0j0hqm6QsajwjbihI3DxW+hv0CGu/hClo9Pg7
VqTRQj6DrYHux4j3SloFQMFT6E7RHTzL6tOIW3ohPqDqjyqs1o4ig56IwjB/R0QnRa5lbP8kZZBK
bjaqlMq8ffoMJkImtrkSH7YnAOJmU29c8g0+8T8tf0/WvGWL0hBkM30HiB0YOOYPd4z7wSyHgDew
9+bkK7uYcTvw1IY9rpyYMVG+F2KV0pJXq7dUqrAh9c5bNRSHWsev9FHOJhlgngeR+pQlkkNmediL
ALQ8rCVkTT0FJwUIuIvZjMzWSnAvEB43G0UucfNK/rFhg4Oi0JxPNFJoLn9aQbMYT7IJq5yTBIK5
63YMrvjpScEMgtUV0sQsbrD5wNze+nsnN65zmh9mbcYgPzX+3XtKBJvh4TpF2vIXveekmkoWUUvz
WRoFBKsDtIIBGIeUs1vG7z+jhWpeeADEG94neCO2WZRHWXhfREkfV4cWB36JB4JEsJ4yl88Qi/J7
uzbebOHZlXDdGACYT6DuQj23qL95gq9Ri5lTxBrE5Q2mb0S/Ri9LX2fxiNfBuFh8QcUfF2Y0wj2U
WUGcjiEpeHLb/NJvb4yiBlvg2/yEhNlO3GD0o1smnc2xSoeAUiscdauhLyvVxTAeG3crnKvC83tw
pXeSv9DAOiDRlCVS2FrC4vz1F6pYZb9QLOl845ApzXz7JXSuo44IMtguSD5fo4O3qvo5a9WRS992
G25O5Iwta4QGN5jCDH0IWKT80d6kgzfEBKow+y5p+dPdgDgbbWJXWMAndNnkohZrAc7CgKuk8ZNz
PupwMYXVO7eQZHIp2YGvuLiphHGTG3+tboMvWDX2Hpa6CJhxLJZBsiZDZk9BEe6PAcOshIfDnbO1
b37x++TEC/FT+5eiC16vY7mGVSyra/C9bDG1gT3SrCNRq1atgBFYqM0PcjQTQuQPCnR8j0u2u3Y9
mLBlJIWvICm020xY7mwkGh9ln/UNy89GiBH19OCERXCjz9bmOrUCT7JvTsqGfkuGP6xY73EbeBnx
Ff2Af6dXnui42bBeNdBCiqR88UXzoLAT8VCTisZqPhXp7tLWxY/hfbQ4tgL7gCJruUABRDpSjsOz
JvNplIwmIe4YCcKICSTk5Bw/Wv5miezpAwHeDMaDxZ5eOR/6WSW86mzKPcn8z2WMzioWI1F7BzWz
qac137JQN+CF986b+zW01CiTBYCeD1uFjMXbtFBjY/sY7wONHRFjaWumgvR37ZH+pmM2PIxk4HGl
FfvZ88PRkcuLGS8fv2L8WjUDORvbzxYRyFM/M96cN9qWD+KyqxweMV1qKay3rF76uOC+PCicd1PE
UET6rrZdtPZAHtxaNmkIZxTh68mtfj4M4hZdIGWDdbeR1bmvBiquzZNhm0Ff29NMRGL2tKbq6SXS
jY3XR9XTV9OwsbHtpfm7B/y+/wzZb5kCe8owMfuAI3G403eXztxElrZHyjfcoQmZOndgCidMZB/D
CD4zoRbywGJA2erU0eMA7WGejkoNn6dizRYPmi4t6Rc2Q2ccprWkoH//qHIKvTa6BzyHulA06Zao
pyT24ZAYhqlzZk3kLEwYcEz1hZcsTtu6lBL/RBLkzy13dt1R0FC2u1C+WxOWz2iL9+RNSvh+JKpR
Qam1U1oCd9ViivZFq6+SG2of8fEW399FEZiGKrAIfltMO15Mea7uvWiHbSeSA/+3AcC+VDVbRC+s
DakqA73lXUYF3WqFkuLKl4fqMElsTF666SRe74F56LLrnmbFuPNo0jywdv+sNHTUkiYudA16bcwc
cvjfS3pmcTf0sc7JPv2czBMh/hFQc6gY/jd5WZHJ+5u9nzELsku+ix0GqPRRIZ78+4cZqR/543/c
oZNR5NL7Y73E1g3C6EhX1P0KQC9RrTwxek0ENc9ehOqkWoS59WXPHvZrV7loX6VE0lw5pZOa86sB
RwFA+XsBF0AIxdwRE4Pgnp9dJ1T5U440Fgn3tbnOfG85gLcTX2Nuy78DOA4dYojEFI/Emw8wux9M
P5Dju7Pqk/EZS7BibwfzHGAtmpGAypmixQqVVrVh4xdBzPWSyLCjuun6H/cnTmTByEniJ8H3cbiH
1Rjv10a1JzhAEGxERkxtDKQw8fKQ9eG2yzWsuWxtQh61m1ZMitKmeg5zGplqErzMtdpLdp9JpOGv
MdKbXw7GxiBN7d2LCio/E2pEYkFfGmleb0jZjWjF1IvvkCarMZPZBEiXZdiv+Tq/LRKP2XSSiJMn
LcaFJqQUhMbNXAWeK8Ptw+0pax5oCQ2T2K9LaDOVOSTy9RWUwye1E8PTv4YyBzQW82abRB9QbI2r
ICzgx+xgbNPXFiWTJAy+J+gBiPC835QAn19VPPRLqn2GwTE+UErGDf4QvHvMpRDHxuNJrTKUpimB
xU+C2ZI1nWARS0nsx/RMjsOtbJmAmsTgtV4zhb8h7Wr3VoJfop5s/lzA1SlUuNNxgTkfJNvcHxhp
OIlVeN01LRPv/vaxd3sNhZekOdXHPKBYfz9VIvfKJ4oeoJAcnKh9mJsOGdWjb4oMSlN5qsKW1znD
ieL+Ra+mwKLTDbgjR0LRNg6dlfmvauh6qy7UdHdPY+suOxiDnf7r+4PM1SZJQKZeDARXZf+bdT0s
wO6WU6jrqoh8RLM2ILKJ2b9h7thqDuAunJSnJCp994GYBTj0kDOn+5Xg3Kj6hHKDpbOaczEH93hR
9pAV0Dct0nNUh4VTP1rAHxlC70dz4HUf0iMidt43xxY+uIcYdkMTGDvHrkJfUbG+wv4uNe3C3o9S
rezg1w7rqYGfYuyO0Cy/l6lS1MJcFF2gZzroihf4SlT5Ff8Oce7vobt/29rD4HbhGFIkjewTjV3B
2gqCshou0etqnOUb4RQmB1peagd0Z0ncUrqO9Ecc+yYLdGu/dtz5fogKb5A1LAz3tUCWUGHbygmT
0Z8wLrnHDbX6qb3MGjnZcsbD9/qlqydgcDqnJKgHGqkrb3OSuuaEHYmC14+pU0hlDj+r9yq9AnOF
7tCa6V0p+QKHzhKRJTehufu4vPNOh0sulJUuY5W/R9MXvgk304g6gwYhnU+gr/NqIR0KzYxOJS/v
GoSzONgfgyhkljIBkHKxiCxlnJXRPSnuE1QaJbaDF/LyvfZQ9gCaO3yNR5MSVKfVI3Xd6EhqEP6p
lEP2KcgD14c8nMRcWa9hQwPeGC+VwxXgsw4Fqnb2esK1rBKCjdWSBRXYqOvWMChxoemJqrPbohPC
p83ksMyB+KLH+ItuLFd9MMivRqu11cae+0M7bs6ZGadMmYoMhvAURPF81IoE/aPW/a+vRAr+JbGW
vYrRSDwYhi7e+tvRuehCQZeKscg+IPcvLQlLulQtrKiy20/hWdeRJuKXTm5pQnUlVIXJ6nkIgQWP
fP2oYq7TVItInB8c+QC82+kXfPPfrHOXz5MffvtkVYE3J/UCjXh1O8ZTKeYHy8TsnQLBtfsCREbG
1hKP3vwKKs/YLNYblOF3Xbx7HivCmo6va720Zt+8v67EajZLFZWgETR/w5wouWIcJir4Kxz+nOae
D39k3Lvzzq6eAdRucc6KcMPxYMRIgH0eWm0DKByZ1MUtcUVNXPMPm//BOYn+FQSsGlUKI4h7094i
7f6paIwpAQU24LBINut6EHu4kXQZLzUSgmjY4Io3EXU8Aceco2oW88d6yF2P9sEvgqvF2QKVOLUk
JEUMo+CzZw6xruDV+8MC46DbxV/jS3vBE1kWanehiL99FKuajf3ytxn7dYvFliOLQbYljGcaAMe2
Hpvv4wdLQ9Z0Ot8pAU7LTYNlP/Fop6QySL+DMQXExuFcEBnKvXQrE+Wo6nxwKtqtf6W8fPApA/Xz
c1yu3or/dcGZ2oiRPJOPGdkCnWVI9AW2pJLKVNuDuwkh42e+aP0y8KpD7gDNczrtnD1BUO2XOVzq
sE/pLYU/u4Q6H/yLKlTvDoz4plHY5lu1Eig6HLD12tVTTJjhFG55K6ZxxpGERKxhXQkzVwt21s4L
LQfUKWVFHkwdEy38m3SWLkPRAqrTiApCpmyV7Q6Dqwlem8Q+OA2SvruR5dmcALllWXPqZWV6/a+W
cTodGNWJtDzFksHVhvtho0vHwHG2LTA7sUR0k+KIhyexHehJ+TEEzhsGAEvgiCjxeGbD7FgcsDKQ
wmGV4HtX7bjzCyf0q7cTDLDNjwCvivFMByjDwLhyAHxcGHXV+Ztzsmw1U4Z5k7uRcVxLko9JOapw
bkplOu6uxT5+K+aq+rRFr/pbgLp1KsQ3XytBR25ai2sFrXaLNSZWS/p+7/73RKl4bl8UL/knIw7G
0kAe7EZOZWCMGhr2rLPeJT8wcTk/zIO5qzEj0sT7AbOHf2Ojr0OjLcjERIMkbRyvy8lXJ6sI7CND
W217dgrZIsKphtn29Hr8Cx4Yv+CLeOXGOo2Aww/VockKlP6yCl9cCgjs/dbGcFiKxrGiOarzKCuM
q8oi7lNErCWSn11sg59jIZg1kMjht0k9fRbsPQrlVqvrkk820+80CiyxzX/iqk08Mk5Wfjk4TnFO
CRwtJi8KkDBM2L/bU48a+QybZ+xUZdTRcGITz2hVYK9WtHRQZxtqi8THcfuwSBlt5a4WpQgANSXA
1rtPrxP5UledVEJVhdqSla1mm0BLCOsokctsoYZtpDvcZJXrxjH+x0GjRSwhGk2mFFSKoAeArMvn
/xXs/rvEfrHN9KoZfCa/Rp5IJXaj3REkMehLaPIg8TDiAVUCAvM+cbw4n2RjEgMg8FAFAmg+6WI/
S2PhqC0tVddZ19Q7o0dI4OClbGqtSkFx4f1CG6Y32QNfSFhNdL1uBz+3vGpT2YIrhzIyrDHTMGai
zXTUj5PEhhynnLCwTo5SaJT3s6DREqAoQeXtqG4QeOBrdAoL76l96ROpZoNE1siSkJ0ITkTmbnTZ
eV0jvp2sl3opL+N/wuOUfJ39IeyFII7sTBaGaImBpo7acppUybaTeIaufYPCsGyHsOg0cXtc+j0X
0QziP6lbSNWclRbh1FuhqKvk18HkwDCdjzk2cmiSnBNRSrA0Qk17X8e6vA16LTYmT3dA4o4+GwV+
EEGqIJ6nVY2GMih2umXwF7C/WKixYNIFydEyUmWepR0tUv1xR8kuK9qixzkXgu3ii2JYpYWjh1Xj
OFgvRDlbVfn9rYn5ZjJkNpCDo3C3Vq6DKKXi3RTKFNzFhfWQVPKRnAOCcO792WRdtS7isqtPlLEI
227HT13qEju6bPUgD8oaegOYsVObGbiV7uKK7O6sHJi/MkI2Fc12hWk7/OPOlP5nsXFGK9zKRoO4
Z6pHTCubxhd0h5wSuRyAbA2wZ5NlrQIdZx0JCATBbK3XbeGvGkSafWRnOM3KPcVOin50sIuoTwZB
ilVSJA4WNT7EkvDUxNpRPl4uwownJEl2v6cqSGglhEjYXWN45vQdX+IKubd+cHpkBbBTS5xShxFe
EomxHFdICqrl2agw6JM1Nn7sgopJJGdpX8JqxyYBSxngc1pvtAcC2PoiJZwnwQobzroRghDKfsr4
knYNUbznKeQPDH5xnQBHnpXQ0rV5k1cCYUFvYGpBIKrLcm8YdGqRpwSKVbZ2THWqAVCPIdMIRSX5
kS6lr4XKx+H6d3l9D60+1pAJbRhMf7xuwd/TqZ9GycO0vzzI448Ok4i62mNYhJkt2zzeiu0u/hqx
a+7vdURt76vCpoGrAuONiNjW11pbnz/NUvY52Nb528vLF/zJZuxvORArrbJyRhcyaE973KyK3blt
sag6k+V8Cb8xdy+gjr28pPfisIH6eIFiPDTD47zuoyw6usm34ROzLvEDIsLK/x/kVugBefoRq1qX
PbaBlOyfrYqC2LOGne+32oyLEP3elOoJQ9kbJjqxEh/ucRzUBVdsuyREYyFgFYuF6r5FburkLLcX
D7dg/aADrrSWk/H2oJADTeO/OIcinWW0xXEtVmVkT7fn20kxw90VhE4JYj6Jcx+H25LjdpgwdMJI
pDwNeZP0LNtbiIP1mV/41Y7LLJ22sVu2eo5mR9Dg4M/O8nx6/AegLHq9stg6doNUc8p38Twopeiu
g8yz14ZXlRPg6EwFohdBBo5yoPWlAMj2tJTV43+jHcGSNvbIHbAyndgB4AsiT14qn7whhodQaFNa
bpf0w/ICmCA6rrxZY8Sxa/AyyEPmp24nSJN4T8CyFqi52hRgpj57dE3CGfyR8y1TcUu1wgiF9ppz
CyVXC5nB7dk039Y5RS6bI2Va7sU0Rt1G7rWFz6pNGdJboCLv2LoO0kf7ykWzXj6bWBQGnR53lXt+
cOvG9cQ5WQpk2xe+ICILRHIR8b2B+UMubv2/Lx924a6MW4AaIlEsV33oOw0q3M8r3LfdclFh3Nmj
tjWY4n52hyn52xG8SLnnqoNmq1ouGKefXIBiiJeXFlrGhnKe0pO05FpYS1gPrUNcR1aHeiv3WavG
AGutBNwqVBAjlvrAvJoFSwsHXmhSm1aiO5wd+AyveXF1Fc9EzQdXd2bYuXyD/2IU9otWlXQfzM5d
jtkWrMKWoVfj8Esu5OA0CZKIfJJjo2YtbbtRPlYcDibyNai7YEN82ee764trSPr4t4V2KxTKwfPq
e8PNpM90gbBZVUD0mhK7DSTur9xoOhxrtZOb9TEaHjgASo1s1x4S120SwCdlacEnUMXenhTrtBAt
K6RJJrPe45tBG4VpuYrfVuKH4Zqq8XEFp5GkB24YHAI+UpEKokNFsgf1Z2YZmIZ/rs4QkUt+9pc2
PZdiEnQaW4fS6IexZu8imJjcbjQGeYU3xD84SSMb+NaLdXwBf+X1F4kVUG1nVEu7G/sEqS+/bM3V
z7zKSVZlBZ83qIPMhVsAMo8KUAwFPvYimPryqQbLMpOqGUw21aYTtYoMNB+PGFhLTOVqx9HesxiK
KSVIuFG6CLonpMItJwouDWrJUA7H1pW0TLEQ7aPCBR2cUSOxV5J6aBK2HL5T1ZqcxErZAnzBdvrc
nSgoFOFCTx6rtLftzsgbFnpw5tKtjaV3RtT8AItTQx4mDqLDph86O5w1JunXa9QDl3t2UOSvmeoL
GBMqCs0gr2aqiVOauvvufWLFDCHFBCI4hQh3fz6gF51JoU0cct+AqbgJEezhgCVt0/mIMwFm5F82
hdLxU4rMCf2HCzs4LqmYbDmIuBnPx586Ni3shNFfuf+RCGcNC89yDVhw/Yn3oxupvnh/6EQgD2Fq
iwh5MDdCHgJ+rTDIw7Pz6ZFZGtsWQETq6yUs3IM9yLUCneq/pWv6NZwD2eh1x7XwsCiH8MZ0HJSh
r8Yu0QkDHl1WIpcZz9jmPBuK0ulj9nN6x+9Jr3Ii6CjAIk/ZRDC0Sd/7iXWIrnFIjmcWClx8WpJP
m5xncWUWdIgH5rQw0vp41UPqTTOopWswDg/dgvZDI+jDW8iIChV3gKDcE+EZv8LESRzeq0iKVL1m
pp6jouCZ8Yk9utXgKo1va4AjsCzQX02y0eok/HUZx4fnYzl0Mm8lyiIskJzuu/IK01icQL0Er1Kr
iL+OUEXAXZ6/GvaX6jauvpV09lcMUpn9Cv7PlLkQ7xZ1zEyH7EDYnvoB4zgXCVcTa20IRl4LxyfQ
CGcscxIaz6OByCMEo5LWnFq7DJ8wqCvYtGW/jDrMTpVrW4VLewdcVcLTjcuhOg6x72KJ+3rVxAD/
KBGN6lve5/+VxoUzbBwfPKAJyJ726cjVacFId/6iEhptMu0Wj9Uz3unt7sKdmAuvSBHk7ZFvzLzg
hb6mpPi6reMrf5IuW/sL4xoGsUUEKvsBXeQLk15DVNCM2/jJ3Xzqouptai0P2bLl49+pauvulngt
Y/WYudWu1KMHfWoBSlLAlAdK0RBfNu3Dazbnu4Yl8kUdLDnxtifjO3WrGz/oMVIw0m1YiOHoIrVN
3dh6+z1pMnJ/Bbea04R4bekTm5sQaDIA3nCrsEba3AHj+pSjecagRposgi60Bq2l3d++5mDWBVm1
S+++cSCuc6wRZelENqmH3xz23+hmYkrIMxRduRlyWwx35OBCn9Z9XrOU4cZuXkybFaZOs6CengKf
wZoiJJHO0azs0fB+s2fR9ZyoEnzyUFzH7r3YAbpcuF6WcAc37gRZkf7RNGMf+e0NSLuTM77GLeDG
PadzRifXZWJxlc7XVwF3IivU9Hzovq66Jw/IFrj4klW/aBldq207FtSlNb8xj+oNQ/DsKKpAjrFW
jUCgH8M0wF4zQZ2G4vFKZqtE1h873VBiGV+LhsDHNXjj1Ppc5S2WTJZmJ/oT34LCo8wHybnfP9Ly
+x8zJlIquMSehZNhQvp6pwn1s+mM5Uy9xNY9oVaPFXj4Dj+AlZyJEhgKVArQvRoSIdYZyjJ8xBn8
cOstBi6QSY8u+SS2WVLt8YfD51WBVoMYwq79PBjV87VAR9ETCgbS5R6nE9Tmd+5bvmVXKAMc8uuD
FIQz+G9MjRbUgiKT/J9EL/a8I96NQU3Jdh+kXv58W2/0ozvKtIp5NKG5qq37gtUzEylZNt9PCBRz
8EkAYDmqVi4e2vi+c1KSWwy8JQNn5rFqyu0hNVvQC/t9jgv2q7lHWpHimTDQMm0Y7GpTmHHZMahr
tJyIJndeLKDMyT9C4X6a/+bc0CSoP3Qo+S/0s5CNaLN4AjEDPZ62CYCSDJYn63KzYf0E1D9VKqeo
VkrDmdF5E1oSFdOfOjIDTDRlxs6Ll8dRsvrtxcZNNlSnTxYeU8otjLHneDURKWhRLJRmhT4tplhz
bbrO+jQEhbNnMbiiqGAc51ATrsoXqKTWG4LiNula+gjphAT7cMxfdqWcffL1UZLV7rUfUbVSTeJM
WzKzbi7DI8kyppXe3DPJ8z/vsoC+xRTJy+qZ3tZhPIsar6zP2GY8Njiwc7nPunweTx+58S+bOjHE
8M4dP9p2pfN7CYLXhs0rBoZfHpX7G/6Aq6QH0PkPjSOsh+cW5P4uNx9S6pnfXbzBcgIa6Tilo5ZS
kZxAEv9CJuvM5z6fYFAbA5UJd+iHvYvBePcKVHBA/6/QCmDOXHOPFKTZBFdkomz0Zi9jJ2cDz3S5
O1oINx1ilrqkVap3N8Mh0dse2SOlTB5OKMw1Sg9nZfpyfcWt+XtztO/no4X7RAaSKLV5JYWsZR3D
DE0wzb/vaKQhVZjYajnHVNegZDUTFbr8Uc9WjbFcV7giU8Rn8ZTfB/27JsAb4mJdkA8wY9beEPWs
ic0bT09lknbLdQKL8Pkvahb2S3ORbX8yWK9kGKZU03KdQROFYFF8hQzEzi8K89aC9Kmi1nz2ddSo
Wi5ZLeMdndIR2EKA6RSXxKGf+36VRGc9t8TmyRLmvpwTOpFj3a5Ib3Sbms6S9C3GLbaPyL35rlGX
9Aa+Gd61OqzDDptR1lsanRaNslxedmYZIaD9XfONmlSxlaJASHr8PVFxEcbVaXH6EhCvStINDwDO
YfoRPK1gHanczktJC9BXw35Wa5HjaImzJy+2uPN/9S/VJ2slaKKXJTJpd7uvwWn73/lMSfQF+dJS
zOOn2IOvESSTjF3fkW+3tt33rrBz0+Pj527h5qx+7kCJpNa/D4rDWUGlI1PWULEfO356s9E7T8dr
ts9K7y3djqgx74DmN0HT3OlqeIbNnOcSb9I1ZH74YA0H7yJWNhVRga+L25H7aJFAxLIbwwd+RU2l
WVUfdonr4gL9CyzzQPIikSHVC704WvOgFw9Ly/9Ck3wXllu0yYEI6rEFBvoEHDA0+S8bJDlc493X
/yhfgay3cezp9qB70mOa8lWQKsrhVOtpP9V7621mMWqHaw7D81MocG40I3KIFET2Uc2PLszomlFx
DeS+kmg/eguhz4elRUoLtmKT2H/8ElaDjYUdcXOR4RzB8qyS/HvtErv4UIWsYc3njHJr0uWQIdAA
w6ipSPa/SUDKeobsNDizf5XQ5+7fr3dPRIIN1wAWoH3X37AGKNzThV9IxOSf1e+FJEo0+wd/oBj8
gQ46E4MxWwsblQ123iDONVgdVTodUtfasXSF+MaSec8/0khcAFH3iCYLH+Dv4ZbVL/EDOA14FUAe
7MOU6BikAQsuB7x7torEA0xPC5+sMDjUqVFeDqddlNhoSo6d9iYlDx5GR+wQjPr3XZZar60fSdUE
P0OTYsgtJvuPHOHhhatUDyuN4acbJBeoeg78+HL+u8IBwW8UWEs7zXyW+UFoATIdIr2N1UI8AH10
1XTqkgS4vL9jPtssJMrcZGxobSAds7DQDqa8dHEMuyuPQnKw8zPJc5iB332omAi5MCgbDx3Xmae3
PLEkF+3971QVeoi5MB+k8BvCMgJveu6O8GfSsv1ZiBl16LA24DSHSv3ehNr4vUAYDp768Ausuq6M
xGB1/yFFFQRGU1z59hf2d+A4Q+Fms/6AmrrRkqZMwDSVSPY8INcWeIr5eVwyinnKPbGfzUIPUhm2
ejFSee0Z+ABHY5cYb80mCkXnzWINoZsd6Ymfumq75SQsmjBDl0iKWI5epknPGl1uynkvP+xl3pcr
Y5Nuc2uDT6UIWZEeVVmgoRtQFqwIkm2augKfAmSZmR/qd8bqQxB5Nb/cFL+atjYtpOhMWYO4oW4g
PVfZh169cacrT1hJnfBYVH4Vk5WO4vTHvKJ4C/7meCwX7jBbdam8CNe5pvhL5qnsi0OmZkwAuXzK
NaZkzDKmXwkh+Kzb1142Sf+sLWUqghQ3txU5BPzFxhPMPhVtiSqtuX6rrsR8DpYD94A1AjaYy3YT
diRrSBRuPkcCjgPUXUxkfkT8u4TLF4C2wPpFXl60KhYCugLUOXPrI5AJl5jHu32kVaWQznybRcp0
4sf2v1Ze2GsKWbJKjelKvRGQzv3qtHTKVqF8zr+5vYnp5XbkajfinIwxeo1UVz5wFxTm022pAMeR
QY/5jK9J4XeEansRTK149ZjqmJYeR34eezaaKRnJEOrVaR+btJh25Siz2bo4PWlwHZanztG4UOT/
HIE6HFdeJSIrQr1r/a3bPetba2AdZ0HZjPvkoe4ruHDVK8swFuu60Mc0ugd7KZUTKCWyn8M6VRHK
10VdqImwP6ONdCF3T6JhoDosF3t6oOH8ivZeJg/SKwPMLKbLqDUdGOZJxTEXyXgYaaLWgRGljQpV
QYGAR8DknD1hdNQ5hkK0FE4eL5JHd4Ar+b2tMLfEoXiJDpwyXLrJ4YjWPDqn7a5QbjLfYXvAOtgN
YqvbjD8SLzCMpv6M9oppGQJxGsgcV7DtQ5D+Lh8lnz8iJ1orJIJmnfIFsOiO+hADzMtw1SWreuue
633KG25iHRyNc3ARIprULwOgV4vJ6r7xzxLuKf2Btgj3z6g6lURT85RpDWic2tnTYA9JgnXVuSUX
XkOyQIhR6qwhlP+1gXlD3G9rycm/VTM/31zNrTDrlnCY6hRBriTDRcGXPFc/Rza0EsBpp4Mm77Vw
drWyM4rUNdv88f3kdAiieQj5i8V1q2bATo+MD0K9jEHZ+tOBkGdJHxgEM9ZAGvRkFhpB26b5pX9s
byA5631md/hPY7snUm5f5Z4RVWcRtrGBJc/FuXbHoLXuCVsbzNcKZiqzKZhhl0yqTiOUdWXQuV3O
2LSQoL6JaNrmTPDA3YBznCclAaEK114HBcJnNNTgQEXHKFkh+6BcLmTUoJVDEYoS6p9SrfErByAH
6B3/spbI5z6+OANOs/wIQBWzrxRpQJdKuaSvpZubhOK90I0CYF8dIcWRZtQynhmeQW5bMu3dcDLm
4UwqFW4viIJoMhV2dGPU9i4S6ODyotrh3u//tB4eRpFLD4xAyM1TfEJQg99wHZmBMxKvOZPE2v5J
bwaglKYIK7HWBoJHXwr5o11nE6D2Rh7YEt8zAkoWVcJBjfgHcEIApzY18U7IQ91CwjP56Ebaa0Cd
AvHKhKddEyvOsXYtCdOFoDTlZ+xjEnck9liAyxFhd4/nL4Ij7xQHU7YwSrX4L5V3VbLH0FASY7mK
HIfATj5f2U/FG2v4NhdCpUwBnXdaD4yMy9+UYuMPagF5NSvkGQwJ/moSt9Wy1OM8QneYmYtNHb1S
C4eMizqXDHsyDmhX+ET0vpZKdnxsIOfYCndtLLhbXobbN4U44f89tsAjrC8QQvJwWA06rDVcmbsD
ogkX/SHwA3LlgZTbwiRWhJ4J0ZFp7AC5164OUOLGEOlA9XhZ7p96SEQR1NmlrAUI7uPxA2s1acy5
/yx/Fw32lqy1aE2pLYfkQdBc7iIa6JHc+i5tiTt8t8uas1hPKmIZrWHxAcYZgubN7v1Tmc3lsw/F
aiw4Uo52TCcWtp18/plo3+juJLahFx7pRPZ5Np/q1tOA3sCEHQL2q1PVbhwRJa0yqI6pDzyMhvPd
Ii+5D6PJsFpOqz0SH+Ur4ehX+8ecsFHicCjM4Ftps8Y7wrqjgvM/1Raz7ZjL9j9qRNGFmWVyN/q0
Q1YHZheLG8/u5xAy3+TkUrNSuBtxzKiaR3AEn4VQ9VE3mz3H8QIBh7ELtZcTsbXfZu3Acm7YP8IR
k5dZtZvC+S70Kmo+k8neCtOyqpzZLiX6800mvFL97/FhF2DcG5VO2fTs99EKTt89ghc2frOsB7+M
Wc8f5mrEovhdkD/k1yZiSKDQHQOX3CAAUi9fmShxYc6sYHaRrjSf5bG85mFjLYHRR25BxBUTHx3S
XvmflCMsWVAw9oV5W1qQ+MatTfQl/fNVRxPdXFVc1odSKLLDiRozmejRU7x5Hn4wLrdpX8JYezPc
FGZzceofdttRQitvD0HlKOS8ZFMQFXG17VCIzWlngmi2+r5qBJFgUpz5gXILcGOe7dbqwYxh0+cX
tvKI5YTBZimqOzhhtqQzEXr4L2v5bxoPXMNo84XNqZtf40PjNDMTDF18GRtOdCKbzHfkxlU41bgv
6673N0c8hR7ojX/cqh45eZoAZgzfoC7u+DO3HWj2s32QE2JkCprMxWYPrlz06InDgHYe0PUPYchu
pavQhPk4C4Fu5351W5KQu+UZD4oETX0cm9E0buqdSwIfU0h+bTPves9HdPR43sd4KiecXq5XzFZc
rHKxx7+t+GMquzrPrcNWcgMWJA23XUI26rEHiysHQ/pA3u0+HVD2OLJPKmdGhEG24ipjqOXwrDfP
QnmPxq2Mhe5YkFTgfZcR9cDhyQXZQn+u0OYVUyl2ZZ65tr6SLLE/ZOweYVCHz/HSIvmYw6/f2XeX
ztd1wC1yua8HQxtJThhtRSoAKTtD206uoRTVLjPfEYjp9oiUwWiZ/eB2lI0HV6YXSIscbapHEvXI
vKw69xSavGovE/qmgxDeBf7JiHoh1AdFsRf6tozOBrE79sVI4I4WjAgU1SFdDYHuC7fu98QYS6qj
mydrwMxvuJRWxEaIySHEmDR8KrbzXC9xJl70JNQy8pZ9uMMNREDmHSLljOzXI4LrpDdDBMR65kYL
bIDwMiSmsuVkcTKYVFbtN/6nPRr6X2F4eiMJ3uTfAIltNyYJ+hu/1w1DTYZGRqRIvFuI2ZACSyhR
Y65pj+XIuXfWJcJ5L9g74NxYeGSRbM1O3XBgrytkuC9Esoj3C5AWBkJabwyhsArnQJxDZuCSODE8
TXMefvXWAVoF/1GGd8TifzVGHNNV4cA2KHjKvbfHUZAw6GwXNRB77tWPtm1jpOw0PzYT/hdMIVwt
6m05a0EONz+p+AmWj6yurjqT3ZWtd+0dL7vOs6lOJtGJF9C5bclv0Kbk6YNs+FjzIjPgAtziytcj
xODzlGzU5+k6HCRANZYiWfJWoH7X1wVfOF0Y99dnrdF3pgPpQT1g2I1sElXthksvVtplk7XyCXAG
s4MFqVwC/+AXeRu+eRohWo30RRqVZFhhRmKVDvWW9NJ2y3v0ya5Pllnencf23A9v69F4tUxn6enK
K49FREoeV3ipy2RrWvgjb1UwMddSJuugNfA4/bzajZUe21Cpd3nROohFJSV0fV1mJZNH55tRGsHh
Zaxa4pMcWdR+W8HdFZ3Tp7wjMvCbtDycqZROV+fHJ9X1pLTrangEaYaC7DI+TJnWslrqaqyNhyKe
yDuUEFmUp2WpS1kC4r/jxN34uxro5eNgbjhgHE+J+kwfCj1SU4jYZPnXMh8O65Y7IhwJe1ufG/8p
Sp1Ro1DBuECbvEYPCJALUfmSSSFmkYy3P/QBe6Ub2B/mp96r00fvgVVEHkqbnrYStl6yOr4hHvJg
T72aY5TzaT7aBsfKM5vVZ5QfliCbVeHBjQ2V3eNT/5XHwUSFLeyWAXfmzGIxsRJv9tEckgprZrWO
ouwCGvjbyk96ajmZyyZ/8siPBjDrJwOtE8nfyr1l0hD4/aGlJshtOQU7235Jh7ZKEip36AO5Y+od
EXmARU2NX3cAPSTD6RJjNZRVgrbpK4NDi4Yff211pC1haZnFRYmUXUO4tZAeCYBqhTZ0diNiLQBh
EqeKsapu5BQ1wnd9tmRSR+EgH9EvE8q8oLTHrPAfL27Eh51Vr46pej+I4AH0GU/8X/NappGRMrCa
TVRqrvZpC/MUhz9T+7btTLnrF42363s0JbgDvWzNnDQkrp3yJWGfajvuAjAjtiLvWs/D2rjXIn9r
IpZu3Of1h/ilWVzrWGEn4p+U4AspDOIG0qNqdHqK5pTpW/W68wgXeGXvK0ua1vwBlMBfYZ6yLEs+
AKTHM6bFqCUu4Z6CMGQklucqAyQDgxLziKwym6iObBOJYp1DKfIQ44l1Jb+TOTmU7gMgr9DMMq1s
108TXbrezJfG+Fc/qhNxmQOh4gLkCrjLSJjZ7pDT5SJtnmLuz+XQ4u52vKeDfbAwDuB3z1DR6DYB
Xeni9dc8IK+sXtDvY5lE+O4xIgFEpngRzQOnoko695G/sMKckva8IWJoWQu3VNz3msUfJuQYrdOO
ySvSNtt9sFGe0J0GftoQZ2koBHZO5Eb8HPzIohph4wafvOIofH7vVNI3WQsBCv7DygqKIhZiJdPd
ektnUQy4QfNtEdi5m48m/LH237seplPwZSXDnLBTwAV1DUaagXhcKQxb3Bqgj9Hit4RNHnxcK7RD
xyLHDuXR2SeVOtiM+HdRn7KpHdB+MF9IbefpgDoQrSoBe+Pun2TcTibc1Hbe956PXsuFB5zdpB3S
uiUc0IXPb58zKhE4iCF3uj3aJ3ZAblGWLRiOdzzH2XT2x2KbzcdRWvK9yo92ldFp2ysbr4eO+V2O
GmLs+3rmX6Cmea4j65hi9Sk4ZccxiI0w7TMtrDl0euRHW5UaDoCmQhmXUsMG6yzAkLCD0XveA9Wn
Z70rZupcnZxAsePzc7bZom12+GM7ZwMRfD15OFsZY65y+ImGFFmo2RkgNcjFj8AhLlgQvfANaP9e
caYbCIFlHYHjM5QqoANVuWQxPqN5fPZiCXSVgXuP7NjBpalgdJnxHBw1VLQbowknRvSsbVZAlmZS
0QnGB9Y83EYVwG8jShutaEAIPOALhJFAD30XkN9yc034kMvItk5m7rbXjJ2z5iyVLEBNzPAEm2MA
MXmz/8NDJ9VK576uT0aWYlLiAktPKXiVJ1l4wrFlOK4SFv3K2kGmU/j7JQuq1BjicqK4Wpk14zhr
Z+baxzKI9kfmTlatRt3jFdsFNhr41NPsvR5BtkNAKaRLIdmeQAniQOxNtFnx0KXl6gt6WLwz2or0
2BOnXBV1DKkcBphf+u3UArj17W1qS+wxlGOuOavw59eSzJYRu7bwzzmDQ+GqTh52Q1KZTeyr/1ZV
REHi60VWcbraun9CL2NnoUWD3cGt7zzKYSWpeWU30ZMQt35pusYMAInn5vTr0LuvjJomFal718z4
FjWnp4Lw44xkLyS0WUtlhgolD56w8z61BRDKqZimwdovdwFAklsq+MAqeMQx36QOCP7v2wj/hyMo
kkJ/HyUrAdX7QS5kSC3VTeBp1+WhQ6uPw09T3jdCOuioFWbQL0ubslBW6uo3eBIK6rxFt/RKOgPJ
ro1KVJcJeheeZAfMOChMXcA4RAHM6trk1uupmrRCVkSugC1Y7mIWqrNc/JRFePdw6IScvH5AYp+l
oRWs5aXTZ82zXCPJk82FyDno3jPVbFi7I5tRYrpxt18hcwM+sDny/Zf1gLEULnt9Zqe+jMmSd3kw
n3e7ReGJbK6pkzNa6d3URi9SoWMg+DezSnX3MHB7Z9LoMYLeDuN6h8xcta4bxBkMMHhbh8zru4a5
xXzmmTV419yVBIusEYyNxlfwD7PKoONoUmw1JE2kGaL8o6Eo7ytorwpaXZR/nd9atxVi+pA+vGTr
70RDx6QPkQNOOYzaYVREN0AXwssbrVz51wtMoqDSUWW2/0q16/WavQ8SVs0MaXD4oY3zv2rPslQG
EgapOeXGwfmIYJsEwBMVJ1IVZFlPMUUFobmCSf1BAm8zRRMh+0Y5ytQVfMwMldDIx91DOwrj1wiv
U0oO/IIiM1vT7C+asp7LW+7GhzR5TaS8jFhWQTP/lqYpHrJ0icuOqIF7qXVai9rfgf/CzuNU8S1q
VJQ1JNWITAK5viWSTpRmFbpFWUA4rGCAEsF5y2TIyujrOa5PYULPGt8aJ1LLj/2lW1ldbY0ryR8n
bizSr2eGD+moC3t3JRtebp0fHQfYkmyV8LxepqAnDrxI7e22wKxUlK4cv3p//2ZrWqDQLRR6q6Vz
hJQA6jo/fCMrSq2eQzf0QVeT0uoscqLUkFTLwJJfAWXJV2vfWDJMAb5I3BLlBPT3zkc1TUgb37LU
IQBUuj70US6vcQ0S0/CWPbxM1omphDN78cPUOZNin47oNp1cyjgaGwSkEdzTP8Q07LHNDydTiZyZ
bd9I45WIVz1gXw8R1ZvrwnF6Puhuji1ykw3rcDX2K+QPnsoTIhEde7vfmDSFJDRMll77mGNmrNXa
G3Dkh1dtMissNGUgfbxiO/n2Rpj/2fyfhfhwDht6YNpAMA2+nRpOMNxopuKCgnO+9NdcHgq07Gq0
APsp86tY6pm5xuJ5JTZ9AmABGs5WIFlKajqkuhvmox4c5G4MXhIKNQJf+SSv24BCSOcPBk+d1BvM
IY6JLdlqY2rXNJqK8tMYVv0swD+l6lANPdJ8Z47he30xoX7Aiimh4tR8079Gx4teqtqEnvbM3PrJ
NiaDLsb3AZWsrIR59zSi5/hsD5h9P+GpR33y4/LKvhIESjyUPMyZCdnh8bmpFervgM1iN7jgJMyE
naGMXVhcu2arJh5DAyUBwbKNsdhQyt6/MzlxZ5ogAuxMncNpDK4AMghM5GAHrLBxMslDpchlHBF3
1oAKWhhzDgCd7Jt4/go2Lb7y7EDIHsg4f5b4Mh2T1BPL2v35mLVKqNkCI0gH0eDSlEOaPgbU5Ejt
SRYuY8JNrWdy8Nrwjc0z8cHUejMM0fswQYrnVcUGnIKMAdQOujZq1oMHUuGDgkLEmIW4Rxl4oXTt
uDLn2HbMMeeOweDmYGp13qFH39TgbVHgUw8TDpKrEg8WJzS2KGdWTOVEYASt+hifDT8ucVC/7oq3
2meXN+c7v8QwSs9rMNf+MGldajl1mtbzsOaW+0MjJq9YfrFOJmag/1QwLVdut8D6WhBFDR7BzDKN
E6qKpVyIe+agMimgIybXYU8I5H/JZEStjjfacEXW22qLR0EoI0O6s+4TwGbTh9wm15+4rjP2Zk/v
ybZ5EqLTHYAsRreuj2wXh+dZNZFV69Dv6K6uuYX5a1bfd4h0P5e9PsATXEpDQCQV330f/AmhEpJb
j0msVVvJ2bfMSXvldIwZ5ZkkcTgGUBjLEgp2VJxFB3yYsiYiV16A4p3pdcRomGjyDBvqb6JgH8SS
gsvVpXsKLzsv0WM937hUPXkmPpgJf/2kChrGk84J3yCAnDWVyno2LH74vFTa8E1i9lucqKgg2QXp
cUxx+cfbo3W5UQVuW/wg4v99C3TmNZ8GxJ5YcIxdi+rVbjqOniGogqTxQ4o5lOjvTkgtY/LRccO2
B8lP/kzcE2hjBEDyjFvndBv0EOhoq32lQQiEdjlUCCnAAi7qdOMtDWE9Lzw6qDnOkiJ8PUDmeUJs
xGSC14Wo9UwHL4mIIY4jNavVUYpjKdlkPES8NkZAvjr9VKPXdAgdwy8saylE5oWvSh7Mc3rkmxUP
0bN7FzVyEnB+tAdOMb+jTi3LC1ud2XbSSVDOGZuj9HNn0IXGPxLstWpNbUovpcj3KJ7mg/D6Y2/H
Pjk5AF2+WE4EUO2Lgh8P6PnaoJoK7/YOMQ3J3BoWnDA+6+uXKHbO2tolE6SPh/XMH2ElCS+JwT2L
ebnuHccDkWAF9KVN3IgSE2D8zmkaG5FiVqk/D6YolHO/sV7N2kyI+dpCpMOaRQMKWu6rQXkEKM8R
+LHCw28ee7r/JXftTjAU8lnIKRpK9acfF2/b1MLrK2Dbv8lqSwQ94rFoYgvAvBcLXmFCdPbg2qlf
yhxvhSAi/Sox6kIJ4ku4kJG+rOttx7hCob+Oqq92waB0CQSIZBJUD7HrbUvFqUASEhzUWJPtSHnc
Sp0waiGrlWoAxqHGftxfbAInzupS6mhI1oAPSdMr0hjPmNkI9lRigx7MahebOabQOnEeNP9yOdgL
2cssxVjRzrK8CUS3KCYAQ57YKQEcN9S9tPzbd6D3qy8bBPBXlPpTKAWzE2rbO01cMwNrN0VLq0+/
+GDfRc1gw+dJHXpuoFLoBXWEkRMZF0f3hGPYtMf/klhgGYvfiqoxGoCPfSwWVJYj2aGVb3gZ4LFh
osb03nNtpMxzdFo6ktm2f8YLcJXUvX95NdEI4D995ew4R580WOtqLvGpvzqT1YGXtdhMdSNAPUYB
sj7iihwIp8KFw8KDaE1H8wWunudDkr4yliTOBeb7TrsGbXTsafXz6qO9zwXW41FxMaVjsUdfu69Q
NjrhQcvGJ4+ma26yL+fHsTcCaCPs8x5+PewVjvjHv6iczwoKRDi9j9AM9+QJH1YSmstrXd9TPND+
SRv/N7ecEKqBUEEf3+hn1bp+m17N2oWkwacyd8AGLfdqHGJXNyjD6gh2p7trjYanuZjWZF/3AAn4
C3WDlOrB1e7XmwV+CXrOURknUBPoRzBmWEbAlaZFxszbqjSER+nMKpm0uqgf8f/7PHw137udQ/G5
TPvnQhd2TSf63lqsQ0/Iz9l8TphbnyXhHX0xSS/CSttr5TOldyAvbgdCS8PGpoTxEfSkZ183HF1S
gmZodjYkoy2SGA1jEreyVObFvmZDDxHIs/cnVm6xwvxjzkndBO/GZ7z3DVvPKYJFoR2r5X5TYQYJ
CC6fEBlRbyHn64nhXYAbPbEF3EQ2oVcc622FHddnx47lxeKEkFq45+I1ZFnI8RVOZOdqMMu3rtMT
4cOKwhQXqe07gqPeG4Qe0h06G/mnWUYy8pVu4oc+kpet+neqTwUeHTjqlqdxRo07vdPP2WiPCRAB
JhRxrhUFVonKy3boH7p2WqoE7sWzo2xpG0p0/sYfqElriW8Zm8W5COj1s1EDHQayoUBpEbXQkONU
tAIU4GVtkNQwFYw8ckN3luY9zfFJkoy8tTOxSGwCkGU4+jb05lb4mXytuQin58ym/QFgtTuiJjhd
MnS2GcGVeCShyKq7AWVJJXlKbmO3hm7HSkzBGZ57ZFs54OHG+49TOwuzJtcD1gUAo1Kf2s0gR4hQ
xyAtaSBejNoNuQMGMlPqCZrjr19JjuyTARMYtDoxcu/dHiItXg/DJscXh2/dgop4wc/ecDZGumy7
zxZlyOd5vEcyFlAi3/B6K8kpEiqH+EHaSO7XR81N+7j46N2N00+CmpYgU+tbdY/ZavOoe0wzEcnc
w0meiTRhXdtw7IvweYhlR3jeGivf+d2qnDgIqEFXypcvv/0OgGiAp/rqq7EQHC5V26SDLauF75+z
6C76ERXo/M7iFAHCzJYb66eqgtjYg4B6Gr53xj8QiVBEXBQG80NvMePU0AJ63/cM6hgJ7yQg5W2H
Q31zBN5Ezl6wOstb7wZ4S5G58OiO4y1UodN0f4q3gx7NR1ZM7pP3Fo8hxtDAGEgM6dmBaTzt0Moa
VnAUuyzvYj+0LXyuhyr5aEyFUYCTXkQbwKF526Ng/u7zK5ho+UbwhR1AjzNgxEFBEJ+35NXXpaow
NQmDlvn8Cmj7fvXXE2kBWSsaSoI5UErZea/VpU/G4o3balgkitTJ38V2FHDZZZgIT43IJfAK+e4R
i/BXBgBAG3ELji9w+POaCQW3EylmRQ3Ef8QxgsXiralhbP32h7089O//wI2AVzceagY7/qi6Qcuq
XgHsnbco5yiCTCqpyTSJ0SOSPNtEhJwjxUV6cND1z8i4dxO7o99g8Gec3KO8iIhxbHqVQO1JZIR+
9ifHDT4ipbHVfW+9Xp+yVqQZy6fL6+Xa8Aq52w1BHWJd2elgwReHmViZwRdGSM1PzkhYVbFnEJUx
SkrPycw/6AFU+qikzd1upyrAdarVnNI3SZys8zF60r6a6vkXg/plnhpNft4rcuAmOX3vPI1RTHjh
NfDPpgfFFpqiA5mZlhfmpzjG5CwnhA6l+TD3xqU8mXKp/t4/Epus5ZuNg0sIVJCv83bLYStVtdVa
deMPAK6xWKa6aq/c+iMW0MRz252wGFCoQCzudw3TlwCESxrbqBN3kV59TaSa6zmjZyreIUQSPpZL
Z29nOBqeUR68ObDvp1fdlvLnlbnw2VZ9gmbYy98cTO5t7yXWKQWP0Pd7YoV+kqywJSHu0RQFZjCT
5qt8AvvHsc8/TGcToWqgdSDSHU3HmhTqLxV0fHLqaUPW7PBGR1WEbFGptmXdl4/VcX40hrDyYa5S
C7Glixp9tGJ8exhbHc5IiBJ+X5QMd6GJe2rNexUnYE6toye2PQatCVDoOtK5OsvEN6RERw/R81Ya
ZoutpjhVa6I01IBe/VnVUHp5Y05seWb0J71TT2uW7BWY9AregIP63I3VEB7Z/GR1WORBfj+q6QlA
tvaNnWw0ZMguPp18145uzbPDuRFOdCpeXF6VclzdufTxSAnZHFvolXh0QjpcP+N4ZrvmieBoD4fE
a3IiDkz+h4ZnvBBtb/mTLQfKzQMC17y76JJr1KB1Itmzz4bBqTP6CEeuc2G0K3JiRE9FPdheUgu6
b/bvBkmgGyBxg5mDgQSpjVQCnTQGITTDHSb36V/9WwibJvquypbM67oD3oYNZP0w00LfyMm1QNNt
yGIM0MGEp4l7epPUTXN4DB2SKTLSL6UyGOQ/9PO2kkChJf/YohkIyuvgCc05gdlbi48exUPkC1UR
i35XaVnkhnAWYcnjkpP2fqCd4+IgxncCXUC3KpwYkjflI9FMK6Zk54NIaceNqYM8w2uObKAHGrYf
HZ/hEt8oLLfis9DNUgsWpcQGR5IVzGnY76Dwk7xRi3lY50l2sSmwH/fm5LEgY6HMGuW1f2e24E1o
chfNKoOtEBdJcoAwyxdRP1Hmou7zoCnKzUBFXLpVPZaO/EpSiXIHaYiiZwh9QaNFKLSeUydTw1TB
RjjvNxZbsT6Q6HNPf02rocxY/kk+5lyia1Ikefo4M97q2ZD5WqmzdqMksPcADkoiFMpuf3K3AIKw
eX4/JYTKMhCG8QJU1HH/bmVDYOUY7czonODGY8sh/LNABV+u6KWLvpJ7di+eXMr3k7bC8D/va7En
Hsy/P6RfCWNjB9w2qSoQv2VOiyO+DOVMy7TMSUkeK950EchzAOI/6ErfF+g7ABdWyuUfwDJdDCaU
CkHD4GtPm9pkbGgvCKhMGApGr2pL0vrzKQD7ghac4moct+7kyZnLRhu3VgoVso8GkXgDX8Kgq8/2
GT0W8IP5iwVkftK3LTCa8NwBeoqT7s2B+HeYeQzM/JdjALqm3gsfeeh0HfvADAWnssKuBq4cRx7E
i2FuPsbXelBcWDk7qRqiS3mUU2CV4w/DnnSZ2qQaT4rEAeCbg2ie8RCt7Xm1ose/rXHVaximydb4
wcN55t0O9mOVR69eWT/amR1KILpvm5V2jp5XZ6sXd6HH/U0NnLMjf0VQi++y0vAbdjOmulp/B+ol
YpR9+NWznuuhrrpmlCAavyFSY+lf4tznvO6/kaOZjsd6nTtbt1k1zB2qbtoMLtMAOG534FcMyvUZ
27uAWTWbYIdW0vCj0IEfpKHYWkq18FadDO0xEseo2Qp9ScgBQrVTo1EnuYm+ASAgYabeb7EHMg/m
+BnFGVJFpZnp/Rqz/vs4297WP7GyazpuoN9N0pl3/mX0hgW0QKZ6iBG8e4XYPlZA44NeYDJzdH0E
5TM6cnpL1WH4uNXgIkACMu743rDLK6fAwnv+nm9tlnQEITrVAlA7OmBZZsisM+kTgnOWnG23szYU
Tc7ImX7tPnLtFel3aOGZ4PHLGQmPL3FCo9gMSQOuyN78LdEhwDwvcVUD3s06XPCeZewNVA2riDV9
mvWTa+qMzEyHIieDtV4GgVwm1AQpvn/cWE5uw/vq0A6FEzY/fuW1g8Fc2ZRlTVtgNI1NQOUCxGc0
a6RVGG1ghDCKFg5SWu2TGAzA1WA6PihPg8D/gGy8k+nWceMP+fzQEbHaA6Tx71h3YBG6WF4Ajm4b
NVoLzJxc0oTI2WqGvGnnr/SMXs94W7lOAXcVSxWj/7OfTZHOoqHLex2jLsP62VRkpBjbNj/xeGQf
92ZDnhWomWdedP5dw+xl/3TszQDNK9+eeSTXymhONKk4ZspyocyfgwuY2t+SF1e+e2DnHAj1t9EM
FhKwHV5cxP9G5wd9m800iiS1/31PaFovFi2FuGXNKmRXS4BCvg+Wh+6kADlcCW7J1kLfuWWb6tjA
wHSMIXhD4o02RqGQbxwzSyUNWQJdxaLyHSKQvQ9t/ES5uKrgEjCn+lRRLAd4XiUSdsMspfNYLL08
1vyVGWCf/hsC5z0Aniv/TocXIiQ3R54Vf/NiVFgHsfpDkSt3w5rOWij+vlRwHaufRBcGtKaglUEe
iqgdj/sbE/2VdRzh+G+773H8r+UO+rkA1ViB9X6eTz3Ro30wHBQ92L7yeZwjyMHKONklOYqifuyT
MYp2AHHeSpCybiXJpGeWHydoYm3UXlvvYvAkFPXJP6psnzhmvcQj8N0fUaMkAXvHohhjFkPmOY9g
L0iqNBdqxND0V9wwliwW29wrQq4SqPMXZmWl6co/7yc11cS5Si3u859SxsAH6TaeVOF2xNGuQwTw
ueqnZquYeppJ2NmjZ/bGvTaGk83fAIoY5DgClr88N2xsYhgntDlubgIZNAJqFfbG4Z/kwPoCmNEe
LBEOUhdmN5uZiz6Qkuo4KhC1JvIsyDsZL1rcVpiNLKs45EwFFNftozPj6mUuHnhF3rAysQVurHBK
Fafp9xBiqIn+5aWW2pdNjrBbo2aSZcsvMY7nitWiYr0nhtTUx8kmazU/gIoiinaHJ8PuxdWM7Qdw
MocXkCV3q5pGWxAdkc92XIBDpgJJyL9dH8BHa59OkdC2G/pdNk98Pcb6Np8rFTsFtPzfuK4+39fr
+xJt2XEAMhhkEx6C8Fqz7Hbt/Vae6ljrudVs3yGWsmBtg+87UC79icjGchz2AmkXdb274AamhOS+
APO1vpVRpPQslfhPh9sfy7e6NxfCRiipTsgVYBoJCwdFwLVEgHi03YiDm5d9sjUxiZEGnjulfzWD
ZG+TCzA6RHCAzSszI9v84CruJYKv1F8h6b/0067m9kSnp3J7oBJwKIx+MJvH80jUlaaG14SfEf5W
E44FT9pTsjarPpAgz/LwO7sxvsdBOL1VcmIHKXQTyT89almHT+HrsvOo3jt+UvQHFqyOTTs2M4nr
N4b1HnxcGOZ4u0SPtqy/HBBX5AqGoTL8lEcL4JYLlLUffQ0VeyN1HIWzLbT7OqdyN4vR8FalPRu4
IFHUxxu9zKv3aUnhFxsj/bF+9z8GGzM1Xh3coIkGq8UD94/E6YlmEUNgbHo+hmC5Qqa4nQGZlwzl
h2744YzDJxihptjWYa4AnNfC3lvJD2vaRHYIN0e123dxOKV1I6p8st/mHsrfopu9zDyGXLzxSf1C
zNM/pK/HuOHccNq5ME6jnnij1lk1qxb0v7VmyVgNYZX9oVkEIDNhZrdFEBvo8AGTC9OVe0JQSlQG
XClRJsWKBKgv79S4r7uLonNK7WI7t5ZvopPxKDdOpzhR+W2eHuSCWYMXhI0rY8AHP3TwOABgPP8U
YXNjxqFvB/QgWyAmF3kCNLkn+6kVm4S3Ka4mN6Nt++FUIquX1MRLjoG2whoF+QHJqtrMXpBp4SkC
mERRJ93teDr3p+u6DlsvbBOkSFVb0n820dacYSSY8Ka2PTWn8uhQMm47OznDhQpFX+jtN6Vq3Gid
jZxiahsJfIN02TCi2JsXx8iOJQhd3mfS4P0LkZZXbSclxeWy82wIieJC0sciZVmfvwdN47qjbADp
SjvkKfoGxtz7JzWGx5IbvgZTqrGzYQuUngqor1wy3DzVXVI9DMprdFoeB77s6DT82c8Dph/faXJY
7ps9r132dbjh2Q86TRFPI+3Wdb9kOnfmSyYpXKR1DgMBkLh6QJ5NsPdpLL0Lk9EZh1mpDez0iu45
QNPi9HImMquXjn+ViBckuVGYqI5cdJ6OvQmBEtQV46dOZs2izwzZvt0aY9iZM02xGh8m10ISWQ68
HwSCkczXj6icX2G7EmhVpdK95KpDB+nvD6CBSZgVyC4dFBnv/YHrr1C8RG6iFp0Anzd5dCyEupMX
cn8u7ue2OT/jwEQLlX3mE313FaPMSw6VNpJnAlkKJbVRa1Z3u8/9/1anwZXnVYZxJUmU/5vVt08r
Gc7gAD0Mtsgy800Qoal2rAMP+LQsaRh1fidRDdLSObYypiUGH9D0pOX3OSR8C2u2c4xqtTwDhzju
crClvMRCbllgz/wGq5jjGndfq/bqg3Z8u/8wIGR1gAD2TkHbnk5jIcCS5qvzWOvQeKudTs53i0er
RgLzZkHUKMLE2C88l/IEgSICph0nJAniDZ5ifH0MoDyOG96klCtRXlPZW7JtwoPqSW07CNP4htQf
r/OItngxXG8jj8B7QPlq47+N+eZ8ucepYDC66YGu3BwHEQvI6VLOjh0gxzS9bSGbGUKhNpWnyAI0
NstQ2C2PKedZnMWcmytdECILkP07cSL5e2uxZxiCIntCUCoSEe3548hHwy2G3lpTTRCCpCxjYi5Q
ZFlIgMz/TMDn1iUkd3J2ZlpuRGTHUuLEkrM6KrtEfcWk/GH3zan+RpHwQMOJI4AbrO0ooAZqAfBl
ZGvP51Q09PHW2bGLtM3efrE8W4btTkBMSXcPIIRs5LDYXQlKI/EIv16FlhAQqEbMlAOqY7m43C3r
w1HdmaqReXL47yhanVq/8eCNRDyydlU3pzmt9ZrplTObiiTbuXQkuxoRDtXQMtRzqebbVXUOgs2r
ZC7FQ3QRW7Zg8xJhaAsqcV0iq9W4k8he1+QgIca8mOr/SVXrD9yo9qk0ynoOb1GbNSWPg1s90ks0
YxBtroHQqrtRHtP1vDraKsBbfFCHfia/K1V9CWYK8Cfc4VNIrPpwi10/ixVM3m/bzr+CjdaFptir
wwfXgjsQnqgILyJ2LPs+SNi1SUfchGlYIIEGJGYNLZHB5R7E3+1rVHoWx4fTsjoLos0ue0ny+8Qx
mE2TBMIen2CHigrY9fBAIPq58T2jLuX+EWz2TPc9ndRh4cX2GnJwOubLoV0h6ZzIKhA6oiFgQXm9
lxAi+AwCYX0Z/UqXYKHiSNAhj+cq2fLr0oVVvGg1ySQ1zFyB02BqR9A/uKdSI5vQGmY8JZ4Zt5pO
CvaA1pRklqpQ7ZFbUZlbZSCRQZXLZ8WE4XMhMQ/kecPTBhrIVPs/8Ev9zA/PxXKPoiR3HaCU4Fj1
d0pjzy85KzADCW9FkkVQNGzE8TxY/lJwYWpUKQvQRD0PdAodo3HWFSM18ww5YUEbC60FW/CUEpFu
EPq1G29RBTN7GIwYGykEWN4LxRVmusB3YMR2QokZsiJyax0f5nVbEjRVoY+dQPTWrL/kfxqOUGAm
mrI6cdwNudvQs4+hvDSkHOwpsmdvoYYZ2qe9K3EOVWl3Czcol2OYQfkHay424e91lYULfQwH+e2X
nxNoLBRGUsmDCO+NCdPXbpAtAXE5y2SlUBxxF1q5J0oCoGLCuDrLhozRWE3damiVhbCX1U2dk0bm
PbYB52XBTsE0J0oDVN0OAY15mFfOeW95zXGmPEKGtqPYZ/kdEXswxs+NhUzOWuuK1e+3+QwD7uJe
kzTXqk7+jRPxmZRSWXrm79ko69NQ6JDtPLBeR/zbhpxqkseoFKfoH8/8dg58PnGT73HLvmprsKkO
xJ+0F/yXde2KSDJ96wmd7X51t+8YLLvm433P6Oij98gK8jiG/5NYaN89oTrb+UYwgA4Lyo5UTvuX
nMnwYwsqDtGdfjuQC1k+mxqdhLxDtptRaJx0Nwqs+7Ksv0G16r0HIVWCcQjogqwi3zmJdBkgQaBU
KHRr3VxW/Mx/pN5oKDApUj5oQneAzezAmW1WX1SxNKWe+xwrhS4OBhX+/45Y9yToYCY/pBN0Z1ar
76l+HryPyG+SAzlHC5oMR1Nr9CtpMhyioWvEBrXaXUhYxb283Ykb3m6rS7GWlWvqfIzOKG//uTwr
kErpTNlW1t37XPlDneaeV1N4VDZy6J1HkLc2OGDqhFkzZn2nKARIAaGVWfjADXAijBNVUdi9BP9i
S3u43icnxUCeqC/w/KLWuru+Yoz3HQPCfeujyY+5a6QMRoTOhz0jn25xElHHODEl94Oo/KaiKrDz
jaDkSZrdiK92jJ6DJSHk6WYBFHRP9ru/UwsqC6zolUhTPBLeG51zo1elVThUSOOFG16C/E4mMOYy
2G5m9s6Yje0pIIPYYtBiHQG1mB46bIU4P/g8g3xGkSV3DvMKSuhRhx4VIcKFxpTCI0iPjDqgbaIG
Dql3jXwZOhEpgw3r7aPmF3Q4Nly3d+YyVQN4MxRIDLA2bdw2NWGZTgRDmODl8ISgKPzFcn/N9X3E
d84In+2C+5tVTLwlVgj7GeFVG3ITW/QmPmSgpyBse/tt0Lkf12KJDOGY0A0QqLUYQRDSAflOtPeo
oItcTMpe3S9qvMwZ/XvDO0ZiS8PP7JMdktA6QTJOHb7Zf4XzT/x15bcyBG6pA3ZXwlwdry7vgVbh
dxs1SBGAla+iXnH6x9d++DPMYXgGvRHXEZpAGnjD3nBDTGdLOSlxiZnVPcT5vcz+7zlv8sIC09Ja
G3nYM2GRUl0EZHSufvK/0VQEAcGTDygEy29Aa+6OMKiUh0G2dPrFcXSPpr0pA1HJ6DLqnm4nxCWL
CWy4Pqy+enT0mUZ1bOLZHuLx1fFyDFcHovtX/jpg5KVfmkI0BIgv/0pCAhaA88UEF8YzOfz2s0/I
8ZuSRRGUoP85ePyswB6dXnzTM9pDP9GljD7Cf9TkkBcJ+y1oPny9gnzUZC6c4ZrRuB9AQSaos1Yh
pfc2yYpB+JQxG4shwClhd9cgoU0Af2QbynNEKTCwlxHwP8TkByDmjK2Cq2Q/xJo9MlK3pfOCJHBt
BJ5j3bKT9oF6D2mtYkHeKc74EoPPiKFiemG800mMSMLwscg0PScW6lEl7BJNqtXpXk0cBxRcp0u9
TYtS5MGyjknAr0KITvHlgwrikFdWTfAtk1sWbcGZbCVTqz7OxMMy0x47RvWf9yld7z2vqpQwFY87
Ck+NRRT8RQ2/enlOqBo0m18TlNjSs/nh6GOXfG06uytuZ0A60TRjcmAfxo2vyDyp1vQKFe7zGSPD
LmcoMuzP1lIButk8WuTf14QxsdXMuI0MmM/x9H0Xm/neK00LLT+VWnXp2GPwzjr9I1YCzrgTyfdb
2uIRdXoPgBe8iyWsHBw2Fy+Ew8r4IXWikfE3WgdH8E0FPK632V9a6/5PuZLEVAD928D9Szbqk3/C
7AvGEgNyYmZ8u3eJOJaACWaq6I4sOMPr9jPf7ckTcJJK/TAw71Ylf+BreBU92gvdckomWErHKbFK
ZTvqYD8rs3sN6MzqakSf4uS/H2+0GpfKWGc5H2o9Z5rOBe4CkLPGOX5TYnJ7CT/j1fNP43KasH+v
vlwX7GIrm99VdRGX3+jmZi05am1GF7A38Jbq1HFWv68OvGUmW+NKqfuuz16mQEQsThCnhBmA5rcV
HRNt2m3rUSd7w5LCkMqq4KGk+vX7vo7KNpqkxxKrI/k0+Eylu1M4AGuOKUL65j0KqBbtxRaFlZ6r
kZcmJamW3aYtD4UoWSIhsGTwpQGwbryfTBWtOMVkHDchCimGb9h3JfpAnyqtAiLEixY02ht7uFlr
L+NfzO04dsvSGd1l1zJ4jixmNLi462FVmTl3CsDQEV0r8WetaHuHdBh9p6nx7wUXn5ftV0NPaOPW
AF1xwgn02HynxhiW1K3hgGUJm7DNt6+GErJRHm3GE2N9Oo7Sq4JZdX+nWrn42j9MnKyWk/pCMEvn
lAZdEJm0iTn8b4lSbHy6QKq/76YrShpAvQ9le2CgKonn/GZI5643SP5JSTCn2RVWKuOBJJ5zID3s
YzlWhTNcyRMU4x1yHnAwawhYyEdmQ31KHaBmgn74xplAXsEHSB/ilquQCsRyup49LBuUFoe54Vv4
jH1XnACvmN2YycPS2i1Hcy2AxgvBm1r7H0IEXMfHEB0pCStMLQo1kTyOBMIg4MaaIIjupJaZTBSB
FOmcqYRxytYMqDIhP7WIaKpzW7fzw4maL9KyKKX46RRW+fpjlzw5kr0zdeR3mjF7BQ0Tb3wznP4w
bMfHnvEgIsp9SiPpovSg1TiTJq2QEFVPyeMST3MkV7jydoNTSVKSSl8QutuGabZhoNhx6Ywj1TvK
ine6hoHRxNTtfXS9w9WjyqUnDxON5vBnIR6ZQa0pbI/OJyaywLSi8HA15qkYx4TH94ook8tDkSx+
CYsq985Poe9oifHC5cpkfKfkkjlMg7hFACkPDNMH+KkEr2IRIgOxzMBfM7TxQzD0koN3isVNg5/8
B25877D+hqTrhrh6CIxBobVqsJpig03k3S4Px1cGPbDZermIYcE1Ow4WWNXY3QsiJwCgXnHNh8QT
elglpad/EdV/O4UiQcjGLOzGab8NaDT8pxNZNQtA8Np3SdFgDbPbTedU/G0QVkm3XPMXQtmA/yRz
dcMmn3AsA8AZsLYOF1KYYBnuNy32OFso391cE1TtrzYpm4RUjKts9ZtAtTWlBTuAJvolaE9hGV2q
MsW1NwqMRLloTHaH8pfDPpiVxEsKlfBhzhYJoR3ba542OlKf+mLEQyteIUANoGATZb7VVVzuZMxl
osMbLDBZw66+DArYXyCOpgF9kaBh9NVJ7g9p3/J4ZEEIV8RcVDYEdmvU04z0BBLe8wkLZXLOsfbM
z1iSSbZqsQw0UH6FuhJPaBNMYUBia4kMk/JR14IWnwSHYp1tmh9p2baOYQoMr/CjWTfKmypymV/B
/JnvsajHwnr+lA4AtdOGF/GTlkvExrvXamMLVmHW7cWVOd8HfjnW1DzQIqvF3N1fdxQ5GuduNVdy
eSLzhxeucy6wK0KoLUek946YekfV6UVR5f0AbfzHRyNSpHdZcfu5q0dhgCIgevrkV+aWQRO85oli
BlimIGgNRnrI3jFCBcw3Ytjms8cKAiTGL+jsuGVlOm2vZq5wZedQRQy6sdLE6iAFvXpqjIHlR/Vp
E8IInmRK9ouFtbG+p+6hmMjWgFetVSNVb9WdqC6CG6/6nuHKEtkHS5wGjGvOyyodxAemLFXWHDK7
NoS/bkiddg3ZD+Mp9e9DAm3SZ1tzSPB4a+yGym8GPx5sPU57lm1xIcqMCC7ZD+zrAHnjtENrx8ym
bpfEDHTzDxe3scK99WMXViO8pEO7knjFBjlJiMSFhKQm2wTJwNLWDklx+HPymSNcl4FjKe4xXXZ6
J70nxuRrsZAlWv3Rr+T8Jjig0OTvDTc9cSKRGuMJTUdACTfTBD6GbhQl8/c5ovJ5ZotQhe3LZqUG
OMDWUZ1kI85VERlLFIvbv3R9SqZdfzAN0jS5Z95FBZqGSSxEpv12L8NB/zvD5IfdVV5wXK0l7oLy
JmKjGKKuu7xudmNug9DIfheOcCBa8rvjCN5GK/RxfHsoAGUChzMcGPAr6yiIH6CnoySi1DsyvRjH
+dj4MWfLKKxQ6wJqpeoxvqbyzo29ySwMlBRE59HLQ6H2x6l98lkEV9MlZdJfqNng7h7BCRLe/QAj
aj1cP+dPA2dHLqhYPr+ASNPheSrXM8haVSt32uqvKk5ulB2c/PuvObW9H8x7W5Q8HO4GFpkrD86C
jDYwbWVrd+4yZu33xS5nC56lzM9A/LghEiiuFd7ZUv1x58lVGL9jHaofreAOIIn5Xblnidee6kyF
sPUWE50cFVfV7UgxZT4YzhZHpU5soV54BtVuzhqeEjws1bE4xvyK9evViOOM4QhNy9uO3Mi+gUDa
mbqqH9V6kuiRK1cseQeLFbThi+ZalTux76y94vHrRgj4CrryuF+Oqy1OGxJBwQkJbXGjqiVOWIMj
ZCBXDcKpQ0oHj0b4A9tln/a/dqv/Xcaib+NZTgfbgy5tT6ThOzhlN1VMIdjKw1ZLf4GUnFkQSC8l
IFOmvVymv829YnBpd/Ku7qeZ1tB+01lnfQofgisOq9oiqMxOIBsGHDDE0TerVrn06fE3gt70ilVg
Oz5cYFoCGv+G/jG7maRZhbvmrRab9UGsrieeLJQeV6WfuKu0vcKk6nAdw5p1YZ5nIoRwWmlTlLh4
UNhF2X1AA3x+mGJphQ7WkAzwCyYd7uPgfYOzx/eXgeVJWK9T7dBRmrzhLz4UfgNQWT2HM1oJDhOk
LN0z6+ZD6eArWjW/UozwT/buQ7PWivxxzXUk4P8l97qB0OeUapDF8lWEUO8hvMR5ruY8T8PR0aBH
w4twsb2AN2T9Ij2XK3RI9Igx5phaDWOOBDPpUskpJ2VEYosspZ2NAqd22hJ/4rmfpDVnor4g4tU5
6UJEmC7W3b+CRAsRNidY6YPn6mSa6BX/L1eesWhrCethDEwmGcqbtrdQpJNlqMJzZM5lWaRTP06p
978RtyXU5g1hH4RWgivf4VdpiljAzzO496F9hRLpzBRKlPMmZWKjY7EefR33WwaSjhIxQcNUqLJa
7fl+sD56U8MnbGmqPwYkPp7sOxL4KP3UDU7/2qERDPaDOBzT3BTlwD6qVtks/kzqtnuUiu9XrImD
fytS2dL3moakwge3EQRzvyNSQw7ZJwuZw4HQCV6B9nDsu7GFhHYFRaJXSIlqB5GEu+7uNr8afSL1
F5eloiu5X2UqaU3ouIQ6aZam6u3cxD5h3lho/Sy8OngmBzSNqWFA3y4TEaSSdETbeDTTZyrWha9I
651dmqXOXiqmqSPy2xCbcl17G02Lmx6kRmF8iSrVgVJkCoOsdgJZysObGmC11uy+F5dmtDzkZkBa
r2KxynZCJT6WAzfSFHBO1+cBXcHQHqHYM/9JJIXG4HJl0BLcWeT6A9drRwAqad8F5MfBc8V4HteP
eYjFhqacevEMn3BC1BFFKu+I2ubWLor1bJrhwWSdqS6yGY1E8aCAOSq49hVrluOazhDiX0d+o0d5
X7iYE6QF+x78X3ZA6WUO4AcvR2WZyES1hCuwPzc4g12wZyxet0Iv2GYXSyGFTf8gkklcZbc3kM5Q
+f095y+WjMvx1aZTHl+kh2KHpSRb8K+9LgrXWwnubIUsqomuZmRmrzasIah1pOnLiMhNXahWBw8V
DPpyw4pkJaKXGFvH9PEXQ+RIilTNWNMYKS+NNR0817isS0NJVfga1eQUjOtc24V7eyJdtUBUUk4D
fnqdrnKzU0cuXTLSu6ilsxPsDa9lyPJPvUggpKpkN2XJRZV8uLAU+pkGF6R20Gxr1C+8OcALfd5W
pWf/WjbJEHr3gbqB4KmlGcebFs0L45ejXuaEEdmYi+fq/IHvWhoi1tdoFBGs4jFiLscedWOIHRD6
QbGK6mPu8K1bJQPLZoMOgm9PaElqblH2ELcR+h6S8Q2PyJXZaJzrml41wbBPPnXjIDfEqfkDX2Xp
3yxw9ZkgJ9klOqsEwzCgV49vZvZhM0VQvtAdeO3Z/AcvwcnOYODGP5Ju4Oc6+yU+J6lVPOzzokIw
oKpbS57f/IOjZgZMFfLVYdtaEmH2jOQtJn76fcrACYkPq0pzgJp60CwJZ5Ig9HpgB5a6KJ5cjKqV
kHHbIWd6cPkGr4WpIe+X1ASM4zH50v7aP94fZTkSuQbr+16M7ryZ+Py2NEm7DTie2+2jxp3mzlSZ
HquWeaRww1OkPVVTTutbxf8DUlSh9KHCgi6uUuBFeiw1ZL3o+PCgQdqD7A/VCHWZ98INS1H3REtg
KucT7kaf8S6v0VTD8vNspUq0kGHjzGJzn5ipx9kqMICpZNYWhGuZrsQgjnsqT4mijEm4qk82eH5Y
dfEbL21BHu4VJM3AZ53AZGRnIF/eNpSsd6yLXQPanWjx9mDwzcSxx1SiToFnZCLKLH0I4emMprfQ
bh9sAU8a/WApXN3yetL3IAJZN6kc1+ZZCJvCuMwDzQmXs6rwfRMeSOLGnYW4OcT+7Yaofy+8nptp
PsWS96IBwuuNxClDl9fB2pOOgPynfmkMMDWaf3C1AWIXVIa9dpjnJc2KilXgXfo22zgMX6Pv21dL
scnqNSwpJ6pPkIyhaC2Fdk9qbvmtDS80Ji6UcUOPtcrhVHK4YtJ7uz0eFZX69PAsRFp6HfDBkQlW
NhwqY1t852R0I8XOionJ7T/dclDAAg4tcIrKRGUaDy/U60T3cwWqdaQI9cVkulyNFEfXQzgjergL
R3izpcxwC/4tc2+4BFnV2KueD6wfOnfzdo5KM9hvjDmD0uchM6nJpJFjOniUapDsBU3O2gXokRXv
Vx2yWM7uq/n1XnraMhBOipWzC/BgQULnZoUr4GMN2Zd/h7kaDxRpK9a0RRPnstIJy9gYG32wgwKO
J8+5OBAXZMdTnzjMZxUyaTToJRi6ZmaHREbxzis2hvR8LxwHklj+/UQWAtEdL7Wcahv0tecIEAyW
4xn8ADR/UtBPbbxjwfr5giiEzRaKokbR4WPnP9W5AlPHAM1P//W+sQQOxK4lS3B0S4eld4uuD9lJ
UiY1tL71X8HTh8peNxYFBdkMOLnnFBBEy4Z6CUCXtOJso1yGfPaZD+M4F//npUTFQ2LtrQAw8SBZ
n/Jd8+Tn62PStw7YhpB2/Apg2D5Q194dW1polCZbcufeCPel1vAFQG4qJYWNhqAOcdU5nfWqcozN
DeZhPCHZ9FxmVE70oFY0UmIlemnf5Ul8OSs8tNFuRtR0K80VgPJqPUWT4h8yKoB2axcJRkqFpXWO
pzmempWKxu+J7CgvYpaxDUQ9PAW+F5AnKc+EyDKKOuHpxEMMjoQuSLqyU65UjRQ879m3Ud4rxrDM
+td33Oig74MmjiTwdyLBmaiCPQJlA4p9hh7FJQzff+ZiJ2FIhfSSIX0p/xuhc7R1MbOkEJQVkKyR
rNU5aLOkays/TkjYs6blW37COwKrpAT0FMBjgNQmqqbytTY6lfPb9UHX116a1MT89Vn1hj4+zdlS
OaANt7Vg6/ZRUvy6ssHBRIjwKuXRVe7kw3KQoOXNznzadFPS//UWVL/B7MQXX17LeAJ0L5i3A0z2
PtvRzy8IFq8mBNBDhfsB+mZm8NliL/QrbU/c88kLhPne/1GkDa13R1uPxbtYMnvR7B/RcB4N6fTX
KiA7uCHugwSDmp7vOuFs8mlwf8zQoE0sYtQrkZAfJ0Gi0Wi7nlDIJyFc03zNWknWqm9Ajxo26WpR
esJBnoLkT/+X8LydrI24c6CDfwjystP3goe9EAYYwIaa8OHwgPDLBR7Yjh/1Bf2Zpzv5y9/GELIQ
kLL1+aDhKtY6MMLU7gzkj/Z297s6pThIZ8uXOEwAqaC5pEWud1umGVkfkfKMmbgXg4jDfZBjUYzs
RAoib7TVnEZuC3C6qb7nbdqmS0xiFa+bp/10ZJ64+ObnAjTuq4WHGjYUn1eMiR0MmRP3CFiYW8oR
J6bANJDjxoOlv5ExDqmZAj1kAn10MNSg8EXIxgOmn/UOfBCpqfkIZOHXojji/6zU6X8AjheYPl7a
6Gib/0iObakTFAxOWBk51PL/DVk34EpDiA/3+KyexLGb+FSmb7cWfb708nYGOYtYVPmQL28XCQgO
/u7Lci2JSk768+m3flFAdrBeLdkf6haikXyx0vB/lzfsm5qWl4tzGzJpKiTLzEdhtZ0kuWMAW2bC
PaptpFXsNZE5sCSB02SOvRsIBB2ozyIaCZMzZZSfUq07mqtzN5C69o1fclENcfoMmH8eBOJZpWwK
cJywI9lfhmRJ9zw20dk/3fVQlpsi1L38e6AqwVVSSx5yXp0RSjSeyIFwhl49omCv4AhV/5Xc2ph8
cKEKSHES9QZiBmGS4pUBOAZRCkfXAMzeCmm1a79hgjAZYznRv6WMtg2r+EAKUlVVLJ8c6i5S7eLY
tH6dDYy4v+Cmg5137nVF4fP1DYuI3DMGSucMKxCgs/jX/Ptr6UT/Y9m9zIyr4SN+SDJArDgp9EaF
LRWLrMXC7uhAIDYDLlCTR7qjM3hJMIzx3RoBGBYVXt8X19TZF2ZcydgdmMPQ103xPlGmtmTDl775
BbYN+lv9aBdJnKT3Xr/lu6lcAG8XSeYNrg1RKG/Q81au8jutV6C7T9C2elY/YEcy4DZJL5fF9SQk
I2zFy1fDWqGxC/TwHTXOiEjpSzAeua0TEejPBsIGaWyk3xkTeAoNOm5rMPnn+PUKt5belOvTHCKw
KSKEKiosy6CgkhITy6LYPvG9WkdvpprsTS400XA3oinsjxgFc55+S7Bfp5QF9pRhK48mj5X19PP2
0Mj84FocDbALVFWcP75TSZ5u+b+yEV4IMOsbUPCJKUKTCB2rb1VXghk8V0BSoUUWtlZZBr8Li2l8
AogY5U8T7S/l5PPawUrQHIQXHqxW65BtOqxbY2r3paTcmQLdN0x7k9ed4KouAhkC0bXYXnKOxm2H
XSd5ZqIzZPd47ZXSvf0uoFBAkHgEa1FwWcts8TIYvCNisT2F3O8PhP32OsR9RzP2bcEBJRt2KJ03
nl1c2hf5EZlgiJIdLFe3FZjBdQoa4NInjcIKKH9PyMWZ0Z06JJbTxgFVWwJZv649MtTkGAn27wbJ
vUr1udLejj/voik1fvfyh+m82CkXSTDwk2JnhlTCqz6nreeb/6SxLN+SQ2/UopE/Lgqs0mSXoF59
3GGr11M6fzCmFPEg71VusFNkf6siW3PSaw4JjT8h5bNQ0T8O3Zwb6RUW2tSTNvGwLXveuaBbf6oh
H3OqPlIk5E+/WsUsbQSSHIacreR3aVbNehc0wrBvfEgi5Qbc4sNiFhpDuqid8ElEYAFm0tnEz2a6
lYt/khlghNXaSBvwsZSJ7cPkwJIrr3tdSxcezWECjd77lnXsA+I4yYuvXDD5u4mVDUorgvOPi8ke
4nTaNt4UZkIqjRT6+Lsj+v3o3w28v20dOAKj4Y0AukxJtJtc0xnZMKsROXjZ51TWUM6iGPj0SJOA
WJ14nnx7DFt3zMs8ozR2DqyKFSvQLQPCieQnhY6kkxT8M9vzVO338qqlqMKjuzc+qGCgcSKbISsu
oxfk7ZrB0vdyqYU5nTjehYjhwPtuAlExuXMDf5oexuZGoahn7lLQOsPTPgb4cXU0RqmMJner1uBw
HWXF704a74GpEdWvH+NniTsJDWSFVgAOU46ewPGhN5u/qJc76CRpc09/DAW09TSQ70pip77XBTNG
r/A+/42gzWwEXNp5sTySe2RSSdmsDryTQyGkQ+qfNz3bLkGq+OZ0wghuJ/n1+pjnkxXkhSVpleEW
tkO55yxmw6fKZJCD3EqdZfamV2WcVUMKaDjYHMoqPxDoOmu915ATgWsJQ4LRE0s1sN7qAH7CUagM
uR2BeWIfg2YAb8JFsNxdBefV3Cr489OIkgK8GCjRfxolhHjlBgPp/tuJ6WdGD9on973SNk47DCzb
dypM2ZVc0NkngUrZAESTpE3qCWsYPkr/8Cvtbl33LjK08sMvQs2wgRYh0mOgh4vjP/KEkKf6hrRI
Q5vyKYQCEKMpAUa0+w9TQP0IDbtGc0P57QHZTKApPQkarbPBhZbRJyJoJkfDJV2wSyUIcoGRvzUf
EsVsdQjx8XXyu1mz2Gl4giHfVyNALJudZkXcGYFeKOYsKWPX3UGmEFl0GNtk4CyBukV8oTMrmlTM
FlbwHksAy3sZene+ilKpwvZv1HcyD8hwEjQyh9N8KmhC0ZQlyZyPmVxuq4F1nHekma2RRBgBr0DT
oqTDQzOhhpHvwB3f/Z3RyeIAjWjjG3FRseFwF+uW2RimpFkUtqS93jjg46IhCM3MYw5gokAyY2Gk
dWZzGL0daonfwYd93O8VRXhBr2XooI9sGPMMa2FoUZNS9EtA35Mvo9SDnMoTgTr/j1TUX7LVqxPW
WNIeh1NLO83+BXWZH240wbPX3sXmfKPLLpdJZzxiXTx2bgMpLNJuC6CCfHTGmfu802+xMxLK+vCJ
8TglHtyCoFsH6rs/DIrN1PV27FM5hZCTD9OP6YpzAfc7eFU0DRACgrqWRPqd8tGgaHS8c1G8ZCSQ
f38+1oCe+09aesvrFu6WovkTryDzK0/FZjMpA6zQpjhwZUarYyVjE5Mso2mmwtNtWWpwz0XBmG/u
EA54nOlBxXzSYkCH765pKG/GjG3nFQKJgN4Tjz80LhCU6yP1dwZXYN/aTZfc27HXVOErGJPKsKL+
vNMBsAS5PSS5mKc6SGdCzi/E/7IS9KD5DZggOneWAwOb2FEunw3YE+75QJ400et7wa5LvQVsfc2z
W8pAPsdLbN+0R+XiyvFZgJuRQMs/n3Zv3SuhN7AfOTQXTxenL6OJASmI1/mSOTTDy/3JVBqPhzi0
cYgqacLVvKsrsNUIsdJNgAWy/ZpZwXvEjFaroUYYDI+IhyIXPzR4x97Rqoh+ahIPk6VSDpLd0aeX
uwm7NoSC2bgbV5uU1QDQ8PC/5ipWFJ8Ubbw4t3Susdw2GUICcTsOIIO6hKKof2xPuknOVZpGFzLL
tBpBDgMgjobH0nwerIL273383uwn2Sb3+uU2VoQAsf+hyxBEhtSxbujQl6FhDvhRBILseNejS3OD
bJJcDHiA5g1IjqbbeTTd/XlUMCQt9LCN49AElyBagXgQUOmabL15fYhwMDvGPZ90kI7OUnE/HEk7
s3680t5K4roXYLfEfXooRjpxxfK4CBRLaqseRgau9D/w1qUGiT+lSFhHYFFwlNjRItJngOZiPYGQ
Hpyv8KqiIF4Sp/39yrGJ/eBkVOeSr3LCEoYCQstJIPT0ASk6X3aoH60dcHIsmNlholdbQgmBtHnd
giGt1+pmtNJx6P4M0f+wlVn0T1bnwYfSUDD6zTVhBTKWYSkh/IhQEGIOecZa+KDyBJrXd2TujpN2
sf1uITES6C8a6eQheBbEG+4+OXuDYhWAJWuyJRaFDdwNYFvC4r/fxhliScM4aNzb7yXqjsT6ZU6z
dtevc5k2RQT+7PvDCnsbNolztYlAYvMb41cYU+R4efQWuGd5q5fkUy/7aistdvnZ2sMGW1uKdP5P
4Q0IJRxGWCIfQuaUCg/DO/wBRVJk4AqGxYicQEeAVgLA9xF4s1r2bJRecUrcAj7Geds2+iB/rKlY
K2b8yAHKRZQ/QgIvpAJyLYrO4IFDxFyfuisMsdG052OAoshO4DagjMbW8eDl1yd3ZPEQcctKZmwR
9CWbfSZisDGShL+3SoLLRkQj3aTSQyE1r3XyaL2hWycphFpcagHhYW3WTSHyTuxSkajqlj39zkuW
/AY3NXLsbEmctTbB9X44SnuR8KCqBN7aav/hGyImybRa6nE0ie5Wg1J79y32lsSWVAWvDY2QEXqN
/t1s1UBhZEuuhesGcb54Qxp7nUredjI1S70FUmTY4V7En/F2ylnfUTEKRJZb+dgcbkxL56zaDpyn
4+MZl0FiuK1G7Qcs5ugSzZDml4qfVkDEH7dsNAxyAUAF702A+zP3DZTUT7Zb8p+xccO2o6I1xfE4
J2q/JTg3Y2wgjMhjAPzYZestxc48mMqT5tdlyJyZkUd3MQXCiojYmIy0qph8s96mfhj5jYOjFBVX
C004Z5h9BQ4ZBiT9fizsSzVDcSvMicNOxTHntpR1mrx93G/1MCHKJhDZT6herqMoSQIjjDKl2abq
rItpmFYUGzvbBZXnchK6GYuk38xco1uqjBk09MMWqZzzI0OVkXNG6fSvDX6eNFK4vXPoFwzbwOkZ
QyQZ7Jm7IWXks2T69F2wVY63X0+g6zi/7iqn19pdVVP0KV4CJiXQ/BlKhmsl/K0kgRlSim8jSBZ1
y2sgX7zuwDcDNqUUdg5f2mFCqGCah1zv/+n6GGdwahOTeo3LaZl6FqfuyWC4ppobB65RM1ezqbNl
5/xvPailyLdD81EeZf8uJJxHLPTmNApWdPJy+0+aRDsBxzXIpgHIPdsmvo+NRiHq0IQi7AkzPycY
6athAOiTnOq8L+Shia7CiWULhmq3WGzzrHy1EvKn7yUBg1qze5d7Qm0/7IC5cH1YKW/maTkkI1Dj
QkYIjy0794u/RmPc2Bt0mg5ptdxqWi3MmL36mH5vh3vhYAoUYs7yTff2muveWx50ANqK2nRcmaYD
9Dj81EEbrZOaamFj65wT9yoazTx45AyENixLxWK+H08tJojlZS2CQRi9cJcS9Bp4QN8B2NYJvVAQ
rTrKjKkcywnSH+Xx6pAUOtTg2bnviRAe7KRTkS+4S+uxI3KDPfZEN0sVD9HevZgbgWcVjGi5YX5D
SDNkKd9Cr2imeEi7SqdTZrWPYRL4mJAqL6kPb3LivYMYVgCu8UIvfBho9bNXDmgUQbq/A1qSv88u
vKLyJ3GmBMXdd6Id8mSuFd5ZtvUbhEJSitHqUUZ49r/9Y12oqTNBQaIjxiYoRrsi1OOr0AcstO1q
43SVV/KYGMl+ahF3Hvl4qQio//Gkw8PV6SLuxPvQ2s9HQusPTCZRK3i4lC9dfw4JF5iwlymRyuBT
hdVCy/kz9InVlolPfeWJUVvTY6D7gx+A32jeRQv2xLYrOKTaGlnmA+CKqzgbsfaGS3pMNELg5/p1
Osqy/ZsIcUmh+mloA821B5Nb01loURU3Nio8A7CQ9x16OnQj6/LtmKdcAu2BCgidVgfcHCN03tVO
cZ3kCdKdN4PRLyx4y7BCEN0WrXMnXduFBq2ZfKhW8QEwaR9cLurfRHpaACtwu32bsAR43RUZneMi
8SdKac5fNTGoG0++YhouNW+eoVytMxTvO2hfvE+HeUtezoZu1AnSwsoCin00Z1aYV83Ba9idiRxk
iHJXlcdUlaT7em3lkC2HnGQ9Eyw7tY73aK2+hJSLr8sMrjbkJJD+yvcskZ7CwKjdpzK4SjaxubD/
k2cyvGNv0tX/iiEbxQlu3Z9lJyxxQdMjJl4XPWMmfmoABMFEU//njNSmdyWAcCUpejaEO7rJhBEm
8jFY7jjbD+lLZXn/nyKiMs3z48aEb8a2biteG/y5CJFocQ4MuEiuX4BLnQOcHhf9SznlM/5Kzhjh
QiLuhVwx5+QRx7mPLenvvSrtIA0yZiFmsrlSZBko+9IIbClG8kqgeN21Hz1XX2lHH1vYmnSx5suH
eLTTC7ARurqNVEBZSCMMPJAg3YWMcYm6kd2622LjbWOsufkRMc1kX8KeALIBd4HTZDjxfWTujGRc
iI7qFjJatyA3EE8baOwn58QX92AGz1rGC8wdYZXkxyumAIiUGEQ0dCgGFnNDWyx96Drx4Acjup8x
BMnU9QkknOskBPrElPkpE8LIwGUq7wLZza48EsLPUbf+s5NG2dIRUNGXH5rvzB1uRSE5O8gn6qt5
95vzmbqW8Kpbv5K8zttLKivcyj0bb1n0jqQu7v1e89P5j67/RYkWwNNUVn5tqRcdLhvJImPepO68
UVBagWPb9v+hwKEp1c1sf4nH4WME1ueXyHwAqAwGJLf76loeJ8Ypa1H/sIui5dItty4fNV/vepKV
+SbEqD2ooD3dz2nXPc5cWZkMsrffFdZqrzoWRR4dwgahe8e8nO546JPjM+nL9FADgfM4CYyiD6W2
nfBOO+KJ9qI/Uv6vUvH2RC9zqF/vZnucHST/thWE7rv76iN6G2hXPlLiq9rLNd4DtJwGRUEPdFjd
41bV0oWtljYwDsRrY0k5lIorD2TA/X5gNgHkEaPpMkDfecitTa1qsfY4JmjtOsf3kByYAG8NReS9
kqnOF8d42HQl8JF1vmAgsJD3clN+y7Tk0HHIuT4d4Cu/snZXaNvOwXu7AIrgeQRaKYqrcl8npS42
s3r0PC2Tjc8466th6rmWvC9udlHOLKdlJuWEHTmqqEsQbS2zy9gYH5HNch2NuPNLgf7KGSo3uJRz
8g80IW7iUOwsbQ0TYC/9BnUKdOGALU8/f9hnmRqCb9DRQSItB5tE5uprrUt+amGgwTmjpTznWpPq
N7nRFRa/jF/aTe2Dakm+bxUd2FDhNf8HhxwJTz98fG7SbwR4yQTJyGvkaIZa4pqSMcKvtUpdXG7Z
+9/MFqo4BhCdVjhu8nU7y00MUr/q9htyjqhA/zJCaHsXKWQTEeETLTRoMKUkJBtJ5hdxdHoFfK4S
6GM6w1gV9YbdFl3n0VglU+wX77AL2uQjKi2ef0XGsB9iEsw2mMQOS8izWsj28492/8CdFHDL6r1f
M0XurYEl5UEEuAYGsjR/5BJdPr9MsdYtUECsqilyFjUZSqkhB6xANhSSHzt5RhyI++gNtiZXIAT5
AEqRLoO7yX7S8BTvWmA38DOrJgnWOuLwUD7JLYkJmg7mn+bv0uY/D3WVk5aA9MvfBY0XnReatlve
nqLfLF+cf2AvD7/UPsj1A78Y2xgyrWEq/m/aJ+hd3OHXJGqGRMqJb4mzu/woYisjtUjHQReuipJK
NJc5GOhwbRdgsTZOo3uXEAoCmRcY6Rsyh+4f6rkeRu8NPBl2mvr3VL09HwYf9ebB0Gmrxb71vzzB
xr7TIl8elIPTrCA1XukYqZZ6bc0cwMk1y3ZW9JzUYUzJYkkEVitIssJmlMJ9T4iY0QS1S/9OsfEJ
FoCFahW+D3NdwEoEgaULlVnfqnXMFVwipmvAoyn7QM2zaWgO7/iN5BwkjuOgOLozZDqpEHq+0tdL
a2GNXLtP56RNJjIpVPTCpA9wFUQoLtHoORMxfDpr5NzzLkRRbi+VipJJqZ/VUWTRrUQmiR63a8RX
fV7YZ4WsymhIE3qw5USnZGRZNPYHBmfIBUrDYnKIBJY4rpmpOdsgyqNzapcepueDO/TAuVTXSdB3
jdtDKioNAQX9mALBGawr/SO4NjmaOuSbaTCtSKMCyZXPNnQY5HzxVgt30/9x75/SkV4IjdYynEzK
G3jmU0m7POGID+BTDTimuFQjnrap4qpAIFWM8NLDC0VH2GYB4CLMrfcg5+xItTpnGZs5xxDYmR6l
x4GhN4/vYJuV0WFDFX+59DScm+PNhcvcAlwldASzwm7q9KZ8K1F1m5NCorGFJzCfjejLAs9Mrnig
AOWMhtRrQOwZZAystNsQLAqBmisQlaHfyOvwqnrMxFREf7hlkV7bo2d9e/OXOylIJCyfAb7PnkhN
aeydm+sCVBwPAo4FhVT8/4ppLx9II/YY8EFNNb36LcDczDuokalPBLJ7j+IjbGeo2OfQZcBdGxMI
ffSMLqapTitHo/zbWXHM7Rv0rMHZF4joOMZGTedK4QoQxo7dgTndlmsub+omiNIAI+/5uN5JgdIo
btNBg9l0izkxxyKSODaktbOQ9IfYZPOngzxJ7QloDlwQp1FFHcADvqRcRRzn2snQ+voOeqvcSaQ9
gPgBDBMgTZEqbEXnMqUXTtIlGat8L4tWOcxPPmqQbPCUZaR35YGEhBRsDi6Oa0simq5+j2xAAvQP
NKNbvz3ngyAHchEPc5E3JOglgXN4CY4MgD+ell1PCNV6ZkF5QX8ibMJolIMrjkKDoE/gr6FfDj5K
tKwhpV5uqkOMxzRRCWX4w8Hxxcc7sFohzJG5PH1YelgJS1eGVXhs24pvwA/GZsa7h4Sd2qKrW2NE
HgUPUc3NFMxCrOFXcgECCvz6zC1fBaibWDlyakQ3gz310eEEPHs66K3yu1ZpcMt7dyzaSybP9CeC
1kxmHrBi5rvSn2uXxmtkwYVTZOs3ARFgfktRj40vaGXJKydvq0hm7ZB7VXuDtuJop5xVYSWXIFkR
iVtKMMVEuVm8TaCLj05SzmgI8zCbWw8kztd3ZgqOwzI7rHtwvFCemg1uCrGRwOwBkLWXgRtZTqrm
crKdFdqtsa5s16wsmquSyO9TSycUhTz4IEY7rSOXkjgoGeUQRc+WDAvckmQxIrDQxl2gFeVg83mB
vSfv0KPMCVVQw/cvDAODyPxQlaoslWgkXspsS1GuArHci6x0VMkri1eTCvKOTmrhlVy80JvA2lvV
HyUu6N0baMnsZEtMnP2Tl4BIIUtkUSFgql6858A7XNGe/piVIlH+KoVFywHfA5fRjyqfz2Qz3Bvl
/BrYNVv640wPopAhk5j1r2mYsDTvZ7Aic1SDIATeQz01HkcnA33FELTEc/jpmqZGthMeyFI/865H
nG4zJ8cEoEyO2orFHFtCsEgrshOJLhRBvufMMgnCd09eJbL0/CC5pfJ9gqbPIxdDQgg4EZZb44Hg
zUjgDCI1LH69/v/1hCa7LOPzGIzq1hff9ACQ6qWiyMHvO9Aq7AwEPAFxcMN45ji+EdKZhYH/0LjB
jV4n2/TmXF4XptkguwrsH8sgKke5SOZSjMgsf6ZCk9/aWws+MdyaWIeRKlJBYAIXJujYfBdziv9l
T1JGAogAnjXBABHw6/jOqGYasy9gPfq+RIP39mQLkl4/mqz0PYHkDvXW+rgCEn/5LgI8QVfnBe7b
lokvwcB5gJUBygoauq56By/EEZ99TY/Saf8gkfYuMx/XFvsNVIwFpTbjnpaC3TudWjsYNGsew1w7
XsvcLQlHm2Kw+OYAhrueqKVimctlzRqG/yepedWDRU4tDZ8D8jQy92Up1O+p/56++VJafFWVPr9B
3Tn3WIlTEe5t7EwjnzmeCqj7xsMtIJHKw/gsDeHDdETTqQtZO6qDfAdgza5Odcp3VbXWbJHSbleC
skFmWe1r3vulA6ejMZUmUirAUlJGfpfUFrmL8GoiDUw3sdRcJANVJrDwroajlrhVUEuVkW5n83Sc
IJ4d7Fv4naJmTOQoWniEkO4H/eFYQrRNK1Z4ebfwXx3/yZFPBsLRDHcQtococdBZDDPAZ/m2pzWk
qAnAGburoYmPOJc8p6liPmNC+aB5Ym3q6LevPZowFuCD/Dvkamdqv4EcE7NPtGAg789e0eqc5X5A
OxstQ1pXk1YEeKChBswkpSSHjP6LRELt8oHy85IVzVq/RU/Ki6VNRXlck4FITfUN4NffFF/UThN4
L6jqTZsl7k4TF8EBd1bp9B8djIbd9WF3aWt4ttP+STfQPfoaVgq2D/Ij69DrgqX2g8bjv9Hf/H+L
zgr5snUzeFknBUUe++ms21tHOsDxvF53gO0pM4xsxtB9aX9fe7xrJJ2PLd19pzWA6FDjOeod4fx7
bUeV83m8g6CsbWgh9foR0Pbs/zjmldNMbvZ6Er8ZVdBLEMfZz0Fuo65y13piqMExhUSUzfeFqgu1
Y3jR/9nQwSPFXV25eoSoDL7OUTAD3+2Q8SmGA+g3YdMIeUPTcMSjDYVtLXnyey2nIBq835vaNLuC
Aeqvhebds6c0mVTBQsBX8eED95tGFZmfiXtvZ8LltNEGUlt3wuoCIuCEqpJqLxaaBFq/28U875tz
YOdvVNcYmm2inSbeq+Io5pwq1ct9EWCJZtDvZdhTNgeu31+XvuBAeGaAT0bqSCN0X4aK8a5NbtoS
/iqKEaZX/3sPFjAyxm0H0dRrSYmbXgA+ahCcQNLdzeNptS+HOBqIS+cRFUMDXFK133gkLQrWsfGI
S+BWCbFDWiaKFK6m5DOQe4OfiptxvbrG0pFL7P5i0a2UxrfDc/L36rDDBo2Vdzsv8wfI1G2GduKE
ju8dHjoV8qcolyu/72w5ZRX10RBBBsaRMRYblVQeWpfvHXnGrEbZ3m1pzBVP0koeXVAqyuNZa4o9
XJh1rOK5oClFnQE2A4jEb0ZsxHRFGtdJqe/Uy/6m31LTUWBKG9vKW1yTupDiEVVWqcsUAv1GJOd8
H5nTRnt4nGz3guZuJUsk50pKge365GNMACP5+yzTZDZEgWJW5M+Tnv0QZ3SOtgo9Nhg/qPcsz/Ce
2ch4aJDukYwKM0rJQko6cHTsPSpep/77SmWgE3QbweZJleVd5UJEC0i5iBOphQACah5JNNqBV57u
2VhnToGzG3vGmy6bitG3KQl5IMaes2u0pDTwEfnCemBnWh09P94VPbUcNTcYl9KUs/RdAGPWpwkL
I6ETh1P7cBxCi8cDhluCI3w3nZ2bQQ+Fv54/7DMSGN5BlYSV2oTTNFzlY4wsjKyqvaQ05fAUxh3n
m3ldsrwf3xqbhNdOyFypLIC+ii3bElknO0mfg2gc5r2EbLxW5TX+YhsDpqyiIjMYeAD9aFIXiaXo
EXc0GOrA0tvl63NSDrGdhSpS9yHNorrubbu0VukjWw/UtkssyYtZ6XwTJu3ZS6RIaI8Z5rBCfJaL
G2hG7X9RqlTWFJwtYx8lLnZp5iQk9WJzYNwvUHFchXPZ/1YVlhQa6Ifz1Z3bcrAFjpzFFLodaHcd
D6YJF2hJUWy0xwko7R8UT2erE5Kcl8Pqh1pjk2QeKWNT5UtXuNntAwrM8BGHyUheqMRjgck1yaOj
qIBDP+0iAT48V+HemPhnllC2gxjN9mCHoSPKJ1mf5ZgJ9ExMjgMXEk9RbdEqoyPknHdXeZatUxl5
GuVzpf2RPB7GLlKr3aB9HK/U8MxDZV34FT+VfV/U8V0v0TQs8XbI4TDL4n2Bc8MElhittf/oFil0
Bru4bAkCYwbt2OqA1iusZVDIK/AekQ5w2eZDWvRafjww2QcrpcZLHbAv8DRVHOb41zjcjpwnQD/B
Feaq1N0H7ergbmYzT78hh5XPLCPOAi4eP2NrfU5r1qB6XVhz3vrzF5QgT7MjgLaqlH0gCfnuoUQ6
bCn+A0TGNUjbqDIMw2rMwfPkGx8UHrWTlgjaQ3JIxuctYMGT4wfP2kp3iDIKWHBuS1fFfFht33Lb
pmgYFW4YLR4bZ7r6T1kNMgSfo4CitXOhXT9Dww4C6jKlP6ZXlsMFzBrasbO3XEBtDZdqvwHoos33
HcJPhcQsFREY9zxQqkUZYoFhDkGMEJAmR3ALljJIB5ljZiM0obEOwyhUBJB44w3UAEPOT+HjOlHA
Js5M/8NPEn4s51SffdAZlfPq8Ll3TvAPhnKANsTuiCHsetsq5GBTQ2bof0H/EucXibN5glWxdWvf
oHiAIe2k5iMrUHfrGLfSR4uBdkvfErEsDsIc8+RQdDoWTrpJxNePKM00a2hfD3ijMA35ADKfw8N0
MFXHel3R7J4qvLEFcs/XQB58NxtBYAm5+jVDS7x4fx6z9woIXTKl+RcnUFXkvwRWKB/ox+x5KHKW
AQl5crTJ2eiY0d/ButMEoWCq/c2RJunlJbF6CS+4Ga2ZbeFv+kNXWWEHAH+YcoI07Zt8qbKJhQq/
2jSXHBvLR9lCNiTR6J+u0jdthF6tuk7LtsRc4sai2ha/YfIT7Kti33mfDUkGm6KNzEuHAxk4fPup
oQUFnalwoF95CT+icaexRLq6qA3soWm3lXIWRr7624+SIebJlLPMuik6VeFMfP+NJ5xxFk21JVLM
ZQMbSVKZ7NdgQk2kPnatKpVJy0C+M2pyyxClO+DN+9dw6cqZ6xRAjUiLfrS05BUwcVl+cOiW/DK1
/UYjZ9U8n80Smo7fZJIvsNHl/9wlUOkas40GA+qalVCppyqUF+1KBJShH33FzaYISL6s3VJ0eBXq
89RFhyW4TVrDph3ddL34oZ7rApQ4Z4iX/1tYaxytT/4z1906sJUmyg47cp7Zqe1fNHBDxuW4YAJ5
hQcRjNK+JAGx6NE3eKPQx1SI5FwDQYBuA2wDsfaM/NfV2bGA4SyhIETIx1EzTv7M+xwA7V3QJHY7
AO49eGeoKILkCQlHsjuqJPrtlmy+42oR3DfdLJ9VK7UgMArQoGqXUw07Z2Va/SYaW3mL6ncS8bc+
6aY3iLZWNPJinCTuzSX8LG1VU2ROdPdpeJlBdSlwZ3BS1SgwAkB/Ha57AjNWxfYV0tBhwQXG9eWU
/SXBQRxkqC6Ara0iY+1QwKpxjnSThyk7E/7XQsrsIV5bJid1UuWslXzIl2xLmYzfj6F0kENuEhlI
MLCXd4cIoQ16BVuIErk57i3E3pPNPampYmi+lVvxY74G4h+XYG8EOeaBEe6L5tPtbgngVWB2Pjn+
OiW7UZ4uGkL6CA/B6aidm+oHsZakco5FIlCyceR4dZDYUwEToKkoITcphOxHX7TrbROLYE/bFYS0
h1f8iz6fbqmN7GO3P7fdxbvQSiyZSdwCvmyJcLE2wBuZBrjbGfdBPO1jyEZ/uPX18x5smEOOCPXf
cMkG6XgeYorEITmsmz2vHNK1iIRUhoTQ0j6aRHlAhGCHVS2LNQWTGbAybnnIZ6Cij6V+SQIsUrLr
RxO+aIxd88uN/KZrFNwAUe4LwZaRjUBH/fVEzlWlZ73BaegiJYoQ6vTzSfYNrnBh1EXdyZAxA52T
yh6rdfw1cOxJpWYlhXnXhEjAwkCmvbcrFVPp1/5iUA90zTH2bDlHqzHtvy33QMj1s2tg7/63J0KY
u/aT15zKBSrBd+y9HXLe0f6ab/XamJXt8Hz2sJqOBgiylbT2SWUuy9q68HbpnYHZT3NJIA/AHcZn
FAa8XiYf2N7TIm+c1XObKzFryWF1WZbOiT/yFp+e9Ga0YFsW8AK7LiZSAR4hs2ZdF848myu3IJbY
J8Yzg6cFa9KrR/05lRg5Vpj9ghk5peid9v9FFBDX24VGid0q+6muXm/u70wHe9jcAAm/peKPQw8s
GDw/GLI0e54mXgk6UH8Z/qUb9qlq2Vm2INzBY+rzfWxH6YNFO8jsnQ4Z7wCWjecEXedcsNTRooTG
yTyd37raFp2/7DeBOMI6TksQZh6wM11e64tJULBS5zdtLi9jF6NlwF5oD6k46ywKJN1uHpUwWAWT
D1GK5tPzq361vgaIdZrn+G949br1Ka5kRPIpS32flrNu7a67S2Tiz4JVnnTmhqG3JUPCJf6OsozD
+7jlsfi8oPVhpgKMtg6kF/F7B6st/9Dp09hSxFRyGztqRGZXDEx48T6RkwzrE7Av1J/2H5AkGNZk
Gw4+gRGAo8XwXAyxGF08QTDiuJlcNUxykb+B2ExyjEQlRBiq1oJaDAR29Hk4zrxNHK2yXctUDISz
1Giz0j85dFmVIt8qIGDtNP83+omL2mwR7/VvHF89WDYnk9yH4HPpXdn+CXd4VMY9+05aoZHvG5Ig
cXEXf991RGnbBvNQufsRXFCz/Fq/Jt+2KLTFl707mEiej/tHvckCjlOfY/iReSJXsPkCwnPSuFag
Mj/rGCx8Hslwnhmatcw0esjP4ejfl9UvJPF8JUA/foJh6LgxPFufbNIQKmNEyyd7hT9TsdvQB7ti
ua0iY6jDuBW11QdKTEBilzgpl7W2llMGR2xZHU01w62jlLuk+0+phq+XFofXLWDmxsXYqlw+5P8l
XlKvzCaCNVDlaY18/c+SQpxmW9p3/ycKnaPzkDddTW1q25iZDeGuLpc1u9BJBkF3qgnIYDGzWpZS
9AqJrsaYGMiB7+/r4+g9CxIOJOjsxVBEvmPhu//uAgqevXo8m2DcoD6cYzP1ClDomXSDG+dPWKXz
YFF9Vv8wPnGQjlLvcgkF0DbgYkuDA685M023jVg3eih8ssrL92MswqYAZvHPBeyjAqb3+tvZsI1e
mRNfovQoty6DVerLIKleNT8v0CHkLsts59H8HmGXDiwDyQ6bdsC5bn1BOjSDqkFlK8CQy299kvfW
bjMWoCplgebIbEGSvUF1rtp/xXVq00/fEntsaJFOerNyN/cWlVvYHaP6wyOchFjC8xqaAhGOQqI2
CSsv3Ou4BdQBmbYEqVNi/DwdgoXy35McUsas2vJ366bvDg2lDUxXbcGgvtl6aZro8I0m9anbYCae
bnyZePKFz37urXCWtC9JhDbXvxqGG+mi2nq1lNJJ0k9+E3at4wnRJVURkaSMtAqlcEMqL3WFMwzE
faEY/lZd1hrAxweslktL0WeIc9EgM/gH9DuEgdnv6BaxemmPquIwHMh6B7qR4r44HnqjztFs4y35
qGdu5BmRn/qDYCHKeVtRIEuXTVbgaU2dwmoIH95gXmUPiiWw+CdnSK7X8z+z2K0250evchE1EqRs
DmmrB/YiTw/cFTUR7LJw3oWs2KLLwZm6X2c3zY3Y/ZZOmykOhKDZjoGx5RYf4DgEnvMqo7+LfCwX
nrOIDxfgw94V/WYCpgMpNanPso7NRxOXzyD37NYcYo8fBAqOb3hdyqgQLxCHN3zxHObhdxAcrw7y
ujkUn9/n59zQNJCArJjeWUiY5oMFYqaRyls6LJDhOktXvIhXCJChPVrCgLn5FHAyTgIKgFw9C91c
E9WzDaJKfv+FiJl69MqHvjrznOwuLIEQtclDkA7QwmZpfwhACYrOxbmORXC3Y0K/vXzCHLLTV4Vt
J1NfimtsS5KlSdOUeptYezE4brek8BLQ+gB71neLDPJJasCC/cO/cokEs0qIzXpVYJK/PTAzcPTm
d3p3/HLU7kLBEd6SIKRKRUmK3xbFwyhmqvVLAeGYN+ewtt33PvLXEZrZSCy2n8tewGp5c7JgA+1Q
TaCEz5NpoQsqLTSXaXBBCO1meu43zz/aECfAlDJWv7yepvlTPCJxtxw7vRRbtHuqWfOmztCQnOvu
rvCPszwFbdUGCEKNKwYbNqoHvXPeXXfP+//O5V55tV3W5swL3RyaaAERK5CCZ0Cr4nt1Y6/Sw5Rb
LnBZUvfKkFVgVA5fk0SHRuYd9+AANtVrEy5BJgv3NrYCuTRU7cQr8JsUeghkwCp7sM+TfRpxppty
q9kndwB1/5NnXa38RTzZwW6Fj0V4yVEacJhVIWYGGsNRa/3OswFAz+U2KpieqeahlP3p6ePBOQBR
m9mVVVGNkpQbM+C6fm9/tAlOXktyvFT4j8SELurnMIU+8xw+FK2NdRe1gAwrQ8u7NWiN9MrmrRxv
kQRGXTbKpDg3ZLnvMY7Xk1T0gb4OEKrPu/0OjyR0rExqLXBv87PdjlA1lofBYzmANo/yP9Zpphiv
V5/PAO7EYokIFZecIv+Ksoeb41wgLj5dYLy6uSlnEM5SDwMp13Uo15rhIEMi0hLIGhEhB+KnTex5
KE7V0mprdVBIUj1nZlMgADi10F1zFiOu8FLz1arVU4b7yeQYQvLP9kEjWnYEUEPeoUAYSDmYDeim
zGu1a/0HZ2AWj2mKcCXZOUR4Ob/ERD8oSn+aq1g58/kcmS86E0oMEuFeZ0Mxss5og7DDhpI+7vrA
7g6IB5bJF71vAkroQPDtC6BUgKD9zYJpDhanvw7rrqZoCIXsmvpopJD0A9/NmAJpEGpjfEZcsQFr
XK6po/UEVh0ms2dAxksVJl739xjiz4SJmXChH2QK9gdO43BdxZ23TpTJG9IOzL/NbZaDQy5Zbwc1
V/NSsgj19JNEBEgp/+8MMSHDSqqfjl2lezVN+JgNzAja5km+w98hoEJM2lHuZnB3xtrvmkGHiSFK
YqmdChIgcRTxsIk21Igbgl5EJkthO0I8XFDR1mIk8ko7L/uziiK1ru/WRv9rDXaxHvLZ3G1mhpDX
BC3CQWNLql5dA7aH3xp6LTQyuHeTCjEDB7yvopowOkYJX7i0d+StkVFvIsxIqhauoOghXEDY0WpE
2QKhjWwnRIn2+BaCL6dr/4J/mARMz7Ilpt5xaP3Ai4uQ9lnKgakZ/NLknSeouwBJoWe3nP1A2NLW
c1/qSq8sA6m/MmwD/c3Gs5dT0o0Hya91ZTb9BbvicCi/nmmR4JKzZx8N47wiS6kZphp3Ru7kPmX7
M3Cz6cSVm/OVb05YqXSzO1sOQSy7GOdUHS7vCr5lEl1sGl5R/uiQznsUHPEH4LJEIcwElpSsg7gR
Nv3GPfSB1DmlkwXy+qFMfg61dWjhQK/z+CdlLZlU1xZqMkwsnj+xfisqqNiwMaSJuRntGmiqToTy
TXTYO855TyMfEsy8JwdTGrFXX+iaAK/xaaJ8eBO71mNQAAHiDPhBHEC99Ws1QuktUJXicQIrwlSR
+/3I7KO7er61tvV/xv18+CzgWJhKmlo6NXyNJsgbs9eOVUgejQGVZfFyMKG+TQuVvVuRh/B954/o
3aojxsAhjQJtYvrUOQJNQkIKKS9rs7ToqPXv5OUG3AQJxf9o3+55ffXBNoHBlTyKeUxLcvq7Qieq
NQOd2H74I485Z7OV6JJjAQrPrYj9pX3jZfG0r0jF3TUDI3j+veRSK5QgrGlq9bWGZFQNrdOBUOTy
3dvdpQAb+JSRT4EmvZ65H3qOBvhBv28cG7C41cirbnnAPqc2X/7xM1cyspGzDz5Evf5Si7j7ZZLU
1qC+TmAxRu0o7qfzD0+BT5QaVH/dpzdLnqK/c91sDEnia8URXkwylBgaNMpTk6J89hzCUFcJDSJs
1ke9m2o4ktCM/Oj8K1L9oDTKOMEzzTbIRWeSTc/HGkxrGzpe1JD/929aGpohHr+GQI3O9gWCSYox
UV3Rv02KC9Pk28nH7Xp/+Rfd+OgkzdPMcLBTs/itQaa23KZ0KsspyeSM5kYQGqbRZC/YCT1FUASQ
pe7noqMJPfkWHbIRlsOpTLhPNUYrHHVMB1jIrDYb6WSguF1rQwUyy+eJC9b3ygweDXfms08qu/Y+
PVwrDQaETeWQMnzYdwhoy686K+6F/OcIMsz4O+zo4RcZv7nQu0Udhb8hCeQNKKDFVnVEdym4VZbn
k+MXrUopj1fieRy/k2UakduCYqII229onAf2onWvUVCRuY/zKIGPj3UeSQaKocBG/N49t41hUjWr
D87XLCqPTycdTsMYEYqB5eRn6WDqQ5oBEYWiywqECw6vJnMJpnmFW0iOClJOHHjF3dhAztCNMEpi
gM1V/7Jqo02Q/v4FGKvjR0J+QYGzPzhjOxXrHyGEzD8hTTM9Q9swVbm/TDDLJlHx+bGkhmUFnzVm
1Zdt34JkvDic3SN+Xl8EYe+j1n9Y53lDW9ZORZQyjE0EnTrt+1DSfgtH4ad7CVQItj4wlZV/7ecc
xMCDS/Zs8IxoPD5U4FT7W988iazHU1FWbvzwgSBHoUABBW+sVBFstes+dcnaTqJLse5Q1oUo/NwA
z0OGeKGbhn81oE3xpAryr+nZYIGgps0HsHW8QNxypsPQoi6y8EHlXQgYDa8Fm3HCk+H9NN/aLq2v
EYRH4jAMhpgPVTmhIaU9JT8bgkYsty7iKq6mEP0Hbozq69KOgCxSS4aTySP6TFwMf0l31rIgUAF1
IeevoyecqWE3TYxROVIJvtw1Q9y9+nShYBDCDbQHZ3yLqU+UVnV4+tEB+tYls9mwKcTNsQoV2yiJ
Zcn3Ksux4fS/zAEJkgOWLilWF0eF9PfSUzzWa3c3JWUsCODngHuRCjKdRIakNFxpz71Tq0uSqWXV
/1P2K2j2ExC5UO1q+xhBa2xvsFcO+oa2skiblc5Rru69mzEmX88yWrNETZne1Et6l9vFs2rSVRe+
MoKKczSzvg1IaHM04o3NoHlgxfUm9Bh6Vrw8x7REqi7wNR65opcAxCYa+kr8PZCEXgFCZ2gBLF7W
wgv8E6lJPRR5dRC1FC38yNa+b4DJKcHhH5zHd7JO2lrQjvVUutciTMHys99wXvD0LxULflHcuGfo
+4hkEVprX2LjIf7sv8VFHUbLh2VlqOXT2SkHEW0gBMjuEO+EmZRIQJxLPjE3x1qdwV6zB4MFXBz+
SGAYmNpZImVgeWITaEtIF9U8v5mk9PzYF0PaSUkNsCU/OTudoQhSvB541A9g8ftRJbxNiBAkJzmw
W3gQLESDJDwxCllTn80ef50AIrDB0P7LP3c5KcxETiG1hnpqP3zVgmNzWS/BYfzp4YGeA22RaR+n
iWGqO12rshM7bB2LvCtWcYEfJSQ004X2S6Huw4B+0qt/KcjB2C466Ywh5M0UhTRi3UX+8uf5AnHl
v4r/5r1Lf+JewhQHgSoqrVeAW8m1bK47i/YGCbVeSekz+tmBSC3rRtyqugJqXzc01H56Geccb+MQ
XCBntf3Z6ruBf4IPx8sKfyRE4bJNQfu1vgQKZ2ipBBss3ZrHfvAsAp8KLanRX6OwoQqCAQOtwIhe
0Qu7I4qNJpVILAnExewmkb30lsxPp2Jpr24HFFsPFHea+O8V5bPrBVkjZWXp2uccOfbOrWkvDoyO
cqrNGzAZkiFqAUDD/9tYhceM9swsXSaEP/Um827VMMyn2o+bKPth2CB+VqDyVcNR40SafN2C84IG
i1coBL5w3td31orPjnYDdTIMwqNi1BUTJPVys1AqeG5vwpkvRuGEoWgGw0snDtoECjeWqb+tvx2u
v/5i2OpV+F24UyURNd6oCHhfD+VHECYvfeEBWDl/+ikC/M7UDqp1/XZQCmEOxuwiubFKQsL0J3co
1fr7Q61fRTKTwVoKsCuFwTXVLxnCEV5Z8wXtBb/m8131QpdBUAkI5B2hT3INlgZfbBm/UOPXXBeu
HenncQ1ygUu48ihZ8xXi903MF9v35XMeSpxU7vX8RWXex7r3Z7X5JP9/3O3bUZskeXS8AGnN3OoD
L5aPHzt8Zluz6L2u6Y+BWegGTgM9K1HHq8qonxWYL+d4o0gPilFc+/kDuQZuDtyxc48oVZMBivL6
cMALSTG+G45F7o8hgi+Zef1CGcl4u67NoXYC/HfBFpOtKJvC2zFJyzkHHTNXURibNJAUkjT93fpK
4gdtyp+UQ0tvO0otREmIJnxuehW06lSm9Abuwk+60Sv9r9y484mn0mcKuz7Vmak5VNbYWAi38ZPh
1p2dbtLh6ib5GzEG3OqWO+D/ItfmN4QPjjGD//TznXa2XoeVFSOYzUNcN2HN1rK60movupVbtHJf
R0o0xthQZqDBfpiC1tW3ugI+7NhupJ/A/4/YQeIroGWawHqNygNY6i2R8ANUUBFa0qCIcPedVaqn
y8AiMm3hmOvcujOFgJGPNcMtvYoA/KJmyq6IiEXIJkF1SEf7VDLYNtYc6LP/L3qt3mUpSeD5IAhl
ejJDzqaGeWXcCwlid71MvzLarxGWGjaIRDyvy2xurAZ5//Lj0NQYVcGPGMYA4+hR1UuiwU25Fo9s
FtjxHO2sRt5f6NDFsbRQ1jsPpPuIT4lRSHELHbZ7IDZCOwbD3Bo7+TGk5EwWGSdaEeWJsIxCFcq/
y/rB5UJBF/WikmGtlGIO39p1AZ6JrWqklexCGzt1Wgz/MuIHWyu73cGi2B8KdAHLeq1ZY+efH8UT
1nVlL3+YycE5N6BFETP3W+alHSrqyvzYRFru/EZBVwZydp4GlztjL5S1MDXydIRxCcCWFfaGEjBN
OIJPih+BJs4F+n2R+wRCa+E9ab/zwZQm5R1n9O5JBLXp51RP9QRnAhmpS2fGfdsxHI2a39Pqq7Dt
0ccRdZSTfAMJwX/OZf1uMtvY0gLoVPPQY3kzQMIchdPWaOjPbUztr47hE3tfleZf4XWwMIvO55Yt
5vHTE+S+bprGt2XrKRtlcpFFrVaw7glmDCSHOI1Dk/o1C10CZftUpf3DV57pLsWqCSOs9nYdT9Hh
cqALGhZ+ZjD9UyaWz99U8FVjtNU9OMgT4++1iXFQQjWtntZB/yK6ASxh8FewzRpRHO2Npusmvg3m
ou6SMK+x9fNq17u6DFojxyCIAolL17SvkIBKRRhADkaF+8GoPkY5ujnq1rGCY24VD2IlbTuOtyBf
7Z0MfnHRqBLZyDlp99L8Qz9RQwCQWwtU48TNirmWNJKeuzhq7s8x0wuaQyWf8Yd4I0fIPiN3lDNt
dg6pw35kF33rKIETno2XWQ9r0K3TbfvoRgVAiWXNiGKY70BlaSLpS/nuKnx7AgGIosJKXaIJSdeT
DmHraE0sd5JsK2JKpbkQK+3Nnas8+PpLoZqWAEBWKe9tZatugqJ62Bz1v3ZZUJwCjrTofAGUC+Ll
8djOOI+DxBLVy5QH4uyg9IR4P90W+Bsf0RBt41LFrHOB3Qew/MwQyzsqjo1MCuhNhqjZS/RHjwPs
0sjUaP2IpTLwwCJz7u0m8WPWONvzU3KwGR3OcnSKUPgkv4JM8vYm41hQ4iL1kN3JwgC+Gy4HCnir
Wc0ew9hDHh8vSluLoCTZwvRH8subZsF898QbE+40KQQXJ8eIHYTwf3n513gtbOT8wKvZsdyLR0GT
XrhYZ9zOxsRkbX7p3+EWsvQ8XlcOCsDxq07MDMtl85Ny++bV/xMvr1ws7FPKa6hfCFsxn86WoB4A
pQ0x7rIMhTDdPt7DDQYcoq4qe2fZZEer0ZmqyTYZXPdbT/Vx/BWrUmrPqHT8BB2N6CdfP2U7Im47
Z/CKW00yp9uh0p0VKn4POlmCDzwqbCZKfDq7zrx1UDpFcgIlZUWHphnwIu9AmkPQ/3sZOh0wi9nn
VHUkv81PtIsxQzD8c2rwhWDz92syxygn4pq6yJ6sitZ5LofuXyqv9znq7YD+ZFjufFmvMn2FJ0AE
+siPiIYyYale4Uo6GJJ69S/GyyiRuIKSyOf8C3/dvpuUUCA/wrL1wSde/VrxOWo6BpFH+XUHkSWX
GxbOwGFH+ig5VGTwbOlTcqRHc8d11gCqtT95zgjQg7ax8rRBcaiayO7MNRMywZaKqBqoJaQn9ZZ1
6wUj9TJbqzttWklJUjOwHGiPKRVqlkEqOGbVADO+SHtPz0Jnyxmm3fzIURQob5xZBRjyswxk2eM+
aBV3uAf+r92AlvkYyTfGpvpT5/tsJj60nWeVwkSBImlHT7rrzITfueCzPyDp+zzcRTZp6eINl2PZ
JzBXqQigwH85e+a9Uf0L/VrGQlg2ZYR9csx1i0+KtURMTnzjtJEU0dbj5cs7L5rYc9paQZt5C/Nt
SK7/umFglJd3AMFDG/x22TkbBHbbdO2PfQUG2qmajr85raVYl36fdIT1A4We14MRVJSzrHdSQMfK
8C3HIt7WbtDckXLyJ7YfBatOMp278kAL7pv9d0CAOrur4oeHQKoVIiTrkFbk2wuqgzzlGSBjNifF
NSuE44+85NwIpaV1U8SnnzjOUd7nULcdLdcWDKFhbEMHTHg+3MV3ajRXbXsMfxgdVLabaicHpgK3
nwGJbY2ItmCWwDvivd0DPT9XQA3dF32aTogHVcHGcKJwrPpQhWXWX2r9i4GRo0YT+nrbktxAAeyx
cVuI4cnIo24yofRXm0hWNxmYFyd1r/ia6778K+8snwi+dpHnbQqkVVeAbRiNLK2W0w+mn/SuCfQ/
aO4ROzvqwCvK0rriCDDsFiK4z84E9qQpWlWuQKj+RYCuwqaRYlN+Vs/57SL5yqWB0SPVnBysb9oV
3FJhVA7CyQ2RvBpOzZSctuSxCUbfNmq3f5Vf/q2q4pbODwot94aGcJZx5cJCoi+R0ajMLkjPkxnk
5M0F/TzydcfvcResCasgqvWUEqN3JGqL2qCOcqIXqd4uesT530I6udGOaZ0Id9vQ6Y0+Z1oCML48
RubiaDYOyfXM+NSC5da8ffMIEgmZJq5GCcw8mvODktKPihbTTn8rP1HOVmnOoqnix2lgtCuPAwqq
G80FdSkMP9rwGKQi3keOfe4oga3ATs+sLSqR0ARTIsQb0YcECwOaxZibjQhjwxhi1NVKFUCaFmBx
pZE6fOPGyrLIcfKvFlAHYvP4oGW6bmsZ2xcURWwJDxk+mVjkXBpgdZfHuZTjBXhCmoYefhWn74e/
740Bwp0YvYsFn0ia3inrRkLR0ZLsoHQA9CTsOr/qv7u/7257gLcaR2kc15FHv8D8B3D3tqtm6QB1
ecVSLx5WohbQSWiUx+I9nDlftoppRhZ5OAw3R4lFXGGno3TpoCLPJM8prjHw7gyjgZ+2bh3J5Qmi
Mi7KNdhDPLs0jmU67Bhfxte7MR1Usbt/m0F+pbr2Ch2+NuDhv5ed+swHt7urPai4bp3alVu+rK3Q
6B1r7TblcV5dAdYbokcOm+3OTp17SL85UX51la5O2ZUloZLm+I2+3WQgdmZ0nSK3yT2eRg2uF5kf
klMIKvxudAKAWLgUaJo0FP4Z+Comw0w0Wu8mgI2iQQ2rZndzOJEoywsPUdG2Und76PtzmeZ6BCN2
+txAXiucO9w/wpvpqiyd8mxES1T/NMWkC0PTJDSy6pUq25REQ7Nekq6NVcGR8t94STItBY220yk0
/Q/vKT1zP2lhHW/Qf6xVtcgyev16eM3Lg96Rv0SXquA3vYJ0XMGSZBVKeiFMuVt3YGXSmd0arKVd
84IxqUTW/JpIolw5m+ZbwdkzLe+8QuHBPm9vNCHBgbbwCGcMDOazFVIDYnXpXJlQhrcUpEHqdUQ8
srJA+Ub4kdug4QJK8xQNAzW/9cXKW7LBCEW3CWOdHgIEFnLbc/3V15QZbX+F3d5HcnYXYdoBRqeg
Yb4X9dEVEo15suqb/xOJVp31I0kZ7RaC+nLRWmIEN0/b1YyqhdjZwtG1vrxSJTtoqx8yKuIbTck5
rUEt4b91th8BS37X0yB+jtAhcR5FGiwRh02XK05VC+KhRz2kHTlTDc4nV8GAlGTJsTAyIaASz/th
eLH+98T3XtpNfIpAT9ORECDTXmk8RbiKs51rHq7K9rIskyD7EXsePHsmoETW+2NklTwAOk5I3Apv
AfanziOgfHz9ZgWcGRwQYnAprGnVSn0F+FdiWECTwr0wGGh1WLX5a1DuqYe+z36NMMw0tPHR1f2d
uPpn6XLRzBGH15uKnWgwm6bsLD+o3v+6ZURV+oQ0wO5NQDXfRv4vLaa+2AZora3N1KnEz1uORC4I
dCYolFA0KE+XCyLasbl1L1wHB0gDn3dIYuR9/k0Ghsi8PB4GXsIhrOaGbQQ1Y8t8H/nurqq/td/z
Mf7n7URFn/ocUmgRNsUI22QbVBx2BbcEHpC07oHWQZs0GfTBWeOuluuNiPD1CyCm01ZZbCxmKukl
4xo2H/b2cwb8C6od6eH771f8pGXP3jcHYXhyzPDzdLfUauGDwx7SRTJFEq2KUVsYefXwSMZnZ1ur
0BsihtYk4E0BkrCC+fwj2NW5A9zY40xRMm1HPSellR4K9uvqjWwDVAg2SqTq4gViv5AL/X6o8Tr/
8TdojjTsVlfmsnjO22gBFYbBXRbObAT4F5zaQeQhPkyLF2WMzT2fzbCpk6TlOqRr8qe4CKfCg71H
wJbi6zTjrYSR3gwUg+yPgFhDeRwa/ObGnM53/vFoFXl5e6cFGxUGe+KBGGfw/zsziNOCL7PX1PZp
dFLTbSnmiXwD0vPDnVDaqoh9pJP6xdsX1y0J1Bebw2khj1NqJkP/ci8OlyNXJHnyixYDlMNlUzC8
ZQ9qUFUDKPOaFiigoybnCfH0OwN8T2v5mfBbrklf38u2fik5GOvy5wUok2fSuBIUmWxVuDI24JpN
5NO/BT+CR8Z0ddc8696Bq16uECCZHeCJ4WDLWoamy+MRhl26bCu0l10JgpahX74DGJV57kAdjvhU
I/x9Uuc8W7HMTuz9PmRo7O3PqIB93Ulb3oVoPH7LCyZQIhmAibE9FFRf/swNWmE9Nx6B7Bmj47Pa
DKccVvs8RI5XBhMEBsOhnjUj/2UjxXyjhBiLwl+D8V+Ndru7tWnUOEnrdZQFtDVFl8yob8InTwU4
2AMPmSRKjm3jCRFr3BnG0p0HXMf8XHz+q8Q3iAlXI+K4DBZaZaihSEtuw5sNVGL4y+f0NJhF3AO4
OMGSTXFF5Fm7gBhYjtW5YLBmcG+gYl5gZUYXgpE3QDYx51nG8Da5I64z2jPjjjitfn0DsL1fF0OW
61p5fjy52uUlnCMbGJSTXun22pLA7Gjjty22fd+cd0vRMXAP4Jf1S7lmgQMHa+SLzFaun1m8I1Qg
OH9t13o3YYyPoQfaPmos4MbsGOul12feA57DcCbXrTa4SvZAR9cxAD39rB4Ng2MvCwdHypCh00Sz
OHVGYS/+vJhhrX/wPMfr1KVlb5c6mabX2oHKhgI0qlYleJKWeMxfY+oKeIytxZPi6otsNqkIyU+O
V1HwZOJhpuYh7EW/Ld14pAawVMl41o6zz7ct8gI/5wz6l0rrU561vDm/d5vCBWK1Wia/Koksq7su
FDV90CPI7hJ+RSzGpF5j0LpLeXp/tYShFomcYjFHR2+xdyLJ3BrLZk9QeB2OWZe45yNAbl678/Mz
JaEL7wuNn+4h8e8jq4JVpqcL4tz7Qd7a6/5yskQYKNtjfnpwSRVCW2AMFcajKvZs1OfTOTt6FDsd
Vb/DiqXZmVnqCYWoK9Dm26AsDiFDxZ3QqHndqZO3L5P1xJzxAOweVjoyonDZpuDn8Rgp9QocJHhC
21XdTDdvJ07YE2+EvCz89AzjvuGZP7j5oAHdG8jEQbo7tMmEFgTIWRTKDKfuzfgJ1+4+gNyOXHmY
vKSDt7UJSOtm9YvyZHqE+rQ03BTFE1fBgeUj2XaQMwJLJN5FO+1pvgJuZ4YOSHHAzHviY+iiolFv
GQhZ4U6dqJnpyzjE88lo8fOKyWq1TjBo78PMb3DvPlSLOsU2DTzWC+32HecqmlAdaeXZb8+F3632
0pz5pt5MUOrI6HLgEWaXFLloRtJLhA2URe7UVZJdnMhU2Va/igLeOnLy31YR9bpOZHx8ECqquA7b
UCPLJ+PxFdFORJlfWxrPx9IVEwHSkSKIkikDr0fcb2JoFZIwP2CZYjllVjoX8AG+EQuh4P0xK0Z8
uW6UqSmOPd7v1dOIsQA62qTYISgRbJXToMrr7NdxB3wAmFuxgjF5I/8crTeNlLsAufla6DCQqlZW
KInOFZ23uUB+AmdcRh23wM87yQYQKUtGTEh0JRfcVoa2BvJLnJaCMMretQJ0fryokTMaY9N1mCCA
nzN6oByay2ElToeVrIiXOxt5DWLnDPD7RKXnrJfHeEhxllKTUGwtZLq6gNjlAHZIfn5e1b2MZPhP
Vbthwg4LLEQhQ7ap1xO/87wbScrxy/9ypaYrjRQYZBHL7NVzfH1xf7gh1y6wpWK+twCxZzXJdVl/
ozI/R9bMpnJDWyS4t58sHiTJEy70Ym5m2NZ9aeqkKQizroynnoykcXvRFm3K0RhVJUO7eS2kVlbU
0FAg4gQMs38u4EEVdAmBiMSHlSiF9TNskYgUQlOSONUuGsFMHIrpHCej2e7AaAbww6gpjrihGaT/
ZTNly83D2VAxAdWUc99fH9hJPKB8DgYODlfZTncZ8AegPF4PifxTavceDTnngLdgg2HeeO42fGl6
GuMVTqVuw5Q+UZZXkLARBcTg/kcQfRa+HIMWbuAjdXP0cZ6t5nDZgr2lIx3taiDjQ7zEl9ehVdU/
UB24vjI/vjl6CUV+gilzN7fl+prR7/+fTtHvyBECVnv+zTv2EF79DPWJXEPgCNiQRv2HSjQLTpi2
sr5QlFIIWIwZmFQzwlYbtqKGxXI66tSUGqQgDJWtxBfNje2k/KPHb3JZqCwjONye1yoRUxELOS3B
Ge5R1viX/YtRfH9euGsxf3q6zdxpYeJKxQjjMUCw25H0yGIkHIOwoHgaHAiLB7yBAuUx15QCL1ir
Olc+dcKgQ4NZ/BhW7ASADF8ApLozlJ881ldHf2pYQyZmCICcMQh5iEUh8USoTf/DW7kxbQk7gDLL
zTJZMVJ+XvhsahogUr9d5MwrePEaP6Py1hDiLcGTHdinJQS4qE9f1fUdRtdDMKD5cdDCf07tLzVf
wKay7ktSA+nv0t7XHIW9FFCO8Um+bFthGGTTcEVR79ICcZWwimmz6YVGmnOb1K/g6/hDsxJvwnMT
4EfuEkBC+F6lpNtT5VcgsAxHqT8/i03SPPDd+7TuXzKOq282Bne+P36zgxaGKMMpt7Qz9MhouZIE
szzChrTJbDleeioJ+gDWheBYEt0oZ7w+rfu+6EDzs/vA6NPc9NaJasyPvEfPx4O1UFfkef5oKbxz
S6uXAYCOi3tAvBeHWOBNKlCxvBwht/0NoCs1w1gMs3mB2SEg87uZJF+18J/bVlmRs+mFSEiKysfp
YbsBfGGyv9zmIWP8mFOja+OIYAcmRRdFn+LiE65+msQ9mHIjeDXtZBPJWRqu9sFwaEKmbU81QJj1
/8qixk/QH45yAgfbRwRzeAtn1e2uBlI2bu+i2nCj5lrTf2r5DOsMp2HZiMhNKdsOP14uPZbulfxT
2Ybf7njbpSGDtYo/pfDhfqSPfN3LU30sJZ4WjQVtMRrAAG27ZIo6xfNdbW02YEfTF+Cuj0EXtCXh
t4hcaCsOxg2vV0JN56ZYVIWx0AxZAfoBhi5M6Mwd5PIBD6Eg4aLc+qFYLE/XA6f1yM+2X/v7whZl
yYOqvdYNrty1ELUR+coYUXJJQYUNkOb6hUJQFK0JIS19ktUPwLbHXXrVGlUESwAA5gN5fbmbv+RU
k4d8Pygl9xyYfvX5ieKgo8bBk7TFw8D9MEbUVws6AEkEo5CunwIQ6QD/nI4zyKduf2/zG/RlFP/n
zinwM3kFn3uwW9c2VXJ4B53Cnip3M9oXhbQ7J4dzuFOZnPjNtsd5+2qdT+9r2P83ApTgy2fWJz5o
VjjnA6TH2LBO62OTLy2xyXUThaqQN+aXkG9xHyvf+6WEHN8wKRjy9Oyph9Gq0TK0umQd5ZhWNomh
u1ASUR4RbRDZlT4zS1xrSwBhAL9O6x6BB/tf9uWBMAaVR+eXBfSSi0JSaicWLFtesoijmTXkrEUB
3+F7WbeJoez+97rT1BlXVXUCPhm6Vv0EePj3Kh1b3LSKGevMW8xTuBsQB8QQXBfuNL8n5r1nkBMM
A3cw9JK9Ny63xK6Qkd53URxduQ83NDV7/FKEFFGsn9tgf1AIEJoElFYYUs/N1E3ofALO7eeCCCM8
c/JNvzCXkdj1DDIa3vnPF0iSiynTvuULDU3ClkEVfRLLtyOCK86NyUw7RnszqNctXlT/vBa5sD5x
4uhDdoFMfw1Pinokeu9G3huqNYxgnOcbc5/KCPfyC0iSTY0lc/vivuj4LV4XlDEwktLV5Zq+bWfA
mvu4cVcqLIkf+njSJOMa15Tw9p6wzJCy/8EL99naQp4dlQSywk3bQCJRMiYcWffY3IW+QwhaArUH
OVXpb3WEwbMWHlmIBG5V+TigQgBDS9mGQVOTbvg7Rp+mSnhRcxvgo3XIEYlA2pLJc3gruzyRfDfz
W8u2Gt5IzW+bGEyzYa4e7uMb9uVr5jBcZ5OsJagt0Nb7HT66vKvdnVL6I+hpK3pnWwxZpqBRBes7
DE4dS0dOeXNWfANp6lilDdXAwKdtff7VMh4poS+VwYSBh0DE8XF2R531d3ROLYu2VDyqr0a9QyyC
EcOm6Z1k4W8fv1vJ2afr6IQj0wjkW1/dV98AAkPtxrsUpmLw89dTRV0HECwfeMlLw3rs6UZL/AeC
3ZcX4VK1EzucBT+OS7ilCHzgQc3wUxqKpP3dSvrc+0SZleFUKul0MboevOJUBRbIv8AmHg6CMEng
3WYXjyk2wVwN+06ZN0KwSzYhaJRpNQqIMSlODBPIg7k7dmgKe5fYTQ9ks12uvHbP3rh72x35HQVU
jt90xPhuFpex+WswiakKloCPquPSRX9apTL4PLHHKEm1SNuM3ofvtz4lbEFN0G7VpFR5prdjev5p
7zVdqs5ctF9kiieAkUIqLdM25INfOlUCvcF+ql/08E263XmNUCTM/wBB1GdDoISziruXxxqr9v6I
XhfuPm8mCg9qrpweMKAh0qWWcsOQWGyI7Pbouls7JJs0cKbe4yctuH65nBuoZIisOnoq8dsWWdsS
EEeXk2UEr/ihtAu6q/blMzt/ruOubcjV3kMVeYiI1sNIGPSvaP12UQmvvJrT5Fjq/CbyGOtFRBBS
Tx2Qjwfl52AQ5BBeKLhgPeZ0IY7l8mZDxF92q12QIp1+sRlPPd0s7hGuDM7ddp2ylaPVrzL38EL2
bd0TVVHTW7f6nSQ8a7wVLvc4VV2AiHwJbYZylFo/O9xleqRdpZWyicugSydzna0XWe6lAd59H3Uj
d3VX1zVHPsSHhILXBI6fwWyBWlXkvElOula0R0Co7xffBMsWKAK33FMQmXPUXtm2htg1j9Bwl4Zy
SCuY1nyD1VW3yCAeXRK7GGEx6MuWO2Jtcxd6sdWkUQMPvDPPFUgWqT1U55AVTdg3ZI0ZRmdsKcUh
qyrlvnkiwismiXYEuEGhQQgTpIgaPh/3gQs37jHVMootzPPWXDVzopOsHAh0whoiLIFrUzOgSsrw
daJxQLvV9WcOOQmeOkwKvKxgL5FFEHMfIIv90kdcvBtsUZJKYq0IWeM++7L9AwjP9+mSdk1t3EOS
iY1xPWjfbIZr+SpIvbtKBnUlCATkTtgljm+1dW9o0Xu8QR8DcfPNlAkEx4pWXPvKd40sNtC67ieR
uR1nlnZFLcxoHHSlz3MyEdl8UV/pBVrkYBiDOlQEMJnUTkx9J0Z0sszrAfhwYXjhsir2tJu1Bnet
oTnxsv4NBaA1i1pKgfabLD6VD5xbIZ0TGP96p7TU2RPip7scIvr5a3j6Yy7OUd1veXSukFJvIWxe
86wHCj6w7JTFOU2tANcbwSB8zNtjAcW5oyC6E2cK1SwWDxjgFN9o5XewaKwFmYCyNvcN5wSRIg5q
ePNpBssMGrVwBKL/RQzug5ukyjIaUZPso3X0dZEC4bqBT8tEv6pdTjssEagFl8shcnH/JbWcv2tp
nq/QU+9WtXZwWfMFRAPSR9q5666O7pA7lYN9jVliIxXtO68eJ5hqRz2N2mXEgAvRnu1P5IVOONID
xne0QxR1dTP2+rynqNbDGyOpyUr5AjjztKr+/WNd2an1dKYHXdh6Aonpf8uh19+MLw7tVJXjnukL
GDlaWZ2jY43tQajXS0JWEuQ96NjcSbIy7nH/VRUCBgpinsTrvcHSZxjZD9yOPCLdSo07YZOEK8ul
gZrByyIv8pfRqBB7kuDPXOdEgX+0tDdVxy2QK4dSTFaUJVSM21ELXxRKtwKsmCKIfU/6H80Ktmhx
EHeCLODQ8yPRdfFtMGqI/ODh4H89L+h5Z23+9CK1CBOAOsNEC2tO3sbAr9SZxF9mstU3RYFUmme/
UKg3tcTZQgBosPD8KRiNnxAhLf6WpNBhMRu/mkiHVWl2eBPu6eYNYGmw+qaQk2X8uq7oJxVjolG8
XwU+3Yw6ztjTMewtIkUd442DhRXF7vfT7KvJPn15xwdBqowlYTRZebFD5j7kobf8FxB6cIkOwU3P
7tz5iABBpKw8143HCWJK54UXsYXxZpMS6Kxg9pgAiso6kxx3+dtD3zcGOSYzUalUbFUP0kTXzTn+
OZ4VgWytNCHS3y+qzhqgUEHq8rQVAsxLooyQ9HTsLfKXCu0dJTTOFSPacTTj+KgcCCeMxirblvC0
SqBRsYgtgtwZUWA1Zn7uvHwtgNjrK+WijssJxS1hFAD5cm+/evkHwNySld/stxriDVySAo5etUZz
tWrrkY/s579U+E06UtUayZGtzNyGDcBtqZcaiHowfoh5GTBY+jNS9+ghbA39hrir99HTCigRfeHa
D28Y/oZC1ZAwx6W+U74KTbmasoc6pNSl51rC0ZDrqZUAcUnnrOt0HqGfXaa0XBdhkOXWh+teehQq
q2uUzaLSzf8z34SLWNtuEc+iRxW52FlCZPb88eGH1plr26d/e+YoC2zUJmEaestvXrhLqe+S8t4P
Xp4DBVgEzrOBpOlripGf2GmH2L7B/pIzBAu3Yni+q4f0SPfcNpJcUFi+9CmOVpPYFs+Dzd7lxZQP
Et9JZP5YUNsNlGVIHW/MVbTsEbEBGmFFSOc5rVdqYpbgKVHPW/tUQwRriiWcnHUsp/Y1iS5UMb/P
HUT2VPmeEbO6gLr6LzEeXnn1h4pTW0897vipSgPuKCdBpXiTsjfTt4EHpW3aJrQUx/epCLrvQ2Aj
8BtZnxrISIx8N50Av5EWZF45MirDKzyQk6XuEPRcuOpI/TEygvcBmhojRNdtSab6MZAgAwHpwu5G
m7hBcZzQEZi+yXs7EVFZxA2y57kDCb5JJuigJ2+arSLFt/sea38GM8KyU+LU4Fn93kTRBYLuuWpL
k9E0ELINIQ8PKpQG2yaALPY4qarRplijcBW9duWvTf8lvGp3JJaCZesmrcY5h4WdmbFsmQ8TumY/
4vLj7qrRJaOCrCjiZIlpEzp3aF6tzrYtscQoEVR4VB49BJkbznZ5FMh2mieCMFwAUJ266GPl09ZM
GcqHvFyqBl7nrP+2wvXUqxG12iJSmoHiCnpQn5Rxhq7wIgfs2MxV4nYH/06SWdZcEx0DsvDGsqcv
cfxrr/evVtXzTpxSqUO3wDknSt7tAip3sSDI9Zlq0T3YSCICpVJaKmm+lhnIBYxdmtsuWLiTZvo4
cR1KWPc/aQgJWHX8eesEs9n5ws6ZVQQ2jhVkjQlGQCt7//dFB8oqcPK0FdPOwiu98ved0ivOECSb
ruL5w+ANLEJnGicfGJDwE+bN83UDRUvM+MPbls62xOT7feOJ+H6unrG4raKm9Ffh0kUuq/uFLdQv
OGCdUfjNDkCDQqOYq571pP7omBgHE6eRIVdjBJ/k6xSwU/zp8n2y8f/y39ERSZPT3xO92OvFrYSU
O7TRspTX8vhVrk0RPXTUcU2bxGOG9AqJ5X4cWCMGVJaUT/tq/3qMGbWwH9JToMlR4tv3MxgZqIVR
pk50u34a0dIU7M6tOF/6dQG9YXqB+5IMRjLR6e4PbtfNtbx0mJ+QedrOwy9gYTluVIkDpsU9Flxb
xkdmAc20jCpEcvL9jhX0xw9PmVPq8uHJlNDtYC9QqU6o7RCdNVIkQE9giX8PooP+8PqrmShDikSk
0joBcnGAYGyerBHAKIM1W+I9mpHMC07CaHgXRXcTcY71weMzaK1mJYXbBdslmj7XJiBl/4Oc7Iur
0IFJPYz9YHYCnjZqUDhAhDdw2Qa4HZEJQPCiK2AP9Iy+y7C0kHVGYAJu6ZTn7m906GAxJNqXgGVy
8/9HT7h0rv9yZX97sbRbFqxEluCJBdGzRnlLfdAfZbfCIHmAsxlYJTu/CPJCy21feS08S7vSVfV5
0yHkKjvThBEeO2COjsaPGHaxFkfFoeYxLoYxozUxVejm6inJRhmtDGEG9gMZuiSsG9PrN9dynOIB
//9PqqJv7C/017VPJK6DQ+Mq5esEbZ9qa52ktT3bDA0VGJVZj9hG8IafY3I0q7BdY5yHhQlrzFb3
HcWdIeMNpkPhxFEiVNJWL0ByAWURvxtT9V3N8logzALhrm0+rc1y0y+zuP5IenocW+oDuEhbJQp7
D5s229/sndGfbmIyzYZ7KrS4joYuTGf/tHBOh4/mounyOLJ/LBeTT83Rtb1yG4v1jMCcMaTUMfbJ
PVyg085/40xZ3CqpUKI2EIOmaAz2vwNMqFHbzl4xW5K2r+rOQJFc+o1yV8BS5WlNLa2ATUBy+ZUi
aKGMOtKJxGFaQijEHMEmengNPmBUwPUWHbBdu5qN9Yn79j/Jhxqwczp49jltYkD+qVGNiUxhngYP
ipXENMhsPm4F3LuIo3tBbh2vEAiA4V5l1p7b+57OXPZBUfy3b2dIT9Hr9oNaNVKWHRcYRxCZ8+KF
6Rv4XZlnmGZWwcFhx73kLQReWM/l5kQTU6Z5jINE3KyDUitLd0dn6MV4fuJNSUSPTy7OhOfXTv/7
ryBfDb5ELa03P5EMiyKfW4+JBGavPbmsfu2f6ZbFFMt/yzIqWLEqJSRy2Q85qSxUksBPsde4ta8n
FgboY+OyXjuYvmOrxmhqSU93+C0UU6vki5t+TxZzydUd9By1ZA2GgzIXNCv7+gbvVeRjT7GdOYMI
guM9ZXdkNNb5S8R0RDLNQMJJ/RN9M7Vp/fm1JBrHZjRz/IL32D3tL6Si18CPNlRjuDhY/XsHht8h
3H88nxttmhTkTE998UcfMVqmdubuK+K5E5QVnt//x7NeH0W1v0r9pfsI+5fpW2I3m0x8A8G1gebz
/q3OhKk4x3nUE7B2XcRGl6lrIBmTtv0tr4xzFoCMOYm/ElGJ9IzWJX8lkcb4WoODKa63GW4Qcvef
JN5URfcjRgEasKN6ZhwxElakq5kvsicDqNaLoS541+n0/ttbrvBfP+gWbUHVQ+YlWikB0friXVXe
xXobs/VuUbyRFLc6QFSNAfCW2LJpkWdSttogggOpFGad8V9HtOCToZxOkrRJrK/PcS03Ock8npFb
eU9rxuQ2dYRHaXOUibYUkokUbgRJTcZxaSw9T7Nl33l+TnJccKE5FWO2O+bgiIXuh97NhmMWipMq
mnTwlTDeK0l0yKnmc19jXaSX7g+gvehzRacSWVqrOtSxZ5uLYyN/fwGopUprqgKQWW1pifqBMmtT
FLcZcXd7RMDTEtyuWeNIcGPV6dD5dvDleNjkUESaAsXWte/iXNvCe3WVcE2+BE6W7LCNNFP9q76H
3AS9puwhKoFTktrQV1GthIDELZw6sc+Q+D2r8muDKXbd9kzSdMkfwTBOHhF8efdblLbB/2tz/T9v
FI+E3ntWgEevJ5hQ2g7uU29JT2a+T8PwVu9hXDwYmYp1CeLb1jtlhJ1AoIb0NtJOQ3P8Zpu3Dy6K
zHOhzVS2imSb0KDkN9CNUxdqkbzKkG5c5uxIF9Eg4nk4aKHIb6SioTzKlJeM/B6avgIpXcYjs5QJ
/hLRnIshCujKXYexT3dfKbYlvjNJ8ZTxj+4Jqd4ZDKdImqyo0C3qIoVzGwoV2hU/MWwRFm0Y1AVM
ZFIT/fsHzIiPktnuJFo2RyKx815T4WhGkKNlssmPs9dQxjJMKxzCE+ky8+6r/IstgTxKpOjczDKD
8//qaH1JFmrhdj7JG1NhZqdtvUlCPnycivENbmuSreZj0Rotz7f34YrCwfHAl7Oi7iKBTSYKRl7z
Ouv2J4CnhOLjxW8EMdSR0rXstxTmDZtJGIThRO3z9QLbA0356SBPbPFM3+S0jj4ET0rln7SVznu5
pfiBZiUgQkSmsnAE3Q+cxG7BGQrqmpnin9fA8QBZR/XkHTDUUEpu4VvnV+t1kVV+jDmvDaOmF0oP
Qrt/nl4rYtjAhZBIAZMvXwmVnXJDmAEHseNRIRdS8hJtQuPv69b2lMGr8qTWRNm5eLJPceUycfKo
BRM4YPfpKrDHK+lJsBKVr2kiSty1AqiwzHX/UyakeOYZZfy5oK7+qPFYaiYlYMqQuV95Cenf4RVI
1syhJzqBXebimO94ChlEmzfcQ5/W27yp6OfCiSETv2Y5MJeHclpK9PatTAp1qhSsow+ZQhGJmEes
htksuz/fXI50z1RybWATqzQASwxlGipguB6wF4bHFSwTcZ65DDR0y/nWSktZ3F+n2GcGZ6hFOxbo
gGWkkXPdF0ExxF8INujLe7Vv1kdokl8+rZXoArw/vr3izuNOG98BMtFYiHeLCDl4AHex9491XgDU
O4pyUjNGG8QOJ9tdA0HDFHHAAai8VcWQhz8bSRpHE2boqFs+Uw5Y2N4olgopRFN9Xc1F/W1/fqNK
U4ODA7COWbEmDRgXH1O8C6eJv9JhP3kZEHl+14m0YwSPS9U5rKiVPqY+v5Vc0FNkAAggetFQFcdA
4IJlECYTSPK82x3K1AHcbXDZZfeNg6Jh4X3LQX18adHMeSPqexY+VSCYJBVVEM3II6Cs0Bee/pWI
GdmYGZPXbVUvjMKJEhvDcMMpvjU76XYPy+Q9JHGT1NAo5zjFhUGyl/afvNIgwAWxeCV+NNSSziEL
v34JWmswnIxabYMnlAlnheK2nYNEIXJHv86rE/5vfucje8RH7rdHJnORujXoYYsZo4MWhUtvs2pR
ujoBkN8uNEKyOU4NMuU5nhBAPOT1uvQf5QZQ5eRBjqmY7MKl2PBYYF4VW8DGaZeYS4q0XXWnAKXF
9QSla+ARS5ffJmFVZjLVh4TT4/GXogdX0oVfT5o52e5Ha7fBZZPUe27i2vAVimcqfzwUoulggOOm
ehIO6YLEpgxKtKtbTgRPWddT5ZYf17YQT+3GB6sNia9QFwyXbArb7mqAsIWQf3REDEKWGgT7P3AF
XoWAMw6jze07HQyFmnhnEVjp4g6pSTeA/cGN+G/Vs/5cJH5qvFZDRKsMxe27eaINN4ha9hcFaCba
QMOD3zf18XugdKIH+H5O5Zl4kSyIYIwk4BWmro05b6RHmUbz+gnz4N3rCg6yIFin8s3+ZqnpRBh2
0hxxrY0BNK/ncwSEnFNjVGI85iTKTKvvhGU+Ng02PcwDmbjdZSJiXFu80VIg6BVlCmiq88t/kvNl
A8ckrEG78xn1vNB5ASTLQQIPMggJqV8uSiELx2om9McGbrue8Z+mLhLlGRi/v4o2gM5zH6CZbiRl
9tO5A5OZZS15u7P9XUOsZPWE1nCJXybPiaXf7B5NqFOyWW8zFEfJ2JD80/RFxAMwvvZ0dJrV+tu7
VYlZfP60D21OobaV0ErGKjgNacVg0wcmI/LcEoiayX4sP6ECGOB8M4obduOj+FOWIu+mTptcAri4
z6lF7RBYck9TJEA5xtkb1eHzKazTciYPc4BDX78hXnVi0w6bGMC419Q0k+y+wNqSw1bUBvP7La62
cJCTWu5ilx4mL0rWjvut7UfcAMkiwboM+RRhaKvezLKiyjD0tn8Ob5v3jOlxQb3+FbqS5EjRon+u
locUcgWpFhFa1T6rja2S4RETBt16bljYPaZaVHMa4zPjmwSqqV/V/eNT1D03fB+AM8AZdJyZLTqR
Gxo6TIM8KOZc98n6ZkP+MbKoQFtL807AUeQYVYjQO4j/wnNCWCr0N+lrN79rUQdxGVbgXSHJgquM
v62PzSnqs0+XLfZEdzWDj3KwS9FXDCpEZwB0Qf2xE+vnStGWW/Dt1LuDv30YdSOdRzE1YgD2XBeo
As5BhcgOY6yetnD/SXJW607e7CLbLd6LIkdGnVQZL9XauDi012uQhI51x7dVDbJTDQ+dHh9cASSk
zK5pmWqS7qmgRKZQCKeFJOGn+fjf4kFQnF3flN0iUkHqx2l62FDEC8MAJTelPUC4ZGQL/MlhHHoL
YmWapNDDqlVavnGzjkhblSNfiNd2AciHFLvbZmoHk0tQpaf4MgBiXhvI4qbWQdp/2jbKEIiPNaYi
SC+/aD5AZSO8dU+ZpvDjiwT7pUJm3Nw0KrS/ZHLngqifT+7CphP/ODkvIXNYoZ/PLgFuaUhLwSPb
AghHbBYYeg44wvq22NAtDZQp++jhQwGnTKIu22lY2bYa/RkQ9RfSm8E8lrOhszoF59Ce24e8UYUf
icTOkNtadrq9Pjjh9g8B17kBdR9C8qevdmAxJW7MSEUFVey2PPNUXQqKE83x0zYdzxM5X/kHrTSs
uz/mCCf9SAtMyaSOUB/fwOhjyGi9zVUOTxASu+KroabcuTgpwrKrbavh2icOaWVPJHSk26HTyYpP
wN63tZqlBBmOTiUtjm9b1hWZJUSxWEJXszArf75K9UCPEOKD/GasaTJyrJTZ/ZXlJ+BHsD6iqMfH
IYkgO61g3msKtyjXEamUYw1moIVAC4q2WHO88sYUorsz8xg2pz7C4zct4GxfhUnT3GIdWA7RU/3H
Scih6EVqih6sYYLoAl8gZlem1ezSUNWRV56+d9KRVfNv31Ih9YFQPk8ajwihGii8NSjgKKfrbuZV
TrirY48cusCUCpLCVYK8Qq28zFHna5l4QNr3IHUAsOv0dAb6WdcyIXi8wqDBE7yumjBcFramF+ke
r4Fq/aGJk/94qs9koSSwIoeflVXSFAKtd5x21gyk1Gco9+xlyAAuJVS5blGL99Paz+ICignzu+I4
ebvgVB22T37kVX1nq05qVq6AjkY9F5hv/B2KDabTZb9S+bfd1wxBolvaPulZ+jCu2CKzNcDb/Ry4
IOukpHPVaFvBG2FUkKX5f2HUCDQzqbUNCmBY2X8tF/z0DaKNdzufUwqrDtDWXfDeHIX43axWLtH5
roepsrplfkFVuVpgDqBzrDEQHYcqN/PcnAkPxWFeLQSyTe7zPXjMobTg6CnjVgMwNhojeASpQoIl
UIS0GJKggOfG7LQOXhnQ02v5p6+vu3affzejgtBxkwP4MA0yabaVOTfuIWNwHbFLOiFwHEt30Yk3
6TfKXL/g27jDgppwwgWFIu5lPcr23A+05bKnhktIBrvbJnF3RPw+rg/ISbXi7SoC5hXNP99jCeoE
+8vwmKBDkd+zaAK6TUQo1pbqFcVrVR+Xop5PQ3SDNvV3JLqafWUY3jvjo4ip1keIcJ8VHoeV683M
zeVOtCqtUn/niRgrtaBnNYbFIcnBjxpAf/J1VjtuvKd35vcP9JRShfnTVCJ41LCyCZoxgGDToODm
ayL8xAZXCu5clNYJDSCHh65BOeSyCkW+1j32kooQrSLsF1xYgSprgSc+rnhqunh6AknunBzDWz5v
RnnsmInJcOS4UtOgJ8aLVPpyVsaw3pMrjGEadpZ5CLjlfE4xc5nuPwPd7gMjB/dyGUGwm6s8An6N
T2sfC6bKCAMLuvNwWWhwVzZtg6fj+mqE6p+vpmGD4CSoUUqtY23QTSTvVA+i5h5vhMEuSIkIzIZ7
CDsZgfQtsIlmdpoHZ85N7euFVBRtKnRS1R+X70ozQORs9PcZ3G+1Hbtir8boaGXaOB2oo60iQ/vn
sSWIy4W/LZRpBj4AjaBk5hREX7HbtDpff2WML8flNa7tlgZZkNbt+ttEOSOtt0BvVVP3i+o9ekhc
uF4JEPK9fVyjCgZ73y5TbhAuO/jgWNgbWo6vDd6D3ODo2OvW/CfvSfVP+fBE0UMqNWYTrcJHl8cU
fkWPn16mcqADYXxPm7VT5qgkEvIQQfNRiewA0tcgPhp1Ui/n9/u86UFgopqYF4eRkzSJGtvsLfT3
layXV2JjWZrGI+AW6s+UsDjHi4nkrKqpTBZ2egtPimNqxWr6lsetWvmOlb8F2/s6jIs/k2WOW6la
pqmhnifts4rRPNvDFPa9FDlTffjcUV1RLDCM67W4eW6J2uf85l+E0WPB0A0XtZ2qU19pt8AFkYX8
Pk1ZRWuQcIWVRD4grrG7UqowKEkM2BcU04z35LehNUcLY5DWwe9eO9//XGOVvrzNtN0vio3VuV8n
bjy5hbgh9gM/wkBuC7Wwg4vLpt0pR8EZFDEnmp5azNG5UVJDiVpVwx2o8AyGV+ymsoWejjzoqZKA
T2yMLAAbbRYzrR5nqJveRLpN+bkKRgvXNMGWwy6lKHpT1zz6AExzjKVfhQVFDS0ZW0xdDk5i+eb9
tSfAhmVyoDDqbj8gWBFk/4fZ/RpcjnFw89XP3Pxc1qbEwFVdopYuRMs8Iuz4TLK54YDkvofZdE46
YtZMUyxBw6f8ZZlXnu6qYbixiAuPdFpbvYBK3zNXVcr+kWtCUkMnwYyuzJIe7Psvtnn9m4ojhsEW
YE3okaW1NPVkzwXQG0XyFeT075cZGzDLDLRuPBXH3Ld2YRypYbDWsaJadspnIx9bL3R7GiaGQVkD
z82QRvV/DcdLNIRPci/u6vaDWL9vtHU/mS5jEUHkxL0TiYr5C0bedJrgv/6M93GZjn9+rA1rVywj
5L6B/L1uWGBRc9w+J7ZIwIin+AlmS0uOFrpm7CeTHu10AcwRUM+yx8W0UWZ2NprQhrI/Yo+F8x7x
8q3xGqCa9KtVzbiXjjGDyvuT5MnS/eaULhiKTpJZGRVwgnrrB9lPTUggdK1HQnorwjUnwPFsLl3f
qm7CmoY/FXSQVUJpfyXIHvvC1b/a6wEzdyVj6ZKrmy9nTZgsiVJw992Q/o45/assNuVSSZDO/PaP
flIlHe++WxBBvHO/cNE7arFosH+F/rRb5TSAHYVRe+WaxGW6KdMJbp9f4dgVtw0y6XfrGNWfDg2A
gw11jxqPYJ+YI5rd8Yv730oMDqW36CQR0O4TzmgZxKiwXA0BWtxD8pfvmXIHnV0AsJCdcoMBoRGr
sTgXzIQIQH95Nv23owcpl7ry4Dd0E/q7WqXPJOdHi35YyxkaRu9OwH5eYqzAYOD3KbbZ5UUkhdfn
cTXinB5hbYW7DjXH95dveFXIH1K62fPLGBi4i5PjYyInwN9kAPNVwP2TQrSbuXPhvNlpFfkjjMpM
OTP/CXFR9kjcWjvN3nE+pUwW/3V5ss9UMH8KrE/pFQfHp/NTExpWVFAwEdoMng0uEOnxRVyClYwX
/ap5GKCGLyUSqR0Q8kUmLTjF939DiLPq2WJ9LZaQA91dyfdmSLV8TEvo1zI5ZdDvzbDhetQzMi72
BT30rufuSeFme0ApS9lgodNpqLJIUKPw1MhJoVGybCTyU2libjVVdE/0GCQe0UZ5Paw0hiIyw9eE
FZ9ldeaiZr6L4kMZZo4IFSfc1Bf4+Tra/jVPQpwzCTgWvduseP86CTJnZwa2O21LV8r6UQjplxIe
UTlQ1YGzbv6AZIie2C1kIevR3HQbYVuwUKIb5cH5LlULX47b+SH8KPsvmVn9WFHCH+DWYTHNRJXR
GiTlyRVxwm0TeF1yWqUATzOll6XZIWPYVYGXMRQLt8SJwQ8/kZXKjL2PENAf7jN29MWh7ycr3lbA
GN4KeLNvpHeqX5nLDBq7912WP/KtnHHW568I6vX1NopR9lIPI7sfoeN7WN67edv8EVY8dwktvM3T
y/IDrd4ZElF5THULtTRO1qwoL6R50MSA62xb2A7yMLdWrJXO2J07ABme5tP2vTifslFRFw+os7fU
ZbwCr+DQ+iWYXX0BdQJ9ldMnywIKEJZ//jVzwClrXHEqhKcP1F21Rj8d0l+/gA3oIyQm7i/68ya3
lOv0QxINVYa4yzdo1xI9nyxhmQqHRtOd7t3FD+V4nSX3RhlGsYTvcZ05yPpdcHdrUT2p0BtIWwy6
LarpiybM/gvA1hOY5292yt3dnIA1N6x58NnGMHZ9VEBAIiWz1EX5akPEi7O2nJDVnSf3RwT5oNDl
SMsiO4ub5UjVME2/ownb3nrvVqgrJdlYw+/ziusSgrYp+bJuMO5l42v+LL2GdXCb1nbwTdC+h5q8
XPm/Z287pTg7ej7dmkZstcm3Wz85WhfkAI1O6L7f4uWrFX0+zW9Q1aKUqlhUCAGDtr4lV0W76pTg
YEm5XvFIAfWvw19cwJK69SS1zpqOLzgDjK0Z69aHAt6+08UZrdEQ/xYidXkS0DvfNgZWpoPpyOQ7
auumG5X6tw81q35KYOlJMKml/6UHO129SQj69r0uzxc8Vd5LRsE5V3MaHIOBNLnF7ZRycHcAKcWC
qCV39FM2BdvuMu3ybap+NcO+Qxk6b6xxhaE9ZmMWa6VHfvUeiR2atNtBLvATgvXQvtVTEdhY2llY
p4f+r8lB/dWeWwBV+36iVoC5Pk7KhcOZmeRy2sFY7f9lvfQPcojllYbIV0sf/8qHeGchkzbEIPJ9
GeZIl6mToZ2Nk35kIqiQwjt2mRDA+MTPUOs/R2pTW1rstIithyzrVf2P67Ga5jB6puzj+z4xBUtp
d5Ye8CUNpKwpqFNGGNA9tOm51Hf806R9snJbmskiD+NTXKdnX/cNlG+7T42qYupGdD1CSl0gyQ3N
oYURXYtVWpz7QdZEJaADRCG0gbVuhWi51YEpP8MjJLqzg0vLZSLCVE+2vafsIRaukW1fAs1iZOtF
/DTksNRin+N2RV7XulPDZddNvj86Gx4H9+w7oIYgnDe9RZC+MpwDNwHJpBcCIVE4dFkqey71PG/k
5VDyyHEwShFNBL09fcf+eYd6xmj2Tymng7IR/yozp/Qzwe4bIn61VsgHCXVlEn8OG7YeStcT5JcT
pGTnL/J9FaMUORKbrJM423M9X4314K+qDX1uun22qv1U8jrWnE0s8Jpevkufciqm2X7jdemDFFaH
kcp2BUAM4Wb0cJEys7ZgeJWliPUjZimO19j5U1Ed1W4flN4JrXCydPIbpJzVumhWaCbWSg/08a/H
qDl8+LpX1aMHxyeun8wa3uHE92OjGR0wy9p6rG/QbzO7lQjMLacwVctX+1RZOnbCIjo21YSdpA9G
9w1UQw+D7HYRLL48dPUzhuMhzzbSOH6m89UeyaGrvIK9gVUKVzNVn7Mb6lvu5H2E7KOcPFMm7hMh
zZnmwhYTJQKCr4m3MfNJ8rfWmbpyLL8aa4+reQ0NHqHFjrl0Rp4SXHzVQuvBzEbTlUHGTBfF8Ort
FfrBZ/2HX7B7PUStLBXnjRbrjtMYANwVV4aMAtBMo96HTm4IW2B8Aeg7C8tAc6T7mGjpqIBa7Zll
aAdVtbV4drhL+RdpsDNcIMCgXvxCVEH2Z/r4YBfEiN8zbsIX1l6CavSzIMsFbZl2cdVaGiR/Tf95
b6HsFMQsb+7HLYNwyVxx7a9XXW8orTKYrEGUqBo2ngJcSu8hf8uQ9C+IdxLxpQDKt+64tiBoI5zH
Ag3mG+5uBvx8bl62Nu48lY/F88IZQvrOHfAgTLEsdxQn72WxYDRl6kpNsPFJj1RBkQM54AmNcaZB
UYqTAbM1MGWoYIACHLE9acArGvRPMuisS+v6syWKQWcHKvSOFQFCTYo3Zh5wd4SKlZSOkRL1t+LH
7E3EHHiJHezJFFaGsOF0+Zlci99TPyReULtmNcNBYCaA8X8DwoQZlLJwKBMPdixw5K8XlyU+zHOh
jgmYqdH1JWObEJBWm+DF1MgegN5Ck+RTMYaI3Fv6L1R0QMqciBRu4xe1R6sLt65IdJQ4M78c+Vh0
p8rC6cij1/bZDexd+u1bw/30WV6BSpgGRCRjKx9w0C/f8K1eUkWm16wgOoI4iKpqHkQyRWKSvd6v
5lnNiE1B8PGMQ2OIh8A8rag9kX3DGUpZ08iRbiBFNiZ1KFa+zORvblatMWt9JPlOFF9EPcDF7ErV
7lqOY3Vc8VOGDaXmrtYokkIJoguc69d1fTbB/WMfF/Ah/oE+DRhNKszeeegt9S4Hx4glLSyFq4ld
dygD3srIK6+x7dQjre6a7iKZioDnI62fNeyldHWD8E+AVk3Oq0sgAizBL7sv7K28+DeQG0PE6RfV
WS/nUKC6BmoI7CUBSRaW7GJMpXwXAnUtwfsz7PhcCJTa6Ck/mtE3KBHSVr27EWoYDy7AWWa3A4bi
ejPUZAnhJwqByiwdug9Zc+N9xPBgx7oQKRgb/5e4UZMv/8nXE8EHTfPnMWfrRlFoN5sGi5kpy/rT
W0pZJyorfnM8iMpHpB2AHBxUbB4cC7f1tCAWvYXA4E8/CQr+LlZvm1M0YRfO3zTl81V+OkkSkhyk
x4usikPyUDwwLYAr5RXNA5yKaZXCvfo68s5n4OOOfllBj2vCvQuG6dPi+kiC1JCheJM8aMNedN3v
jH9lYkb5SgrnAcZ8OhaSFHQ/exLvVxKdMXot+IJ3hIFROjVkZDRSJTrVxCphAGW5pK56HWAB2N90
rGZZNSQ7Se1OR5PCffagWZ19L5Kw5FwOzfVSPZ34QebIeZE3Nk0c2yWphEMkrO3H/QXID5xCOKY8
KZfO7/wQkwhbHH0p576UCCw8jS/nzoTq/b1CPTBpmvKnzaOyrf8q2NfoIpz/4AWofI+9Mp2X1rJ7
OAJGOGCq3jr/Ekdq3/4D89A89CCie9qHSnWH+/qwVgNawTicBRUhdYFYXO5UUQ0Mo4iyXNpLDwx8
5gFMYi+XIAk56w2S4QTAHZmxtnfgbySjQSq0KSVjSNMi96mBcMFs5RNt3L6YCZZ1qdqb6qN5jNLf
uOX/yCoSJfVF6StTs9BFbWuGa0fn5KMW4Y7sCTZrnv0CeNIdeEizru9abc1wszZ2KJ8bED41Yqd9
G+ewrITdVq/5ayS/frkT3IdUvgLxioTvhPwP8jCv2wRREiRKstp9lQfTBf+VLSVsfCs/IdEXG29r
NeoT9z2xa3PeNPlOQ9yJug5dENMOV5cgxsACyaW41nF1ZAil6aWWUJsxb68zIYV36Qrdy0zFLyGM
6I1js3wBS+YdOTuHbfDIECUEAdW6rzuCNRM1FX8XO3cEOOpg0Imah5xbwKIs6Z2a9W29mLzFPq4b
jlXhe4ovqKACc7ev+um1RDClfpBgQrDNrHl+LBZNBXDK+tT/1Q6wCzz3BC6K31BaTJk+BKRL+GC/
d/+GZ9SlxbBYzWsv+P/AlNrb3FNzfvIuC7an83UqgTnlyZsUm06+6vIDplKxeGiZezU7/STnGT2s
6r9UxGhDOsjIkFzs85JvKB81YjiwJhIQGyxY3q9naQ61+MActUHxPjxE1dFZsqaGUaGQdJp5bGg/
joEQ8RcLwcd+dfjfU1hHyRhwbHKlLDXGXli9GvX8ldIHi8oC2Al1edkEa8oWLrRxSeJdc/qnmXFR
h18d3JleOwP455zsKvgElTkHZKCJ9ap5DlBTimQwjAtSFl8siTQKCt0ZhU6gl0wIvrhsm8qu2PwS
dCDhqWbp+SUgWfAFbFeJ+rUAsKB1nPmn2p1UHaDIZkkKTHHqazOkfdC+MPtfTTMNn/QMwSDuRI4t
6il4eifaTUOBxTIIas8HCU+ULLsR7gaRJqNUPYKdqiBRcIBLfywQREWscJShp12MAENG6tXaXk+h
/RoZWmPV2kFgTdzrGVnXZkt2fVMxTj4/NL/Io/kZNCJwt6OkoqrX2h+iFCPMebap3CjdUEV9KtuZ
WD+jwoTUnuiYtnz+lCFuCowNoomNh+yqAjGKpl8g1iBewLiBmnaeOOFDRnnI7Y2UMYk+rIOKijNz
W3yl8QFzzx6BHb3MtRkBkq4fFlLHhv93osDrNAdE7xmnOakryDPXbVJcV3ZEhuC9g7WDU13MHWgS
qB6+JxtY5fChkg1SyGHAs248wuzyxkVLVBAhpv64ydVawvY/iCeqX8bG43sOyvAbOI/M4wzvhXLF
0wrPZIBC6bHKXxLso+kmbGSpQ6u3kIuJBkeQ6y0YdguQVbEkbKa/OZOto3anvC+8KoxRxZNj16hp
/jrwNJuJuxXu2JytdEHsV52vpRLCixZgd6JWYfwOOCZBzeDK55H3E00pGp0lxC0nMSdzQcMB3VtU
x8LOD3vNHFnKWv3R3tYQO9GV5hMofaAXFPjaKsXgSCQFUbgvwOaWfAA3jzl9gi5ZW7U4mFTzfjpb
Yp28zbxxusKqSjnq2bmBa4Jb0NH/tO8/a2vH6MzqXWVihtWtWowJE4poC0s+xPE3X+m+qh9AhTuh
hr2ypJSuogUPDpuxoKWoE2h0g8EIQJus7pbxoXgsyni+QcKb1kBgG1FnKPz1XiB08jrlOZ6ktB/i
l97Uzuzpt+/IUS/Q+Z7eE9BY/2muuBEi+v3aKDYVvFU2/MDAmsh3xWVqGcyeHp+uhg75KM7g8+fU
jyea+jUq2pmuh/bdrX+TqW1CceTbxu95yMJgI9IQr+Ez9UVSiTAhDx9Hnib0uFBb91OMGZjTW1tR
H8Ij/9V67BOaY94fMxx32NvDyQ14YMFMWggHr956adpWCLqH2BHPn4dq8SXwoWeJAduK4RiLL3lK
UKyDv8pwgFhs0bSP/sQpEdy3sAv9+2i5/mT3F8vngBrdF+Sa5Ps0mHdz7IO7jeYreTo6s90gOoyn
+6vxX7zDHsp1a88ULBGdKOY+DeoDFFUDnC/Xlb/DsS2C9biaYOLy/Jp25ugyoshUVDnqAHCVYy0N
XBlJ+S5BISa0/acGGRfv+dgaVQoWUxNuwSN8K4LlekK1LSttqMNf25pLBd5bFIfhVqueSLO3+TMn
+6y9xDybs0vzSA+M5aEczlnkZ6eHqYzKGPhFKyRdDUvwYZcylSRiW+X7tMZUXiFebUn0NqnvluJq
xPZE02JOCvY8rqQBQ+A7iOLRuKeNuw+tngEs4ZK9AgeUAMQ5RqmtfyT8YD0SIypAidBeKuW4HcJc
0pvZkHwqxGHfiCx7+LaY4x/21YySM6JPXznF4xPkpyNaH6aa55k6khVs6vmGbiaQQtn0rGxhbcNy
uBC2JSpvmcZWQCu+fqGR5oBQHF53CbEOTx7IViBk7Rv7zsc3cCh80Y7BQx6ea0wJ89iYgL2Xu99z
ry1GDFr4DHkm6qof9wmFSopDYV5o6Un25dDM+l8bbM0u9q9Cl5VsTnEl81YaXNV6+srRh+SFB9Sj
xbaZesxuUamX+Xw2/Z2VUAoxrP00PlRX4OP/bNqBQuA7ANzMuO+K0gzG7JQcqtYFtUESAIH28sMZ
940M8O1DOZ0NaIANC6uypG9eQyIRYYvQAGaW73ociCQPxrFdgOi9imCj7+V2dUnT0WYDGclWlguz
Xxo0//cdY2TVNfxDntoWjzX6cP1mmuwOfhiAfhYdWHYoaxGkK7LxOKqH34DVA7lrEo5kLolYfDg3
l4inlzzt9mZLODgx3cNsOI2k1S+gertGG98WcQdVWR4rapCPmcEW6mdZl+N5R5mgzCuN0PIPR3W/
EOS4E6EQ4pPA6D4kCja9yARIkeenPlpOhbBY2yZF69br3RCd31a+alx/jrMtdmLqO1ETo0idnJzx
5WHq4jJ5OfA+DOEtAQUOF8kaJvecnehdtK0Pkg1BwNkApPnV3caf4M+0SH/PqcKccE74/XjMkQN8
bdKsYoc3IP2CY4qMkdlyFEIjf7fhU7e/mF7L4WACI7JUAt8d9C+afUGl03JG5Dh/+Cn0CaONsNX9
s2DU7mGo3lbpY68hot3b1L+gSS1NyiJO91RIolH7YDkgqIdE32Z++vlkAxS3ye8548gUgNOANdOT
UTu1YYNPnl6jmsiQPWe4hW2M7MgaIl7LX60bfD/E1AGsMlRSnGVAEqEETeG4h71d/gLbatOGcsO6
klZezAqvFlihGWWm3b/8sfYNLx0eoHKe09UPycpzo+TAsx0cNGskN/Hgub4pJohsmtmCvzfgm9zc
uS1Lo7ybLP8AW7CeGGuI63W7gHIvGXN4DaX+qEY1W4xJaB36oU2IM8720vcbAmG/h5piDv18WmFW
lR9OnI/lZrFAb5ShZYGBtr/P/C7ElpEeUXerOlpp9xAaOCN7BrYMdjbeJ8vrQmoNH0MBKusrLJ3d
Sy+DpqbGZOWGkRpuPauzWA/DVrJjehh6WCQPjZ/LkmW5wsnCXfvlaCCY6Tn+AWmLD941hukSTmcN
UIAjfVWXuY97C8uTpRrYU6C1tZILZcl1oNbr0HYpsUaxEpW/bk/0sfcGZgpkt2gCQX1XZozyrr1T
gFjSr+vo4e8BV40TIEcMZZIJT46DdL+uYV+fsIsw7R+DrYfHmdVrLEGABHlgyiKAYEef3lY1KvXj
t8UXKEc2QaTnxRmZIjTyxIWCawLevmsh/bOrMwIsVa73t6S6IwZrpiAy6oMdVSJNwC+adSY1OmHO
WV5PHI4gY4cQZowfCbmE06633oDzWdGz1wjcB6suYgx26CMIXSyEVj5w22ERkCngcFgpNX1uxhpm
Yk8nG3wtYZ9koxo9k2GjN8NyPEMKNR0jZblsu7cMACiU/TBFbU/zDjLoOZuYch3kLFxeb3v5wGf/
OKdGsb7ns1FGOOdo7WBfbvJfnAGV4o7bOSTotnKF5erMgsT+/mfOP60cwASwfirJNABYjdmBVkkm
OHI9TmHXpvHvr+jD+GR/paWkty5OYcpK0qTx4DVNB4E8bvubt/PCjSRGqPKJg3a2l4S+3x6LdlD6
xcJ9Ur243bxX+lIUFElrQGtsvY+/QQUxQIGZXZ2eH7lrl85XprONE8CgwOF8gK3F+z7OqOJ3s8Xc
SpHdhfvJF80q9X/eB0tEoWUbBs3n6hgz5q+9ZK9mZxOrTUMwLSMJy7XWLeX334+74K5wjELoruC5
dF3RGGqdnYUNdO7JAP+sWPPQkUrELkCpphgaR8MSZ8cwzNK4HSyeKW9L0HNtZq6Ei++ZH549ZvdP
R34rgFE6U9Di0y0DV0daYyeBJ1N6e33ZVsiOiGWxbtbFZ836FKZfVth0hiF7o64+h11iltooYXtT
UkmqF80tABkeWAwobLCpe/50kepMFCkfLHlOXaRcOrNElIZ9E55VUKE+VSCU41S7Ic4gwpLbylab
JV4KQ1gsTgfC5PZ4xvMN5ycxbpVucQe62iqeE1lXou9W5u0tV/27l1dy+DpMEWBjPp3n6alPMF6U
ZqbvUh+MiRyJHegRjSHVgMd5hciADRf+XGET9T+zaffINXEKmKuTVQ7Yrjjaz4lpaA5vVaIIhNjT
xn/NFeLclvBIZf57yHz0LYiaGU4qqEoiwW/kCrFkER+4PQ9vZmZ3QsYFMLsxYT8pYoTi2x6VS6HZ
QPgAub9bNhsvySa+C6T6IYYhnRvrzOvDpUHHWCWxTPnp4WbiQcCZaXog9mG625iG3WInTMtWCZer
OOqa3MWsXPQo5eMjOROKGTvqXs2rFIi4ey8rUTkS0gs+LnLgVjRHfoXhgdoI5/I/DNugBjJWTVar
6si/fzaAuBjYecISH6z3yXz2nm1N/A4ON8Jf240nNO7XCFo0Ze2pxaBbBUzRrYVGjDCJJDfkHLRt
GAXnLh5V4L9HhNlMR4ii+j8ZXUyH+NuYOJmozHTWj7bG8v8sZQrdFMKm387usw3X7zoveBpaxscd
dfDFOikmrgx7iy4WWWZ6Ox4H5XW/vSPJwuV8l5EKKPqbGcmBNQrJ2H7O7PGzxM2BiIMSOYTHAs0u
ZPOsGLV1HPIET4nGdLL7NpQRnOEk4zAalulvAJq24H12leCctT/ed4imRtLU8pjP/NjfLzCSZuu7
1e+v11eDpuZt3996dOKhnFHYYgQemJ3baYUmdog+Y074uDLEgu8JBH8NtEBxOETqQZy4wcrV+djD
q3qFpgq3XVmupC6iknCBzyhaYJEB2/2sRDONGdR310732tr1KRbaz8YFDN+iyjY+9Ae4b09H82ao
voK7nbOmXNp3xjBnY7Eh8gdUIyTwOT1uEp7fXzFNsexXbDzb4Q0NvTvkEFvu1/GlIrRguFzCdTik
EIBBwTgKX57MKoV6ABlc+qEOSBx2mWJzvuctipJEsP+8y9CRQTt5WWQhMh/DBuexs058F0KtyQP2
zigWWmA90/eNh/jkxWrpujZJ+IgLzQwOdn4sAA8TO3JR3KClq8HqAs+UfREmkjJDN+MJo6YlI7Ed
QfQ8AqxdihKj/JTKKEB4g4I1SBDs7sjTs6oRQMlf5Xf9y/Jj+Pb9RirOlb3LcQiM57G13PfN9L+d
0wiJw6D9nHeitNN3X8rIiFe/7y+bzq0uEelIDWQfKzleeC4SlOKBBE5JDsupNiTaiHA0e3tRkfvA
kR6ZLLqu6u20ZXMiAWT9IoiYb7CR0UsBOoPWjpk4Xjy1vEyJcqMrvdIkGLO16IMnHypRQZwY6NUk
xNhvpIYnAFuBWf6StSUmBw0T23dQWvjfAKI6G8jsnDFH7nuFIqLlFhdxrwL0rUSO8pvTvsA8VUw2
W3pMPC3UJRtXW6gqrlNqDalhTiHiyvYNB0ZOemzfiJIYsNzvLq5WNjrqXBRrgpXGifS2JQeXurZd
GLpmNcjTYpnYAVKmusvcCqW1Kc+JRDeXhXvsEs0/6iUnQJq53getTntl0OvZ1O3Dmz030mkKLHOI
UdJoG3uHeh7HMCAEi7WKkNdjrY4yWYlf3WYaKhjWCjkIn6koavUHmIsKBpRQ1YzJMgGSFJsuCM4x
EkKEcBnkwpakmjn7FM5uOLuUUKw/GF6joln8UKfARuE5GfKiTIzQ0pepKQyWRrmHsmGfImzOFbzP
nq34lQ3Ku+zv5g5/+iKfxzJei7iWK0GG8TUr8Ml9YfKYfZhY2FxuHzX51RjRvcLcVPU7qYaKXvGa
zZmMvb119Q5gaBoOAwIK33BrY32YiXYhty8+h1q30Aiex2zQfiC6Xw7WAUYJbZEBdMxjsJMHF7Uk
dltqOaDgEZzuYSjV7nlCjafTzMl2Q2Yuin6XAhKQqcu80agqcZ4AuJtnI5V7GfU0MxVMGCE8Q3SX
nj3Ok+3MYzEGH0WlTLAv5YMtF801nbiOa/KDk9E77MUnCStT0Jxm4a1gRzVAh0j56EkE5+RgI2ug
smyPIGm5Xz8ohgrN5pAZ1CpcwEdl2TSG81dGxBoVu5EE/gHjuGQDLSplFDjn31qevU6bgYqP5nAD
y662vPA/ZrNoeBTJV9vv5bNJRUIy9dhUEtJkMt3EQMuQSfoUKIO5aOGHg2R/L8enctV8j/uA6lFm
RxxNYQoM+FyoIeun9mtUFIDtbBQwEeZVf7b7VGODHMptdo9LCrownz75ggXdvcS7YGTO+P/t02ld
5aA6m2Ej8ZP3m5RjnP8uRHP2Ki/qZFo1BXWq8bSghBSypPFXYM/jykJOlYvQn06AUNDKvE6SwsA3
hMnL8qDcybALxSZAGz+F6LNvX2wBOUDp2OqfsljTeWe2dTX86n4aESaNN6dIa7fwW+LFHkY1cyn8
fnI7UQdxiYnM8kOy1T1shOYowVBIsnHH6VmFVhaoY60sTdw/jeXfPDWdC2i9/AEB8Ua9EtTTK8U9
klS7/Z0GGTClc3MeKKlcLFPJ2UP5+70MAJ4PKKk3TgT53XMdhX9bP4RdOAH3Ndrv5xzV3+X9uSlV
lIE+arW6XvfS4SD/nay1mYYInd5YH53K0aEZUIcs2ASjWIusB5c5+FwIco8D5ABTVLv6gCTrg1BL
abAMCrJnVBy6I0gWEOh2tVdvSykOahXI016AzS+ysXsNV/REXuJsRXwjuCoqym5Kmwx69xPgLwDL
8HEWUevMEERJcxiRMkIOMMMcTsX8s1pXaIO+lCqmppV9OQBlPyejm795eJOZGY8PBjcboQbYL570
tjmCffkEGmQ8+dTMgHCAfh8lq/xkCa70M9b8rOne3cMTo7djl/u9lfrx0AFoPNmJzkLfNvel5I1m
gHkFa/KvAb7Hvf85vNJ4MD3DHVvFkMJHl52AB0xvUdBF7fr7NhHwvmZABd+GOk5ximlZr088X9UL
35okLQqRTGTTzHnAIDWfej3KLYgO9uJvgOack44fFU9lkx6s6FkGXJdXX9kdQMQijD2D9cTj5yj4
lLs5xSlfwTex0oPNl3eJTzBEF2xpT6nqL2MswZzmK0Qy5WzzCfb0e+jpXhelmHWviVlfv/49XdGX
Ln9h8JXmYOZSwBg9CMJawiP4EmgnDNy/TeUvXYJdOBmBo0xk5khVR1LqD9rG7UfM5X+Y33sGbsCL
UhYVsF5yRqxY04+Zip4EfNLG17vKgGXRZVxMhh6ot4BfPqWMcJq2YspUL2h7h16UoB0UpAgTD+yS
1pYPOHXAnoIvRTgrZETglKkojTFRMO0abDvHnArxCV2nIFR1UrbBqeErhv+i9O8u2sMHZSFJ9RYk
kGn5KnkeYqQjQ7lXzp6y8frR5jzZJn9LVjwAcX8Z1P6uZFO6KvTpGo8VjAEKNEnY4oGN5ZzMMYYo
Q30czFScNK5XYoB367NdoNZkjbJmJtdNXRuchTr/aKldkizvScCn0SJpi7j0lnKbJXtTI/gTU3hR
yX7flkKYhxmo/EU9IXN1Q1vLVVaGyyNGvEKQMSU9hKTmUtkAty6e8d11iaLl2FGO4bDnv8pHLL7H
8GBqi0b8mk5fa54xuUZSC/FCXQcH6EtaTSrJZ06lRF4kXkmGdIPB+mvWMh8s5K6ZxSnm1bzxKDQn
98P430of+aswli6jZNh/solhkv/CZWWpI7Khkcrj2ePjn8XE3SoZZF9msnQlwz4riEG2/zw2qEUw
DNB87kZ+D2FM1bPis2W8d9l3r8sxDTnkiojhpq/6kAN2i7iQ+Pp9fFhXbIiJYFoNEYYC4tVNLhgT
3CHUwrjCtzymsC6byj2G3YAKpgnTHZKKiGFKZ4q2ajzfPZVNvgyQLs/nkGwRxT8S4aM9ftSTyEko
GBFgo19ujT9Mb1HCW5Puml8N0DiFqnlFxvsUCGWLVJ0Z37MFRl0GCe0myf026wWzYIr315oF0Mr+
+OrZFV9YamRIN2RQGG8xNU22Od+llM/Ibhf/BApyW+7Yc5/fCGiTst6NK5u9hlLJL1XRCSD8sd6i
6VlWlDezVcQXRP7zQlsFYckCAQgFXLyVUpZGCRp3XmZMSJOqYsZlj5XAtCHB6XL/OOD4JcTovnBz
ILMeMOLD2xkWmt030llWOhUPHVTjVx0lCBAOjpJkmAa+fIhtkp0unxzwHzRepGA0n2NKNJxCr3ap
YasekRxqwHJVQ8KsO+6uqth1MgriGYfOtqfSEFEtF6PXVT06y4Ip5JTnEHCIJIDcghE13B8lcius
hNblc2fuGebjua1H3ImDWIbOP6mmm4X/1utlcNfy0bYT9jBuQiMVumGA/BaKLqTFik2swJy7HTbx
hXspHFmjn2UBmBkQZYUGZJmRzEAjdKXdd+gUVCPx2gc0ig/E1JZPzre9N0Mal3kMpXAw7imv/xbn
c6vO/PSACWPO+Gx5c3vMQnEK5TkIg4zTtAdmUM/CLU2/Jq/QIbow6pw9r2m5DGU4qT4TVNtp7qso
Xl95MIedbOrblIzRc5SIp6FC7JMEpFdecuT+rksoeVHH/ds8EyNLPuvcNg2KuYlN6WGkE3ZV94wy
7kg0/erwF0Sc9VZwTDUHDmZnqMoH7o62pz3psK2KoA1936/DIPovu1bjVUbqaIR6vYqCpmFM7/V9
h2uoSepfZpdSWddPqGLXN5REsViOEm/HCKNpoxyUv/AzD8JN80U21UPEcaO9CaDPJuwPI1CaSmLp
+q30BNjzTfJbvJoVvSf0a5iqCy6Adr1NGMn6SmECBEJpZgZce/Y25WcqAkc7N8P5boKvsPE+t0cP
R96kMIuM990ZBC4pDKWYP6jFE7Ti2sW5HZFdXdEjm9GKhJLeXMzBMZpxt7L5trmahBfLy25NU26G
e/U4uyvMGRIMtqsbpBkh4ovIOPZvhKRR0v2uFuyjb8hC4tFV/qbCBnnSpWFHwL0Pg2p0sGjSVWcl
7cgTrNjE1Y7o8B/7deWZpWpF/MkgJv6x+SccC72vZjkp73H4pDU/wVXUJ1sKZAUl6uQr7F+M7BRu
RSL0Y2pHwlwnFrrAYvoZVoePJr3UPjjTRvlTwqVuTfiWKScWN7hNmxO3mV9k/4f6U3MpFTMaSZHj
SWKOnxeOok71byzMZkaVleno9ek5RntTcvRFx5GhDsKqM1ekoRCtgE2Sq1YSWOm+CPcO/mpor9Xx
wQ0PGXdK7ycoq8XfYECBCk6gZIr0EiriIHgUPnqTqklkG/v9vdHCTOC3XtQvOfQ7UGB0y0JuDsh5
c3rTJQtAOaC57XGuxpcO4vi54KBedWBbxw1gPp3JLmwIvX4bwN2Vg59unSndeZBO7sJC97BonklL
T/VH3u1YJKAn6T6m7V16Kwem6Y/FXMg5Caee1JOhjm/b8fLD0DJBuFa89dwrvdGkK56WKTfayq54
imkEMYzrD4pKJI38V9nYXkFCxXxbZgof1kb5rOfqOnmlapdBKDqSLTF2Td4mrfNpZDR7RM80x9Ws
Z0aX3Q8Q1CShBGdklfVXUy7yEtuBWNkAFANDWpFvK6EL86f6aGyz4L888If9tcMlogk7QarH1vm5
HFNVfmBjXpDFADSvwErMQK2aJlclUtw9yQGmMGq7266bT8gEC9FLXe1vOgceNmEUPzyiNXVQgPhC
OCgseT1uUNajxeF4pIP9kNK+qiM04Jr4H4o6YKorAZ+TKS3Hk53Urb8e7Fid+EIozoXTqm3mCfop
+3fUJph7FoZBIAF37xRVMF2waOCyA54vqx5CHUg7GyeuHaX+UYld40zQ+OWhbGTC84gXvNFpQQ6L
StWweZFIXr5jYqAJGi1hd+KK75w8ynKtKp7J564fHXnupHWE8fVNxfWpJ5pcYfHh6RL7G+sKxedg
ELGie6MEYQMj205Wqt8+lexcYbO1Trspx9qTyoyh5Y75vNYnxf2+K0vnlFIBhYrbi4/Y9rnI5shk
W8NdlcrhzOR9thRDacmSNG+XNOg9pOZj7qNKseE7JusLrqzhOWfWO7BmyC9uKnyMpCSojlO+s/7a
jy7vjBuNdksc8Tf3KuGH4+40q3hoowkEw432pxVQw1Awv4c50dwYeekRGhRwQi73DCD4NhyXucy1
RplhDmti/NGiPAI5W53pWDxGlfyFZMaKwgzzXcK8TBNpYb3E9LtD2QOItihHHql9061yu5Er04cW
NUu7nxH+2whxxIF1gEEKefaEyHW8A2Ct2lsONspSR65o5vPo9iW8+tqkL+Y/sXd33Sh8B4K2dWpY
KlY//+1MBVm3D1jar+Xv7PCrbJx36WC4lbPCnlVLi6/wpCwbBrewIlbM+xcYRjDgikK+yeC6SvqS
Slf2voizMAUC1LU+91z3kAYyuEYOGsKH9o6NBzF5cNrwi7MMj0X/khu89//9JXJOMqpztkMx+rfO
04vPA2hKHOZZVofo4gws1PM3nUT6f/nVGXBQNQqW03012rdfoRrMsstq/wfs2LLJ65jHHWhWfz8f
CRxZiTUk2o4Qfkn8z3KptetI8yfQdOOlzh7XhM6rKz67symGEQiuy6CM8nVdFhI1nhKpVqYN7jrs
AiNpiBKOxqRtBK/fWFEJ1Ln8kmpJaF4YTmQmsRKE64paH/60HVLVV4KGQYFuKq5s0XpR3eHdq4zS
DKnr4Rq1wstaOzgs1whbxV9x4xvCEfvia1CyxqEd1lFzlOTO/TKPVkm0oE0vDJZOvbyq1oBbuqYM
YZdENFrdHQegitNJYsqIWNdz42gGwS0fdzntXcaB3xg0H5FIHzJR5K1P8nxp76W/jFs+BB6H6i8M
Yx1bvLtKtCiKvnCUv/azZbvtUVJxG+LB1qn0QfV0JhdZwDIQEvZirhPnQ3cMgAjT0lh5g1Rugn04
fqxK9Qv/LdQvoG/T5wJHmWWyJKOzkldghm2BZTx7Gks5HlTiXX/GZzoohi6rlMpCjv86+T3SVpCk
9N6OlYu0zzQWNkEUHBXenaBPIXWxZT5/9suj+YT5/RpZ3O9LxMjCqWJMR0biUA+CljOBKC12ySE0
1luqRG/6PhUut7HgtazKEr/thWT8IQpa/zttRv9lNToFYDqWLTVvGtBsWOLRC2yQRVRWRG7KoQ/a
n+9i1vyGgKVaKN1o0s7BOWoYAz8qJ4bnm1oKkHG+ue7UkWXFxr/sCmJhsC/P9g0I/FrMau2/IpvZ
ftPobCN9hTrAi/nf2nrlI8+z0spRSAzLWjQP++phWoPEZIFMJ79ds06P7cL7sdjMgC5YLGwl/LCv
E4PmwBq/eP+TQkrWuhZ+SLJ/6Vb/ORBM1ntWlhg0DysxhuFXxWoAU0LBUItvpy3nk5ubhi89e6bN
nYufFua2U0Acve3QUzDnggNUvCElzNH3B31gZFZiyszA0XBGIx19ZsWjMuZR4Uvh5tIjBsEnKfl2
BEzhDx+zFGt2JkajhOAVZPNKZnTbSOBOp2/47EccLC+U1o6FRR393+DJwTonGJU80uQrQB3edafJ
0fmtec5he65tof+ffILYWNKFDKbglzIoiFMFWKjgJPYDhVqGGCmQ+6kdL1CangUWFpNzVLTVDnHH
vPFOEE8L+tQj2kKL/8WOqFdSQN1oLPeiAT1im4VGAqmU6ypOwLOUrGkkonr+bNApigThrwqTzYSH
L48a4j2XT6OIVA29XYwyfccI4CuQVDmHUCjF83B2rV3cfUOH49Hu0BR+s1SR6zHh0CxdNEJh51PP
c2Mebs2vSPsXBtmphFi7UVQtywwuYJS4AU7L7/FRrBQaAu/fntrfwwmCn8sqnn8uJR1HhR46n2vP
X17HpfHDyyN6XSm6CY2Yu6kdW4nNktXZ+/VVT9m/Q9lp76JuW/v6aBzZGWYmgRs/WWOuFVzovc9/
Khr3hv3/MSUHrGzhxeAlBx/W3P8YW5jzST8AQaiK7bTQ45ekpyJDzWf+pe5zvn3j73cYcIlD6YHe
yl6CzDwxK0RsmufvazgHg5lUsrq65VrFcOj3RSV1CMCAqBt/hPDSUnX685brjkePvwOd7ymMqSgn
PNrNy63K8BTFXTDQ2bbUEwejAoJfWjfqTLB+f1iUg6NdBVYbH2tTmaxhOOUaGoT/sgWZI7f5lrn9
gQR4pc3Lb17e+UkFkUm3fGCKBctOeulRP+x9irMuX7IHjYISb8EMVoTE6QleDqEZogi3TT1+tA6B
QORF4VFQeCj0Uzk4+8SffCnNMyYZYKGtGEzVGvVkrLVQXU6WSaKqhOkRRJ4aMEHRn8eyRLC+ZabR
GXFxqzTcgCpkyqb3DkPfQYNrxwF45i1KUK6is3/TwbugnCQKCu5MR9dgzK6Szj1f9+5RkKTOLM1k
MSGqkW72fZV/C/wc8jU7PSeD635zssurz2VAIokc2G6Qj2f9tqfe56mLk6xcVZV3HbwLW8PJ3FAc
lQWThcAGXSnnQL50W88qdpUN62O/bJlvQDYzLmiaw/A9N4cKqN5e/+bA/kbiJ296gQ+o5m9BpUVD
deF6+Z+p16sk0sGabegbm8xnLsYYB0rofpJE9B7uNezMrf6+CBQ5ZU9wB1GQD3MOe1wFtqwGnbK2
a6u+6BYKI4mEh1IIvHYmqtiixRo4VYmH3sC99Mwk4Y5wvjYqNCOpok+9zk2cKRgbsNgIqYNKEx9F
xUXnuIbgieVAKSZ+CtpklsiYV23+XjeQWNt+FsV8qjR77OH4t4GlebpNpiaZWdCSkAk007zm9wSL
TIDPEfCZGtpsF+ninudmXWCLxcRcmCHcxrY7maF8iNjTCGRr/lKaSlj/J7rJK7xVIMaFwGJ+mFiC
mLsjniL4sqvfjYs/dlVrAHZ4R21BnSwyMRklnYL9/vwftEhxby/o1eA0ErzjpxWWX5ccQgPs2t3c
kciHoN9r46dbkJ3g6NWwwZXTmC8Sk+JmsxjYISIF7aDxtp0al39nDqVprxBhCvsv23PR3mHnrxes
buuR4sQxlIHEprj5X3GgjohSppwHtSHGMgARb95q7ULcNDE4V+CmR51XIS1M34NJMblQHftXDCcM
Ekz06n7g7biRqKpzpw9U0NAG1BF5vbMGcWEIHoM8o+Ab0mnbavszB27pjwYMFAoYe1g2EHdxnp28
YCXvYG7r6QHf2J0oU3E44DyJw9MlHZgIdbV0hb3Gc1760e9bczplcDNCDjkvdjii+GU4tuzgNUJg
djktkRZqgajJoNCmA6yFXoiATPu4111oo8RgFUnOzIa+ynbrkR8pDGsUoxkDBbz3nrQovChbTi6p
3je6z18ssbuhImKrhZN3wAqWOZ3B6YMofzqVi1xuKRKvJAUg2ZWQZQhNQhz2Km4jUY6oc/z19fHq
Zr2pv7Bxh5QxX8IDQX2eEMgTwWwN86c7hcGhrP9VyqrERSeLr3Ro+2aSCEIPFF46Rwj2m1tMcMM6
U3mULn5NvMWcKLdgQ2FwXuG2wCPQcNQf2Nld3tinI/ywdfd8o8be3UsTL8VjwxpGjAzjXLuRQeyG
yPI1C23y6a3fSGhsghTZWA66jBPgHRFBZFpGPO9h/ZP/WVnQsxBX0Cl56uS7zFW8UXoJxNtXAilX
DeZ/3r3BmS5ohXCWGpqZARsbsIB30Cmg3ZpI5F+/l6I6t5Nesiu2DdIZke694V1K1yufvmmLj2z7
MPlY/KzNaJW5tN7n2ZSMzSaWrTpnmklRqlnmTX0flka5BHAFbyY5+J9J1cPoIHoK6lTyW9la9eD0
KEIhQyJ7SFLF+q2D3h4dEuS5Lebo2VVH/dr8M6I9S6Ket9g+UqI8cl3tfed0Sg8iII4VRIzKg4KN
yLGau4VFtNLAV+alYToaWmmx1143trqQhas/BNq7MnvwWBsvwzlNVnUesWjsoVHI1bUIvS53PrRp
UHzUL0JJv2yXQKWFOYVTeP5eMZ1b8VXC+ZoGaQjV6Rrhtis/BH3IORjHxbhSjMc2U589WSA6wu5Z
obpFFcr3YNFDthmCXuOPfXMY0XfaFOpp7QiFHqTQwdowvmSbYyk+iCiw1apa+QAM8a3bFpvq1axI
uLNBH602IXfoS3tZh4m8zsYd/QeY3hCrDz9idprg89xp6PkMkWD4G22VkLEmP+EFqXXjDdK0Zqgk
nNaUEE22iZchFnlYEGr1kTJ1vqVuUEehjG9x5nvSP/tr3g3WCtP+AbbnWD2XNRoOXChrKxvAOal2
9S9R2qh2RAIKT2My88NkKYpz2jkfVRza5tp5jYbHgTpnMqcesHXcVqnm9ZWU/TvCDcRQvDiYzKWg
x7ArodPZKWxlCm6DYFRFCcuLOhynnvPbPPEJiLNhm9drTvEI3DkYUweLlbvSOgvpZylzIqIrXSQ+
cjGKzMZGD5w1VxUOx+N+nsSVuqp25jQJ69rBIpOGIiHRcltMNjepUnwYR8/Z40JDTvbh12TXFN+8
Uz8541x1uXNTbtGr9O1SFq+w8YSrb3u3iiBn0fhKRokz45R1eCeYyBrv01Tb/cRyaiwceZ3M6xln
v+OjXzW+Oojb1FD8GLgCf0Xi7ZU1Unn67u17ZDAWrZY3q77q6Tn72zWMtwX3+XDnzxIsuouXI8vQ
Fc6JZQRjxcvvhqUR2F8hR9BppU03I7pv9AuETZQDfPPrmu/XCfe5doYoLJj48tOSeQaTY6Q/rSdE
TMv08NSE2tOzONHoEqrA0VITlKt23V0RvjIR05uQOJRoOYKv4StjtswSkjk4C+WhgAE31E8GolWH
g1hRj9W8r8e8Ei31jjdBU/KqFg1XS2Cp78gWXbriVldn75+6EurzzcGGP+LxAHXLOjI0kmzVWzbe
FNVyYX5pJhwjgGeeK8ahHnA4ihowtRdMY8Za5jjEu1MgQQ8Rj/+oNw1M3Am49coIrLQMM1KrjqXm
c7dvwqKdo5FHCm/Yn39UdSizFi8fu6sHVkDPlx0w76pNrLJu7rZ59WwgJ5x0VN4rDFJTcKDPl3xJ
yy6fQeCB2bd9ZMI4Gpw9+Iszm3y4hsUiC62BnY+OLX6TUxaI1CalRFdGEG7J5rqRd181yBK2Ykxc
Ygq6Jn5oazvlqhmJ2FHcmJK9P6exuGZPiOAdS1ZKWK2u3QwSZevBE4y40yrF2GlZsun63bhbP+qm
epaMFBaNZmEXAXH4BOOhSb89v7ZLXpwxDGviBMegAOmxh4WCQ/Qn0DnAiEpl3rnjFnZWbZ3jgwMR
v8e4PzkzC9kAI99T7zn0jVZBYrsvvMEgiiXLtMmX4+DDUp88H8CHl5Y5+R0m9Eb/D7Vy/PUwEjY4
ODvNJeLo49b+tqxShyJLT90CDNDljPHs6NRWD1vJrxm0czKS7ZAwpcUHkVsr808S/eLhCtaTHM9F
k8ifxRzE0ulEFyMXXEc0Z/BiKiR/cGBgDgcCCzU3uxc38Yo/vqyHtCwZShgg1Sf/sMIUoIafmOAy
z6rVBH+OVdbL3IjhbpDoef8URI4INDBwBvBc95dOwGqSPyOtTINF1DeJa/Ln+/q5RJ7CA+G8sfb2
MIPiL/blTJw2tZJ0MqfHy48n7OfozChO30RP7hcA3F+4Fh3QA7Eq5RABQboLBgMXaezfX3vNW3E2
7md0DMfAuqLhjhPGgPky91eWnfJoTdQWlmRuPRXDcQY5BNsZV6hLqIDtWe3Sz0jT5tYNY9BqcWih
W/Jc2casDBPLGaQwOPwjolAvin0iAfS8qkUeL0yJ9iF5sFtmtWa2R+/5vo0lzE0VErTT9qMat7Xe
h+SVWRhxfpMhBkCgDtzuzVuE62wTgOl3wqrFOLkkcRqfN22ozCDXBKgZcj7isZBbGuv9fkHCUyXz
McymvzgpDQ2ak9kVbD1082CU1DnFdx6c7u2FI83Po65X9NqIWYcA41ObYOj77kaoV0+TyopFZRTm
yslJTRW9ta9dlLep1878PgibHGIZjn7zgTBGTKmB64ohifj8mQtSucTW1QGbE6KX09up0BUOo8Lz
eHLQiOZRMtlg8f32P5CW5V9IsFd6HOM89GROPuIJ516DEUSyhxLjQ3/3J51Tc+mJpCUj3SpxDd+r
ix+DZoUoE2ieBRAArdLNXpnn1j8025nX/Mk8ubFzswQAmKOJtPckEkweIJT0fFkqFBHtWXUpoz3y
/qzr3INLgUjkI3eX3ATwDLnMEKeHujnAvhT5DDYQHibhZfwbwCegCS+xf4/kFUO2FUNsQQPWStR5
cE5FEWsRtwFZpTpX7j7XYaFRYSHpKe7+ZANTIGHCc1MJa4HgUJVp1dsBrz3eNGhDTeSiuIGhiTDh
pramBFLh0rgAlhEy+AbrckQO4rCrLa4G94sbGpBVVXnMXYSfe0k/OksvJfeZ44h0tk3fCwIEYAtr
ZWlEmcf1j8dR27a9WBfzjOwZBHgXeDiaqObWehNJ/JNmcrP1jUmhG4aWGg9Pt4ZBDQSUIJb4RNpv
MP0JpD4dypKb0/RtEcOUV024m39XaGF7K5ERMcXzC1J7NpuGIQXJ00wrjIQS/4M+E7I6FU6SCb7s
hO70x9QJ+WOIWJgCTnJUfkGaGCCigaU/JyNFD/mZQfR9IgSFQpqb0jHLp4hK5D9JqMgoGkKsE55O
KJrPnk8RucEskqavrP1JViU99FCjbHTG3EY1mCamPfZF0+B3mRrWiDC0Ljbsc4cGqvtRT6Sg71uv
oPSYMtcZeu8PSwmvVkwZxqLZ8ZZ27ZSPEUwHKekK277GCDPoZxMWqMG2oPij+Whv0+d4YBdmYiXh
DoEg9Uc3oCkJi+rOEcbuPD6BqDedC01PeNSBZ8A1lF0UrqsFVD6/N7iw9Epkt6TB/dd9Q7yeVvLa
8RbJDgqw7uHXyzn4FLuREKiQVlT59FX529FFRyRY/zfauQ/ZugBdLzdj5PNWk4UZw/iHaCT1EOVO
56Uc5X3MHq0NeZC8sS8IdfLHmI/ttQOKuiMT/FkK1CY+IW8QsTuIMkQQhXSsSDj2+pKcHJrMc3Xc
2o3Efc+GYF8PQecakGUvaHZ5FqayNdYrunLLg66+LZ6r3o4G1+Gkwi+1Sls3mcnz88WtEQzFk+Fe
Axlj5UxItBr63Cn+E1gHPNQQbWxl5N/3qGzuus+K+XU0YZOey+RQm35OnR8HCTglt4A7RQg8Zpt+
nQF89vJrH4WJgFCmnHQC6o7Fb5lorc1aC8nqdliplU0vRnr6WgKCj4VUzfc4u52KCZ4ILFb1EYJ/
C6PeT1qon+T73d5ZKcKS0KOFgB5uTZhkC74AONjRriHysSavfp2AttfP2EsBEN3f6g6TfKX3TfSc
ZK68x0W3+hHZyluSTReKRemP0QAcdvz2lJ9/kXOnqTl7xYhnt5nnlMxg5odibSXQzo0qJk/vq7N8
iCf7si5+M5pb0o0touIqXL/qxbi5hM49/r+6vCyl5TkEn4/eGLhYZKl1o/WTnsdC0p/GEjfYz2vC
FAC7jePQcKbtcqBKgOpjzaVcz7VSa6D0xrtiSwNi+vN77eb0na+5LYZzd3Pn6kk2uhfz/krbe1wB
baVtLSYi2RyIdauhBVtqJkeYDsQQz9hB3+ujb4exZwnSJ6AJ2s2M762Aw+MAnhNTKihSwgiboTar
oQqUzee2EE7MBhKYdhEp637rHskwyTzn6rRPcOFmGxDu5rrTUEjA3icZWODnSjQChHN3seA/MJK0
ymqDf3AOol8C0U5Ajwzq7b3Am5IpCcu2/CaC/OV0uzIDLHQOXIrWxqi6cLhLTWImzSVFoJ+uc+NH
A75cp2FO8s6wCm0aQj/q/8+bSIsyaTo6r9m2eDkhehq6UWeo3yVK3dkvQdQCe08ngmEyIIAGzbdF
dYXJMEjJ4jr7q94pDlvxINFE+bAZFmGAnQPW+g67yIP5t0SlnjaI1f3Ty9wjuAcM2h837lLi7uQB
B5x/IJJkPF1jaU2ZiknZOQxvJ34fQrVVPk1qfyaBN553joaWFosUjO+WHcEq8xiKeWbYNuGnh6vC
7S9YQA4pWLi8/8g3Yg5NrwLa6aiogr5UlVSqlgso+DqZBoYjJ/C/6D9MSuMbTfpIk1C0sVpqILVE
zlhzR6oJ1t7md/1dkZNCBl8uCvXOR8Bo5I7dpfKo5MEwRcvm9auV0yzZ9KPAUmyPmk7OJU15gDrM
1SgyseCn1XE9E7q+LfXU1ANvXnzEceE7wCAXyYwBw+pXmN1c+Bu0MaYweDbNYD+jJITc3nPy1rjT
nNXSUfOe08cUaw0jcojRt3F+wo50og48DTiHdcedRnYUZCWuu6qm6Q3EwQrSRouKoOYyHSAp4FO6
k6hSwuYd100picYe8XaQqeEO/UEu3+T2OfLguAzWtYD5e1wCDrRtl7xp6DqFCk68+MkIkppNoEyH
2lj+S+Uzi+ckamyxCJ/K6D6w/LeLVl1uNycouA5pCAgeXoNqcKsiceEdnEUWeF72r/rhd2Rpekq5
w7MA4vMRl3riuidbxFMSzm727GMtrTbLWzdbe0bHO1BdaeUWlPqihqBD9kZQXFzWALFSwfuW9KOZ
AlyK8ylOUEtGZn39bJ2pmPrLYyXNI7kBn1t+VGWwkXnt+B2uCnCMCdGTd+GA00nvpQ20iLKXFqNO
h92+4cHl/9TPt6RaP2W+ka5VBNLChTLRORCSHW5bSguqpUw8IT6x/RR06CSt3LHaZqprWau0PvqA
burFaWIM0NXaCeS1YFQQB1KWQcnu4u2g7mMgaq+zzn4hGAXCBoXMkXjAvDdsmS/Te2OOaJ6PaTRP
iXyVXG68p7lXsqBIgrlUWHou4UUUoayDUXt1gEXSIP0xjXdEi1jrCFRlDEjhizSPxqVbu7fEr6ew
5l1w4BGUrpR7K4pM7KJKxvGn6bZn7lmU0HT7uVzFpzbfYYZ/mJHS8ORb1kEwCwEitoNO2kqaWQVS
lNyHemUsC6pSizaXd2N/O27ojFsNkddfS/lzhEf1rifUtWHHrWIbVlEdtfWNILg2CTx3xSwBS0EA
37Y7piMqQdNjeHdIj0ydBUCtIIySLHZbDoEyGJJBL90fi64q+TeB2QlLtLeFrX/4Q+BKz37TzdDq
Dmqx9vkKvr5MR/sZnbhiJ5KzdPo6eI9V0cHXqtx1qeAelSqj9ywPnNiYdfokUDIuqHoX5cH5JUvW
ojkxIayRkuVuxFj5AlRjHxHMR2qNmcu80CPAfk8YX6+yBLaF7U0NVgfuU6d+fGNmLkokZcOLMPrQ
r/IcL6PwCkbDBvbXm7akh7AzVIUvgAm8G+8KfNOv+mu3ZKFIzUzimKI9YbLDx2irKeQx0z7SFJi/
5J6Fc1ykjm9QzoZvyuDdFi6oPGF7cYF3GBKAqyPA59aNzKB1BmaxXAn24YGr5F7n16pE5YafbkiS
Jc6UAAJY6NZQTd6BwmpRYURJpRVVoKkimNQuCfEEWqwtzbzMzoODM8MWYgjljKwzzCCJR+/O0qFV
7eJFGj4aZDrapNb3guaEMEzB8jrJUr6r4RFOZoTnPs22fpybb8TbkDYsbEjjHCdMwNDNfIl0muvy
IJxvcEY9xcjTL5MmVhChMhSMHm1my3gVY78bzQmX6kIWgd6FPvLo61btFv6wYg86gr6NfrtMhVRd
dezIDsMTlYv2/f6arE+pX9Wg8sE9iG60rkauUJEu6OyTBvYhm+5SYRHrw9u5QirA2/fzIooNo0kY
iLJZhVGkr8cgUfW72LQiWiCAmpsmBZ65DP5EEuEJsYIpydWxN8ybAlUiyh+CS9bzGmLZCrowDquj
CcYKkIZ9hB9+3qVmleLWwWt3BlfYy19B0KsmZbtS5b6saH4MTSg5BGWXoML8eg9Q28z5r1U4pVq2
SdcdOGzwrXASaRGZQ4KTNkHPiNAmnRkaoRp8eDAllhz6rxPMwLxnx98+Dy6wUqO4eI+Pe033Ppx4
bItK3FLtYp1masOYJcSJawZDqsf2Vy51x3UWdn8fZFfxxhLzDqG3EXkAJCfcQgowp8mMTx/xTsaE
/LycLtB6F34mcMnh7xuQluOBXCX6W1CHFWNvtWzeUX3p8Vd/KY2zhs0Kfein2hSy9ou3r6bTNOFo
i0E6QEUgY9x1nZ2yHCqvRPniaWNBjVXzjXZe+HmJmMBGDHp3FUgvgPrAGVuAu4z5bMOiapJ3vMwV
9prASzB/t47hg6KFnJfRKUvXL9ZKXoFkH2y2zccDv6+FBvKy8Zfh2H7ja77RECOSoIOgf5ON+1vi
rf0c/qBv5Y3qj/6vbsjcLO8XYTtdDlV5kmuerw4z/4x/rUAJ7M1Q6XgNS6ZC+OfHcyat0A1JZz5M
o/CgLfUcz9oyJQ8U7W3MWWgAw1I0za+uYpeatcKlAB64UbUAF4ftaxoL7/nsoiv6fnJfX2TMVmYv
QOVEGGBLcwPdkawerYp34N1xS1UtgzwUGxcFysOK+rKLydVUzj6DDHLoX1zjA1NKZrenmOg3qa3a
vmAVtyKAlO9vkOTWcALmq+iMDmssJwEWYAlPRdHGzY0RGCktjssQV3WZau/mSiVLwMYYb2v5Icke
9EZCNa8pmAwj8mNcGRKUSVWlGPUDEX0Frb1w4nCarU16RTKekcEbgMu3WQwQBLFZfshCtD1psvhA
TF4srfa7sorqC/qwAgY6rQXuvV0smyNcIcMXLJGjtczXYaqcf+M8uU0L7s9TY2aJNSYF4dgEwSh4
Inea4DsrqC7UfyWEYRez6TFvOj6gr6qYgI2ibLKpC/AE+3pX/UEHjA5udmHfGuSQFXnpZAbg05X4
GJ67hPZh/yiwgR2jZu6GZfvH/oRz00jLsPOP/DTyOrIdexBG1dX8EczDnm1Xuxjel+sttFgMy6Wi
dmKsAFX/A5em0F8HQLg7EoV7fDaEvkEyxzSqNRNobCqGuJAThFRR8KJDDwPCg8Wz37oftofNKbeU
Rj+dJ0fGdLB6DVi1Pa/Z/9QQC1Jo1qizfIvnM/3kPXe9ZOfA49yp8a/qgQi4SWqxm+wvhaV3C4xR
+m4LDgLOKIQO2BWRfSuxRuKcRBttbpKWGRtPV6S1Tax/pUMWaGpELhBa5a9vGaRmRKfJQL0jZxLy
0OcyD6jDrnYQDHbge0HawKwdbkx6aT5H+FDtot1EvtuJYGEWjpWBbAWjxqar/QErbj3QojdJcFIf
Zax8Nssg00Bu7RBCtyFD2Gg9Ht+sB0D3rzsbo/CQwFaCJJRrdesyVvjfXgc5kezSiLp07+xVtanF
b3e23xoKMU60NDhhcAX57AByEeFI9NUQX0Q3q+tDeZeAv/CR2apl/wM5kjdQc7QSd8y95HwChKnf
dPlJPlfIW20B+uLMA6gF+BJjq41J/PD6jY2XK4ppXGoM47P93UPuLF9OL/Wi8bX6IPRhkQXKwts3
DBXk3XIc/hI3OAbexHNJj65cBUncE5MhOXxFrI6WbTwAZH7p0vtnNNg0BUC9NMjPqpFDEdku6k5s
F8ZKTrHhCzD539xdw8EmE2Qrf79w6/fty5vmA8R8eTBOBf5kQrdcOjU6ylOn6ztUINIxMMAHIkwZ
jvDLIZLXC4zOkI3e4S+SnqpMEBR/W5EWTGqU9YRHmUzOV4jwHlFLm9OKslbnKHbaXmobDiyePmDY
4clPVlSdHLxEKBThDPOwm9a6TkqzZ2cx2zyvzbxJ7UZQK/hg2gbF4rjHnfP+0Vfjyo4rInLEa6z8
odr/JeWLa8zznPipEPKKlP5uaE0gkNL82qKELezsdS9g+nFTxGwLJXq/aGe/ibNzeNmQVXwdNYvD
y3/F2qaZr9B60XD7iVDjZ0QcooA3dwcrFst2Wjp/IK9vEPgsBr1m6nSCbjSnw9rcw6mvzT/JTqyc
Oqvnj3CvwJE/QYXHwBgOUE2j6Q2rUP4mHy43rd3INb3u001eAamWAAyi1sbA3SPu/ymHxAmMqRkU
phia6C8JNNKzEfWxmc4NAuH6MOU0Vrj8DX5vYZZmpDuweCNhYqZntzzWBJe5wC15k0zGyGBPdj7s
mZ2HnqGQIpaJU8872SoW6inIIWvbEbjNtXJOodQyC5cjtX9X3dOW3LmHXREVhxh4o42aSF3ycGfy
Or2uwOKDPhyFUlsCiyeUVLVyGq+WEnthMy6DwfT/gHCtoG2hwo1IpZq9Qkz+PDjMvBF38UOQ7t1V
YMzk9IbxHZuhGw7KUXiakICdfnPrnB7S5U4AOksnbl0OOpPbvOrMYzi1/CIvpUJmX1rBvJRF1UM7
7e1+vlBy+Y+QXjjjbEVneqSeQUKv+Y4JpbSLddmS8gfTwuTTqJS/r67lUDn4EXS/RZwUZLRLGXi5
U5bIs2KuRbYYa+Po0vqN4QJSeNNUcN3/C/8Z33BYbMaEsYgid0nSQqOkmJmeDR0qabDZQCfqCX2l
Z2ubwVu9K0Xbg4OsL+mCvo3gzDxVWZmtW/NAz3tl8AH1OcTY284AnXGdaSLVIAAfsbzipaghA/fA
8aBsRtsrckUG37CP/lT95hmqvtNUS8rvm/5L54WaSXZrQEwMGq1ESoudNW+ydH3IvPetcEsauH/I
sNV/UR1UYgDqCV+wpqbUjLrbOEVfAzV8kY6KTZdb/AkW8TQo14isU9E4RsO05mQhA4UJzIgeM9vb
2P19g6ZZtaeWJ8tZYtOmh6H7gGvccihMrEkJmmwhUB2R4IzcVpiV8ExUlAm5rxdh8yjvZMqA6bda
nz6asSsZyPJ+NUVV2UnIwP8C3RvTF0nfiY3BpuIUjwcojJ08Nb5vnY/+71SvdxLcvE9RNSPVS4TN
MJVyGqupuP3OhNfw51IPZsJPUpPGXRr00ghRzsf9xRqAD3t/79k08cJqZQlwFFHdXVcQD9E7+nmQ
Q3S4gRbsP0qu/ma2yEKNF2oiNZPpnCt/MEgwKHh80iAZPQxh1Dh9qJjYFEJG5unZs9rEzubgEYyX
nOJF6NCEvmJsovPBlkXODgMycseB3nxUIldIjJSnxp/he5I/3PWCnH9/c75ml9MRN84pyQbwLKtU
UZ43mzWjEzzjt+UTG4Aftk61gN0GuzGVTLesyp9/kg2ZBIxvszsGDfiHbswpqFsNuvUHlAkGf5LG
hesk7IEFDPl4aZL25GutpgsGanBQDoxkYtSop3j09yAUusTw+ogyFxAkygr5egG7CjZjxvVdw56X
OA9CZbwBkjMMLFczZgwmDxRlKQrWOsqL1G88x3e9jIPQ/iaVOer9Tn9pyW1PbjLuYwR8F01d3cP5
U2hEGZ2NmX7eDXroef5iJrlYyxKT3Hc2PYMYU6L5FB1ajBXnQMGQU4brQMq72lMlOCDUGf5440Je
zJ5z+sulBdHDx3FoY4jBL18NmmxTIA53WmBjOpfevIOyhTwP2LLbT+8jCUdb3lr2p2hMTcMjwsOg
sythIVdyAyugCczqiE2Oh2OtGldayYiP7T7kc2X1ecP+1UqxBSeP5fXy+GvFkRmlUa/n2wVey9Nt
H4avGUP2c0QRge5bLU8mIb31JX0n+r2c0GNxFAQcomxBi87HB0+IVpWhkc/qPxZUcNUw6P2zFzHv
7YTo6pr4T/5zbzM9WqxbMHS7xXqV2PCkNBk5RxbpM6vlLV4KrLm+hazyGhau0tlvZirq3g8XXBcZ
EsbCUUoaVqVSC810U1dhDgQJNMTqWbcbJRBluyz5114DxfqB+4xDiv5xfYkYJWTYDPtcCxVLbps9
lS772+alHcYVNcMzysC5Y6QR1g+5nsbSLrzKqx3gudOm8mwvElQ3hCHuhpynrcCj3bIc2csg8o0V
Zsg3NdIVmm9QYjl3Fvy8K+4pVJaCX2wlbStKIoQ1PA7rvL5RhZfCwBMuFFT+WKtXf3gOu1LetkfO
X9Q6tRpazFNj4gs2mBAWJd5cpZC6JWk9tWOZWSbFggKg+aPoDhbZNjvKfNhwc5KWsPvn/iA/YC8Z
skYBfMdL7UB7Vn2oGOy1sGJuEbHB6S4hkiRN60WfzQ+Y4IY0mSiSp1VVC6MIsKh6hZUuJSYxdkM8
4zYKK+ul75lOFNGx59Fv6V7/I0/QezK4KDZbnC0TLLw2aoSOnroEDCpPJvGS4jK3KPae6vw/ZKy2
3mkYbq6BGvA1i8P7siUdwcb0c6zsIrs8FrFTD9HfuQdh+YTNRMOyJS2v7OG+F23rSIgTeLnAuf6m
l7oWisyyJU8ffhZi2zwpVN9Sr2O/OovARjj0XTjDHbZCQYnPfP4UuviG0jdPyzQExKz9eWuIDfSe
M1pAc1428Ef824ISW25wz5MyxDSqZCF1NbbKYaeoEEsABUxOsWxMqCgIvYfJdY6xUJBMd0McIDDB
kQEKq99G7rkWmJguVbde4cZiDYknhTRMTfbQF4lFa4oib6csn648VTwgtUG5PTm9N0jFZkaRX3um
njBAlrW2lq4a+GjtYw8XLmjNtEzt/i7Dit2En8RUHL15TxweVC6D5G6h8k0x9N7AMIITsHU29ctM
scPJul53RpTOoWYyc0wuKxIncSNEJUJySlQE0x60FrGL7sCmEJJs7nS2M2y5nyVjNaLEyWijykfy
0UBzY2xhZuIGhdy1GGo95YDsghEj7SzboSnQzxMDkGbN2/NmmcYvKFn9l8gAvElkseT8ONtEp2z2
FAgkKN+lPItI+HYlMDwE3XZ8oyKrITzQASIbNz4FGwzQsXJuS0blQrG1KP26WC1nsvJ8qZom3qXo
tF+1ikP221NMPBLaMiaVlR2L40qn5nzDkDALEjSDFo/+CDXTqxCUZsG5+3dHuBa7zwEkRw+0ILg2
0B0nXlZeT/hJjRvKe1yIm7eJKRdZkdVyEze+Lr3VjlZ7a5CcVes7AA77fsChtYVP7a84PEAqwOX/
xncyF8s3/AZK8mv8ouMJtBqxBWBnNkHDwWMLEBaAadu74Dd/l+C4iBgu8/6lcZez844ojrWRnptK
q+lrVGU78QbwjUvNV2dLJ6mcoQZbvmo8ZOh0nFXJNb+Kj1tD2UFeXSfrcQnWOKWV9JcN4tL1X6VX
Ab2AEA7g7MyFhPJ8LRu4JU8HIs1uPZmRzP6PS7DLZLJef3QLGTb5Yur68T+7S7BgOYhhld9rqjnO
N9nWh2C3k8euH2UpDE2YJe8UX3WbCjND6xCFaLGgmJwFXzPdTE5sFc6IxV5jwLXFD0RXQJqLGn9B
8ocmLALzhExqxUa3zawLqb/73QehDa89P1JW13hHCBoeTDVsrU7HdXlX3EM3ThqdK8kQfo+1K1+F
tz4UUvZGcv2z98rpUK1NG5xTiMI+xvIAYmEKCkIu8B3gmU4J6GBdegcedPO7D/kcWrbyx3U+Kasj
h4n0aXXKSgmfwIV9tekrJ7j5HSQG39f5putbPwHHi11U8PxguaDb5ahRxhsCDtTNOFieodMrciOg
C2D2vYwgaCYgYQS0LpLZ/Z8k5bLrfvFvrRGmZbTe9+O7tAOmDlcE6/wihGdG6i/dMSH+Da64/Wu8
mTmPFMx6T0L6qgh7C7LXM437/qK3FkBdjTX7eNMaJu9yeduTIEZ+WvOfkBoiEgyBgvpcfrqXeQkh
sM00+lI+RuFJ1MLveJazhSQ51xF/jsTLjLkBMQOUE7Djj9MgwjQsedI8Vr6xadvsrq9lg7ONEABj
5Q76KJuckRfymcLyva10Ph8nvVR3RG419s4T1OsE9LB8zbknBjT317jHZmZZ9pYeThFYkFNFTfqh
ZhEuVhFvsQC1zbs+yXaVMmHcrdZFsn9LsSMPyh60YQ/upRQGNY5iEhfl45T6ho5Bns70+GVwH8mz
oFzS/2c1DlygKusHAWwpi8N/GrhaQznZRxzPt/J59Np7KJBG2TwcyU52wKskbLn3twzhP5/BWL0R
PzrWkNEo/v6IE246V8SAYdTi7XB5eJkNBQX+Hts61ODx+d9wBEqdvlK74NCnhbmJJYYuQLcLp+GK
i0d/eX0m1AgnvHWDGYynXV9B/LAOMIXC0eKQGGjGzT2W8l434SJiZP/MOH3TODsMtRUQShPCe1wv
ehPFaBgXDs6sUuhyfp9DFQwjOD7dfVyxiUblbguQFIQ8+5G9P07t0PB2NHwPTgsqNUkfPh19nOi7
Hf0+a0cpMvu/tkeDOsm8wuTuGKuYz6/g49qwlnGMb8DuUZGNoODQiRPq7wWItRhov2za2GGWiM0d
O+HDRGvWSJ8eB1avpEH4iw7Md3+cm7RmnIXgllWswhheSEvF0skp7vgzUWC2TaybwLArP3mVrXsF
pSDflwZQ7jtOzZlXygRoucCkGUZan0q7eF7USDtkza2l92a0lbcPAPNHt0i7IvVUMMMX7HrdqyY0
S+hqmTQivUtPm8AEGnijSNugyaFZMKppEmLvEzEXnS5rSP/JuuPg866wf89bUs8o6gafbXy47LQD
tlSPruTDweOyfX8/QLVOv2I0NsO0KcdKCOPRixrpXFhAcooKeQ9e2MH+nwlXUrx0otW1q4bOztk6
/3kXVmpIxT7DVU5kmVUBQXNxyCtp46+InInL76mumBX1skqrxKUE0YBN1i9OmxLjaPxG2IuV7TfD
Wi44B4NtjMIQY0bxCNwolnWrPCa0F3oNxPse2oSXbb2i2nl84xDV0XSsWs/R+Ab56MmcAHpGrW0m
sPWDEqqY84NmBFSySl2tWky8Z6fZ9/WhtKH0mdVMjBSDyu0MFiS8WJrL+txVbIXYgpgmBfG+rtKM
KwFo9KgKhx6uyC9nDH1Gece6rdEEIKNnzIgsqpv3gljU9lU16h2fvZsnA9sxJlUWdc3KdRneOWa6
auCWABWh8lsYLAVEyCMtQNvKwZSsnooKkgMGXdCiLj4ZgMiPuOBA28gLDvedDysWYJMnbBLBybIn
v18UR4MvaYB8NAxchORqRhj0vyGVWCAPyjc3fpXMWRkLnnZuj+rHDUbxOrkkgqb4PtNbXJbUXgN6
aGApPttvkdF67dvicPuQG06GOlyGJ+/NVEZyMIg1z3kVYMvuu/pGYslafWPSx2SGICL9LKAo5qC1
rnPB2V7/5aK3CbKy2YskOioe5vIlosCqtU0giBiQKc6M2/PynJv7wo/bObmZ4Q773zCTGQENogeb
TkC1plsAtawuXkqHLPl9BJWO4g30ypMoqBUKkiWBxwSEh5aP0xpvSduMVSO4XKXHDGLWTnuaCCRO
bYRQpeNt+AbwxL3FrKxLA9YCgTYjSfHsSVYdRD4ntlLKQ3EJgVAzbpg03xVp7A8OwbLbeFwekSJL
Ut5vf5E2v04YESgdRDi3DOQhFtLBhvQ4BDjcUJR2RYGrnsFwYkhzSnmGPJ8vp1vuhPgKSL0dVS8m
AC9jTWkUmZeS5RTX+y96NIQWGesOYldLFHk4BbfmPVUz2lsthT1wE+e2ze3FqprCGOOG9L3bZiIq
DOCK5mJuIh7/iQGKOARey40AtWfHDjImD9Pln660N+S9YeWC24B1m4SgA4ZCFWf6MRDxw4yKeda/
YweQGbrqZbBBT60WJ6Wu7CCWP7yrPx9w9IeLSeUAEXsyrj8GSr9QzIVCCL5uHmvASM1HzWqu2VQR
dCQEYBumZMpUSzWarMT8YRUwst6b95n3KwliH+8gRGJNmXaD34TlPhHeoXnwnQYRYW7SekutdKX9
A3d6xzVmRgFfKUG4pMkjqA/fvoSnx03DS2WSUQWdYGXW9beTHANHecCqFR9tcvf6QnK/ROjh4x/G
zZ0SBE1gokHbtescMMDMCr+EVUdasotqPWp0vLG5MhtpLhx/40EhpztdQ4O3ff9kIAPJ68LTz1sM
PFgKUj7LBasoD0KaNYuo7LyEVEYBYYE2Bpv0SoXrx+WTp9dQTB8GQcFVn7Ic4sKF/CkmvEqF3xA6
3rJEPAp893VZOToQb10L/ZJfb8A5Xxf98bbmCyyk/QjMX6IENxQ1vQGYuof0ciw2RI2cb+LJOjS8
7/CM9dRoyTqRDS8H3K7sRSWnnoDZCuD+GMSx76+dvMBtPatZ/RPkN43RVHD4tfu7MfBvAW29XCZM
fCZJU6PuwAXJHMPRO66jUOSiql9r7s2ptPq01PtuX9ts3ehcJXgl3LQIgjPyOhX4AwhjRKIFCeD2
hrtpD9FhdAGYuBFYsVBXjFqUzqrO+JQj54xzTHTPCul4p5NYbN/RuxFB7IoAPgj6wkAuy1UHwVGk
T2KjoF1/BivayiEykOOWZ4pQyRDihnbaSlzC007p0FgAKlwXSAezn6EkwFz09fSqTTv8RZVTEGT1
47zSpT8YHrC+LUvb9pZSP2W5gM20KW2C46MfkhsU7J9q4Rm5dAKwUqGHUYXWZPtGIMMyHVJ6VW7+
isbfraSGPBfs6mRhjDEedaaeIPDh0hTuVpqD1/JzQnEZuFyITILnRLNa6SzaotGDlq/r1vODT2Vu
XIZICgymv7vIupHRDZdd5Rrd4BrLVcWP6NSlAzqADBKIq64vVanA/66/0ZfynWcfF0jDB+DsAuwA
l5CzHOPzFdOnaYqOVks/myAYGrTWdjRtxL3eqiK+OjGJuCHaR+Zdrj2PN6MxplFB/LxI2SIsKvWL
0MQg8tVImDmywK7aMvLgzOtPin8v1BO+9uC7BnxAhZSp1s+rmuny8Z15K4Ysj0h7FKVCWamndit2
EarA61D/i31xv6PiJvA+1m3T62KPv4r6/4+cB8X+L735QUH/q+Cowll9JM4b4MTufbGD+BgZ0w+s
8I9E6OKpMeggsXazqUa7NWDnVZ54vGsyJBV+T/gKnCvr+6j5bzNluyihKWrid98boiMeON9izI9i
ziou7nXx/ds+EPGmzgKZ61jsEu1ZR9fVO07hcUP3Q87C5CBrYKAEMmGOGqSUYxS81b5sFdrt32m6
1m2O9HF7N+HUxKCG6hCJQoRjyLTNGLdyIHI8M5GYPnTTjKDsl3f5TUV5DZnHlJPpcDMFFP+Smmpf
Jo/I8x8aqnUSk3ZV9rn+C5XNu3yZ+PhYvRDJrBJnzVB0DrQqKCQtydPa8Vg921CDpzJuzbN6vZqp
1LkY76jrotWtBM0lbxxHY1o5hSkl5LPw0f3ytnlnji1o5D8TDeSLCofrFOyTrFkjvr9+tlOQJYtd
aYEVfCwuZi2GinSrDB4ukjxEqHVjdANfhks1ritfm3aTDxM30GnO4c48uFVzVp4fdfwM+R2qwrjP
6ZTYLKnnol10ZApMcA3y+ycO/Iz9qKW6L5RFAOSEmsjxhK4hiaHHkuOCrGpihYT/FUj9aZCvPkxI
V9UTWGEWY3/l9Gj/YjEIZZa7c74Df6LfwqIDxnq0yFmSz8Qoh6BkBgcDIaQ+2w6r2xmZMFJJd9Yd
UHcNGAcbXV0qylRFS2HAu5u8CRdskIHohfylcCSOuCKLDdkcVO0ba8ZBxQLQMCqUaUsvD+HjjSNo
uG/mjuT6p8JEEiF3a+3sF856qdsBNewklWnpRQPEhvrpzQ24KZnsGssoRyd2SxViiVU/HFkxh3KZ
PChnLAUbZY58dgzyjE5dxCJ/6h1oTxWg0XMWUtJJIB69s077vqbpsnKXVfeURZREJaB/efAS7qVV
QStiJYNzL56XoWEoicWgv1MNdr//d1Os0hzyM4ILXdIJ4hsApraf/UL/cm3hqoPZlPGLlXhDHRiR
eJ8717wHTbtSsMfy8s/RTgvEL6MrLHal4olcj3NzzQdUkzCy/xM/hlXAeptuXflpUub0taFUcBBA
jW1IBYvBLDHy5c1QIQ0xBzzXsGlznAvhzKSM5rSvCZyOfBRrzji/bmO+jAL8Zr8kSBeh9sZxL3vN
6VP4wmOCGJGtmhhlXn0VFHlrf1nttt4sh14OsDhQ6bxRtKMTMYOO1pwEw/X79f5h39mqckgwmMF4
25rThl918fzz6pqL+GRB9VjJb0Rb3qx86I7mLlPdVZeIKRtKnQbsR79A68u3mhWrQlKzAasXA2C+
CKPbNrVCLzZetM08JE3qswumZlQTINbOWmDlhXPvBGdACl6kiLYQX7kNkemiUpLKG3HOoKiQVsKl
Q64hF9ThtshE2qzZvuEaWhQBhl0WVKdJj9pDOrM4Lvs8NOKv5ODmGyKykEUFx55l84HFmXYI65RW
Vgo1iMxZWM86juZv70DcpP75j8SOJLIWPaeCEjUBoMLtKILUKxhyvo1m2Z0253p++alVf4NrBCpY
U6cPQSsQqsNtcigJRdaerbONthKMkh7nFWsYvgngmOX8hg+aX621HgLcKSXWXdGZ0vrD9cEKjoEF
Zs+NCtL2nlpRekY/CTAq95rSrBvlZvgulnbCTsGgykwO4m5nMGJIFLhBZ6u/IyASlxxi+dWWgGb9
SlrN9hfiChzrUXrhoO3IJOKUsPZwwdQaJVApk5bC1crU71pSlFDUHivYHBKSy1ghy777j+OVWqeB
jx8LeFAZz97n05BeNsfUZXq05Eh6st7KbUSc5KzOZXB6HNC3BJjIGdn3Ri9XQGfUtpqLVuxP5N3j
coIKQaM9UaOiyBlfcv8AiXGyh1PSWorkRcKJtXNTNOknujqISh0G+58fgSmx381D8mlD1zn1SkOo
Tl17L42FxamCd19SU9xCZp7j+RinBtvJZqzmwAgh8sTbYGEEGnIUVpLJzfwdW7FJVMXiUk9MOY0x
574K+WcFfCjbgWhfdMeMSCRbeZf2/KaSkXTPhZWePo0G8B0R/ze/5wqf9qw2oW+dUH0Ns75uqjQo
p8Cq8Y3TttCXKvivBq8qiMZwTAfunQ3BzInZsHIMPOiv4LKY2UhStNDw/M3VIUHsJ4m4q9k2K7PA
8lrni8RZL+Dd6Snvai7HY2RPj6PYXAUksT6gQJLveJ4bJEksmUpESmwltAB2fO3hKqauabdIriUe
2odvSCqhzeVYyFz1rWpGEk2JxZitgN9j582LbIowQlnDxXh1Lo+lJCm533b3ze6g+UU38VDvs0mh
sJ5vL6DcObm2hXFVP7KQ3xVkANKxBByH9/iSmvSA59GS9NDcEugVPPoA3Q2e3cN8PTZW6ijVDep1
Lyk0pIFespqUFf+VHGql2a50OELV0hoFV8kLOKOCi7SVXu7t7AOwmU6D0sJPsoqhJtLGOPhFCPop
2P1Hv8POytSZw872XNTmyhV38miw6HbKKwhK0JTldEDbfXl5DejnD93JBK0Vyz5F3SWhE3uuAZk9
yNi9v0DP4Rh3Tr2L5+wHqh0RMpJnJ27ysY99lJj0t0qyVS23DwLz4j9+O7rD90xjJIANpU2qlnke
n3wp7I3v/bFsq0hFrJhQtnHgdriwwbOk/o0ainzEZqMHFNX4H9OUgyMYrUSnsoCBk/MSbboVoODh
yTu/8CBTqEP+sJcQOEFNa1NvcwPPCztq4fxWCS90EMq/wm4P9eefA9miFbxKt13KhAq+hbBY6XU8
rKdiJbtcCE5b0Tt9GM1CJi+iW39gjZ/DsT6K9VQssLK52ChgtXy+U8fdeFzZJjAs9ks9jqnySxQF
3/JZCkl7X9i7BlxZ4ld3ZByO4par7ulk4xN32m89+nzSuC1fL9w6s1MUrYMyPBr52Dh1bMoM4FvD
ujKdXTgv039gNdmIUPFDwioqoU5cg1o2cluA1PKpsGHfNhMuYYAemVn/mvze6xHC/J2bovxUGQYL
kP340TQr9gIe6aWSbM1TtzDj5gGb5s/Ns7UI0mLEmgP8dLGpHAm2EbsdYCQbas7gBDS0FSV8FYWp
duOmCZeU9xbBQ/gG2fCVfllDMQlvO4YVYKSqH2JUvTXEr0+IEOfu/PUbEeBZLuJsLbBTs7G6YmFV
xA1nyaz8cfXrCj78qPOhEUfDoPXaPP3941kqpqFTA5Ozw8ynms3jehEU+MrRwwUhrgfhM8TAHh2D
LZQpxJ0PxuORPutzmRne9emw9dlLm2aORez8V9xJEzKGV2CcZFOPj7iWYHPZXFwjplYnIEqC7ZbK
tx/+fjSpQsaJLlqatZayYFv4zi1WL2n/gXYZxX3R9TAh1dbTjcXsCyF3ZZ7INKNvAIbDq73Mof8+
wbsF2Oi6An9vQcVy14lABPTCjLw1hI9+pvKBOD5v0+57C9H5/JEco1QL2j2EUjrIoW4rYjtgt9Ws
5iFUrmoSWID3Wso+qT/pebTK1V3LOCKDKLbmOOpXucY1LqdgAdS/KPZx0azAO2oICYB/OiSPXZgf
oSKYZ/8dXBbbzqylsdBq3ukcD/cxys5zyLIhrvtOKUTX0aHgnwexv7GCRdDNKkT0ZMid/NJZxqZ+
7fKOwkp0bf5nBhEHxXyujhehd0V0GYGXjiw3SJ/ZhQiZeGQkpMl9p/tDeOUFIU+X5Kam1lncIsL/
zdy7Afh/hD4K1MKtj/p2lKD2Ub7aK/rfXGTpbS/6O9UMMdtd0O/ejL/mFrLqrm1bneFobGduD9fP
yeh5UHN429fLWZuyuf+h9Wqkid7Zg1NXJ7PSHV/9pPr3mQ4eG3iOXwnlSBpL2uBrQRadvjz301uL
O+5At7cs0E39DcZOIocIDexmJJCrruDmlHHjAw5sS+b/JqBGlU+PHR8ADqGEaP9Lo6xFuwpSHE4e
qCP+VuvJwv1LrUdnD27b/bKOXNOct9DrQdhysnTrGoCbc/4jTIj6pyGbHSgnNJUd8kxhc02pg9Ff
RsUAu8ifN2fZp6z8JfCxzzc6RuvsiOGdtGh/FhUZQLV1Uxi0RT1ci2LGjJkmz5rPg6pcfL9ehCjh
mCrOXYYms+bfSvCCSctM/ffhhnwajiZCvF68TGr6UE76rl0EVgu+LMC64OAz0PiJo+w6LoCNkZAc
ULAOtT/XGs9X9oi1g1WzZgwR4GQkbc/h6fbtNXrwU9xZ6VQ99MrWRT4FqcmNkvSx7Noi0EFEweps
3HZwuhuIaYgJrB8HPjzvIBS8Ob0FMNlS9/3pFitjqiHyyGOEj0JEyryddFYWIdsyvbvBWAFXNfic
WWLRp97wRaLJHC14oWJzIlbpv/d1zZ9Plimjc41c07u7rM5GEixcmofX+dOrdwSw8bjTrvGKC0TE
r4nN9SrJco7iO11JogDbGRd/CLU6dwMPt2UMUIgA11Q0DonrLwGr9lC+VIxX5Q8nWpm2dyr6s+me
kvQr4z/2EWeSMakN+v89iME+4m5+/T8V4Z4kddHJYNIqqlJrI8jsTcmY06iRzY2FFEVVV5Uk0iCS
x4Jl31ltTxwQR/Sa9ACZTgvNuwOlWR0f9mfYjaPQ9PJldf4Ea+f4EwUCyCKN/25Xi7zBHBtYrKVW
qEaSxAarUbmX0xM56gAgWKAxNp5Bd4uWej1rSFUirnjj0sKWqHhO0BFyFpvlETIZl7PjKQ/Q8rLf
UFjtpxTSe3qDg+iM75rjhZuvuGgoUQypHrF+Rqn9qEjXQBofKIIec8fU9zD+TVLX0V0eWIOJwPvl
LpWesYNkIl/aHxdWnnYrn2Iknsev6cES7UPFK2et5RelIwkYPyPtA9LyKx1CXGMfxK2g0L/LLvJe
7nCjjZRZwzdeSIRkYlK1VglyvG3NLx6wkWIJPAfjT2xFRYTKVH2A3zf0QbAB5ukNikJ6/3XqCtrk
hiAYPrs49hkSmFrJCvLmIrzD2WrziraSU5Uqz58bMaPbkQCt0EWpTpDQ6m7pWN8O+R2IkjBXjeXS
ds3BOFmW9QvtUClCghU+Zck5E0AzM7iNE5SCNvp7C9XsWYgwxxg6ZXgIk9oqVK7nUBDuE1FHC6H0
n9N3QdF1/Hl63pBgV0fNgkIY75j0BjUBO8T5NNOflSbHBfTpYqoXIC8dIyYmDsd5JHId2d8AbPwr
HqAmTxSUZvbNxE23Nfp/ue/wdu9PMxNAYF/lvtAtTE5rsYbIggzqUJntq0aU4vwFpVjm33D2pOvc
+ZKOoWq2OIOJUOcxU9smNUre5f0Olf4TCoq8WAhmZcSQzzA+OTKm3OrunWGmPJ5irb1JPfTfSUbt
d/T7lNHbXQLXG7JBjaSjoZ96+HkREnvHTrwoPIGG0wgGRrSH3x0yGc0TWXtxJ1b8y7kOAYoRNh81
Kq/i402T1Z2ThxgAAzt6F/g1fw+gOZqDtAzE2ggtC8egkYZd0Zsq2KrMr1/KWwtNdx9/nxwynsCq
h9Cxg9dgB3NpgyYPexZ/1Rr9zC1JRwELg7ZDFnazb/FT7sGy1OLye7bH9vL92mhHFtZinsqYTny6
IxieCEB4N5eCpFA5KDWdDMcWBbevyvuzL1QUOhUynXlEJgyl3+Jks9Jc1qlWnzRb55RJHvfk9lM8
hwwbFhvHmGxcuToWkt8DKG46vmJhWVUpjTYcv4Lg074AtIBdjxQAowFU5EV6cU2lLMziLFcqbY5/
Z2ZpSP3qJFMDWx9gnuPbBVvrNxBbVIFkpPfu3Yfcsh3aiuF5uq6WFV8P1tje0TAbrIPTKBA9X+lT
BK1bboRzasOjQCz+RO7+sCf/cNtX1yqIh3d3fIrgmrX2qYJTpraD+wYzTTRmrfh8TX82ZMlamcxu
keD7q1xop1hZZNQ2XPkil3qQYGjllE9L2nS4fHVSxHsqerfrRqvnayWPnItvG5dcoKduW1Q4FjRk
Kdr6/xua8veys3idfVFVxeG+zoJua9RE/CI661twMozOKzSHnlXXmiOyZP3fUeLolABGjBPKzRWg
VD6jJbjplwghy3sgJ6dB73TLcyCfPoczdNZ6aA5rHI1VXw3ItX8iZyoY8RbTrKAkvoK0Yep1v1QF
sLij+OP3KDsOoYUMMizJEye0JZrVJzFUoi8mfCZv2v537+IW175ccE8+N72kGxq0ANS+uc2EmTT4
07RoynTJo1UnEE+UoOCze/cyhXYM7rV/zbvR4VNm14UFudli9/2fNi8MeXIUPdaLqeGckFKL/9wN
XvuesplhXruLzhVgqkcLfM8ZgKuXDrMXAuZmkbyoWHeywie2Pv/XC2vxwWjcUK4Dy7pfcnziAdaT
RyMv9MYtu3+yo3quZIxL7TM0ZKNX/nK6NW4njS5p9m11zAxG+UFeyvtaJRFuT8yjA+qyVR9YYhZD
OW5eFtUn3uWLrIoPpi+h+RZpTMUKYen9VeyUC7zKNPkOzOF/ZnxGbcfEZGvqGI9o843qIg/sG6kR
jtrGPsI4tQB19mlEKUywoR5o82TaYM1fTPY/sO9zksPgV86aeiEI7v1IZC1D1Ez4wRNte227ehI3
OnxdmOlslZo4SetQWpvTQWjGDTWgjMG98RzXbZKAaww5oA7wCSKNYSqhpzjq+wxCQLsd/mBZrt0S
WjJlrRTDRQ34IZikMNv3KqVKD6uTWnK+sGbakS4onRMTcoGtU5PSsj1IGl2vqWenCFxe02eS7fL0
CP2XzKnxSG2z6I3gMKHnwuvaG/JfKzCxz/GGs6Ae28SQ1SJEscQCjbIPF0zccP+AL1bSbUBpk+08
z1qFRIwKWLGmaOLfQT9w1cJ1UpbgkymoDmvenrWqwOjX+h4gb8LHrvdStt+mgGzF6m6ts3Y2sa5p
v3VUuh05Pno3/pE/d5/yHg7wY9PYlG/9rfZVefqlZsqaRLZqKO9OPFNDXT7egqPfp8/VtGRPuyYl
Ztg6HsgyUVZm2khxokiO+Q+sCtFkBwHge/hGaEawvGP8iAWSjZcKDB4ktJn8B5LlQy6aZNSbvS0x
nxTamM13I+pGAJgNVk4i0LLQ6M+PfHi6E7nbrdkA0cQj3GBj/VWkUC9/CGsQwo+hM/Ssy7yHGTXm
9g2IqNzI1KKgzXbVnsXzM5SXy+voDWV/UbEii9qia0yrImfQwU/dg5Nn8Z5pDWZafM38dtf8P0n1
kV4yN+AdVGtTSGxQzsOUwpOIkiPqwmMBK/ssWLHQ6EaD83dih+zXw2RF5Pu5RTtF3F1OoF3qnGKS
o6ouBCuWx5zFDK84DkQlGGyDLR/XQdkhrtuDUzZkMQ0OiceJYuJlsWffqeIK+CoQXUa+Q+FhTJVc
AcrzCGbo7LpjgrUYWbRbhD+CuLIu/7K+yYaQoEaRlkgCkYMFiFgyTOnew6pIL7OBheAKdE2RdUJL
SrblxmAiHZQxorK2NEarCKZKKGNiAllnEasdQScK1NRf7RwVjPaKmz4pGBm1v3ey/NPlCcA0RlKH
FpreOuxhSJTgcQ/4Jcy+Tzsxx81+fxiym99/VRZd4NH+EaxZczUXqPVHa61FSXBQk0N0F8bXsF3F
K/CaAGHRAy0IBisnivOS9/CZ2BRBmUogKjn/29NRW4WSzZDBaUJG76rlDBEoE1+UcF89pwKLDmZe
OQkYdam1e6iwq5ztACQYlTNTsjbmQJzkO6srF35fn+BlVVutq5V36JW9CkoY0fe5sfF7jOOgzijI
FiGTfAFYkqdc1vO/valjLgWthHhQwU/lHakOyv1pICvW4eb+Wy3VSWK0X9C2fduJvYv+4CiWJS8p
UK0TL4uIZz9udVQvBPPh8IZTqZ3AF6Vjrt5BNtqFkKXAfO3lDYfdD6SUOpTASzBy8lq2O9Lv3wXi
JgOG9Oz31mi1vXsYI52GxSUfcd1PLpvP13VHYsdDK411fzNVtpZbiqrivXVCX6UC/DoYilCN1dO/
+QgEgWgKrjoeeH6PaTFf3KlYHAT/UGDF09tF83S1qWv7ft0fAlds52XRdt+K9urrMTizt0HDoiQw
BMArkNv7vCinPnucKC0BbPtlxvT/crF/wgXynXceNV1E49ZoRApXzjfJ32zbYc9UYhBYpjfiL/k8
+CfzbyqrQrnxe9YH6AJP88HvZVLJT9zkS3vzMB4YU335lDWKF9Yr40WOqT1uqX8Ju7vbIpjj85A5
qlcC0b83wSJCUpWtp4R9pmNMnTefeVqvwy57tw+2OyqeX6FuFurS8PuVRrZVh90k7EkuLFJbcsXd
Ap7wp4vJ6QNioO7J3Clju6vD3fP21S2zyk27CW/3o+jeawchv9mgyafAZZWFmRVJVn4Z8zcwF9mS
tGfO0i/D+IQS55+uknqjf0H8jE5vLaq8KllEWt4RbBatx0hWBn9fxMqFT3D8ACe/NabfAMur8K67
gWlWlD57MRUg9FeDijefjlPsRPANgXHzfNrF0pMAFeTEzcMEcc2jxLv4f29ma1hgSLGdhwpIN6LD
DJ1PXRWsftC5tqNtb8ck7kZpxRmRKW4omyQ5qyMZsn7C67yisgoo4mrvM5IOaZNZ09u2lC0w/+F4
GaoA0shgcd/twfXi+ltc1Nh9spBquSMqCbHa7+zzUhJyxWBnLpHZ4ZCvk4K1hDXnvRxDNTaIUvn0
7QEKYaII6WSimLob0cysjUP+vX3f3R+vPKgN//ah1AOEMXIwQ38nroBxMirbhdywqt2Rvpjs/qY9
l4N+eiRFKZPs+6V63M/utCwESQqaLJP+oKrD9ym23JQ5Qy6LV4lN20ujpURgByt8G2xflbb+xeRN
7FXXJmhmKwFhgCQ6iCWGmNiNrZbbLKFczczt4Rpgmf2ok2OmICVARJdgf9Ju782Z5IToE1D1VpXk
Gez8vNLlF/acmUHBhit0SV4UWakvUQP+GLYI6G5uLNhFiqNc9BexqFmDxco9cFdwulmyXqnc9PfR
9suRBjdLjU1zk2hirSOzhgBAXDnBt4FsX5vyxcoS5YaflnL5hhl0boMtS5HM0d9lOICLFLlVygcz
MHhBoKBXyazs6ea7z+PuYKEEFUUoFHainHdWXjRSTDM5lE78AAxSind4QyHucJkpNGJ/sjRPFRaz
dc3pOqpSD5rQONtGcUoo08tbD6dUcG4BJehKa+g3Yg3QTLzhw3/qLKBkk8rEYFvNq4StMX9CURcN
hr22sSACDh/b0q29wuA+3as/4aU6v2zwBRfm+HpZBcxsAoQmuCytlrPGkH+dotPmaAhHRcmz3R7u
f6KnsFrcBRX3cz32H/EOr0rU308HdJwzK4UmC25xMwGD5AFr/vWDwcXn2DqqSTvci9TEqRxj2aY+
r6AJuyECN49C/NUYqlK2StVcHdT+/QAYdnAxOjgP2xbsfUZmL2i24md8yzAFvrIMFKrJeHrYswzQ
NSA7HKHr60Y42H9Jsz9jvIK8S96rIVNdhl1RlO3pjGHyz5dvrD2DitYLBj6x9oHh6rReIuMCvwsF
wWhx99yzRT42uMcfdskPxE6fjXXmYahVsmO9U2qBRzc675giBFrNIicw2/+4L0B6/xpxizJvId6W
whulEklHIDcdsAK66mDP+TVJUS2SbEp6p+6Pc7re3N3JnElI9Svnjl11I8ujA0eOyTtioPXZS+b8
ksre5YdKQJ/d6mzw4Ck/F/0OlmYP9JZ299e8Omo7IAV45eh/RPZJiR+eDqFLKLffU01MxiluK/FJ
wWNDF016aYsYvnim5MfUINX9bXHuf4divRt9dGMZad5UrGBxk+CVOv5ye2snTUbDNGNnW4tgLTgC
LYh55Sd+IwrKa6i4df8522FjRaXLmzk3+r7I0vS4DgRWkRVXJyosr4pZojJEgrYRNV3bAWTwb5Eq
lIokMaCbbNEzifJF7g+MKCuBYV34+5aDs7PL3TJBqKIuLwIDhX3z//rkZZ7D5LF+gJUFkl3VY4F5
R27vVUolhKG2lFTqY8CgYUpYGCbA5409BaO3ideXW9b8dHNdaTS1KNxsDXYNQ5YRvgWXMH8Zlvmc
cavjbZNy0oJdpFgamOQmsvudQIvXCuBi054Cxt8vguM4HYydpQfrj2QYYvSantb7Qfoeyn0LL9zY
C9JNnp6KvltXPn5dBP+5WUYZnhSVZhrwI3d47dmxmVIiZavMN4pn6iQvWUyVVrZOMHZc9HFmMqGE
B8w5wai5oE1LpPV+8WhAznDVAl/EEHlq2SoE+Tkbs7sC4sd+TOXWSTLGybpN4kQG6aBoFg9N0WeT
emxI/uemxYm9nrB6+yC+m1LDgMPYkJdcxO/7HMt1I5XpIfECTUR+B0mFUQsKfUnOHghTosXjgnFK
RSaKc0fAlRDRbzrdD4yFricnqtW4g7ujj/GVkElme02RZ1jm5ri99t4XgrPDQh7wH2NjuOr/nEFG
GeFjgYKKT3Jip4yUJJJlkNi6MfX5SlYJpNgBXqSNDQBPKSjR5s8at9A0jRc510gkNyWHoepgMYnb
sBhvifqyI14JEvq8piRhNzLxG72cF1nE1uZ+/v+7mw9/rrLoKvF2khlW3RRlRGEPlIWeH+4FcxSD
1LXfk5lLQIOMrLMH5zOGzbkcJ2vq3sWWouZ7dmWw2jEFsFv8NR+Mnj0swS/r56lgiDnY0QtBWdec
yeiSIcbW6MEWS7GpQWDuF2UQPGKeusVFrDGAeoVrTwDGpr+nTKyNvmz6IDMMBzRPIKYT7dH+s8pn
MMa6as7LqOVK34xzAFggMnvUhaVzfNncNJt8u/9IOrnX+a+CahuK+ie9VAVifWmJNOUkQFkFOOEh
QRzKFxWnBCr+PwaKVeYQXOk9Vm7y6lNqV2CLf8+hhifyqS6L+iwhbgQECnCON0m1esBkCNbC36Df
AKTvAQGdi2VwTOdt/I/07Jg63xLBEzpiLZi49Ug1gFa94yZ2ohnkPPgSdjr8CLU0UDETeloZkCGU
hCjtyJvoROSXeWOn1ZR8HqhjcsAk2CxzEbuvqc8NkDfJecy+U9DRRoLhniBOocbqyaH4KBh19PD2
kxBzPDwqiciig2o0APfQ+ZlbCPYlx0KQ/nf23lllufNbnHwtNVUu2W9uA4XtXhDLjRpSnbHwaIWW
QSDoDM6vFRo04/ylcpTcQVX8u4NDZsxOzTHbO1EOI3X3190l0m0l2QpIUonhUJgzUhFw8BrPbIva
ILZCP5sNC7zG7rbDhJCQp0gpPOUWSpqK1xP2c97DkqoXhYV2ovqhkpjvqu3MY6njBG2fxyKVeR0q
QzDnQD81o4KtR/KeFwjS334Lzcls+UmBxyT+WBkBEljlK1LqZwGA0tGPL81jc0ini7DLCCf/UuXp
Rztqskv/KSvE7ZYHNC59k4MM5YJZVgKqVIgQw0rBxUrrbOdsDt2NI7nz5RaSJBl1zVg8Bxx0CWZg
fruzocROgz56p+jxOdJx9amhCHBs6non/ef8/7E061zSIqYzlkS+06AnBAof0qEqPWJFc68l/drz
Mv1mdroxHHZipfTHFn3Dk4pKMlpR2dokqSGTqEdhjwqPaFjJ3sUVY1vqKVrfs28RfUquAvDxqFPy
9DoXgXM+mIg2KnvfhODxl7tuadao6KuJ93KUPOVm/VBmdeEkee8dASUoQs2klvRHGevIu2EVkgGe
KUk4mnCHYNoj+GgWHHzfbYFGtDMqh2WxOsCR9foOnv/xPuEoleeBKlrQYfPB8/WlT8RVUU+SlnZq
nO08ppv4Ls48HVvZcHg2j3XMLiPzdRSdxpz3qmHrStU7ou5QatqnuvKBCiZuLLNwET0fNMRoSbgR
5zt/KIGINXDK4B11XUpc34Bu1oqV73h2RSg0Kt3ydxIdQeLmFNeUFSwPFeQepuq5IMZ2Hvbw4vA9
qMLTKE3iYcR8Nk8BSYRYgWhzwkWxwYjoEh4bQY/dmVR3eWJBCQQHIr2UhHdU7TWZD6AcANvxH7Td
NKtX2Ii7KvOhyUtDU6/oCXTU4buHSiM+x9VftqAfXfbxYmSv0WdIBZe55VgQK6m4nhgYJA2tZOAt
9w1T9lN0sMnzsN7VFr5g9tSsJJ4Tyn1dV/Lhf4T77mv2dtzrX/2MQptjP0MtDBrszwGgrBWNaZ4J
by++pPq6waaFouVqiPMHAV1IEkEdw1knd4LA+yN51zNX77188omDnaKAeCI38P928LSsyNYo08aM
VW/GimN2aI3Olhn4HRhKczCM8dTFrKvIUBsf++OsXcmE+udidKAzT0czETVWlXIwMmBDP+tdqHro
KX/d1SQNNjQdDb2DNvs9l/eCInmmN0WxQgu3JyLqT5g/bef12VuVa7wzXX/DZtCfhYPP+zMnEz5c
8JVUWwOHE/e8klGskoiUsiMtN54BV9Q+7qVD0r49JmrtAb6I6SSsgM0ZMzrLipQ2Qqed4rSL3VpQ
fD11Sp72xq0wHQ5xARMLz2Ji1la9qysXuXPM/XcPJaeatyLvQhQf28kUivfRlo30u5EZOp0FJhhP
O/yKw+1n6rQhXnixtwFmePpuznpacMTUymUXJXk3yQsUwha9A2/1CE+qc0VMU5OZ9IeARHeEIsfz
XEefQfmQaVyVb8H9XNYsy73m6MA18dKLYLcgffPq10PeGZydwt+HWHA5+W3rD5M9lqUMJLGXF9Op
0sqy9SrYl6Sn/Hw7Cr/bN4oo0F2HXUZbGkfgmvgRv3gwbxTDXAUVVekUF2yflAgV5TXQhj3AMLNb
3q/e6+2yQ2MPIYO1/QzanBSu8GML4wZjtrbyJlKFj4UT/IZ0tTrSgZ/0V33/em8//FiNpukMu5qH
XGIPEnBHNm2lzGKfubd4y4YdSbiOfjSYKuRBMmNLNyom3tktP/zY0N7mKZyNfCx2r1Tf6xRYWVvu
hKHyyRdsLm+Qfy6QkoG1OCIKeTsygAsQ9B5UANwajnhidHGaadcJa9IPuBuCAN0TxLuxhDaYDVn8
zB3PRwpuWrQMKxDZyT/1idg82iUJTggnip1vzjFoaf1Ml2N0iiZHkFHSbEP+4cceD7/LECl0gRHt
0oxhqs97LlWIwJfKZwGPixEYc91kiRmN5h5wiZmtcyprqN+MXdPh5R35kd3bxnY9gxzQQ1OB4fHH
NavtKcVmpy6ElQ/sgYrV/gtL80iAmtLeCK0tG4gRCPRAyyY5MAD2voaKv71iUZsMdaHoPRhQHsfD
XgWD0KNnJFlO0xcQcOZoHKltP87oTzZAcG6ZtXqA9SidSVseW6O5H1zRlZSjqjSqNS+OVTlJNU6A
0vWkj6HypVHGYDXwFrBXKv+nbzDayDLi7tXFIRwpWM5WAsHAvkwRsOpY4yZVfNLEer09aLURTlZc
7Ao0aBsf6dhNfBsODPwM7DhJuEEyn/U1ErXeo02l9FG95AoCSfnX5fXAs5/wUQodXFFSVyb2kh/m
Zf4zre9s5MeXLpTlV4Xtxi0SOSKojVh2FgwcgrQ/BrP+7xaBT2U0e2RRMGgLsgmwCulC91dQo650
TlcSr/aILoBYXUwJZxaKRPGrFQpRi1DtkKGpfi54Wh11TC6mUvvG2s8+r4noL3oanYHKYDvqgRYK
LS/y8sHTi4HIZMDW+16C5OX9gGq39Z7kB3qhkRbbLZLI6QnT0TiverisEqru7VZC8m1fY0vVfo/h
/neTIzqLyA9onW4j5QQu7YgFDUG+lJ1bsjBddM6CEYGTEX/9fo0kbQ6oecm1gotYUB0+fz9Wygj5
T/sz4MSjH6lpQVb7/33xBqL0BOLXSmQ3ooYknYH8TKBJk9uTSX0u4xsWiRgcpSPRSvR/7uQsvfBT
ZMmcM8tLxiuVj80ZdR0g6UGLRPAd0BOKUC09jEkAlLyt/P/p9WFdzXFxGde28Qc+Euo7tm2Q0CdN
/8/Q7lds9uDhaV01114hMK+BIdNGA/Zhp/QiaRE2F6T7SsdAHxFo3po62u1L2OgTBeV2P0s7OG4t
G/GY5XI27IBGwB5WtR4f7Za2cvy26prNKVB49Wd6sRYLIgkJDwqPraLYiD4/YX7oXEv9nv26YV2f
unnquIUu68nMU7KZkwmPtllB2a9RU9fNA7lFrmyUm5ZmeF97MlmXPPgkaYext6ef5UyrbYZQK0Ck
wocITq5NX7/TP8v+AZNk0auQE/+DS6c3Z9q0+X5RSY96MK0PnCYXispdLcOEW6xpeCYbyy/u4w9g
0NBzHOw6klEdihoPnDsMC+GleT4UfWnys4ce68E0fhm+W+J9PJ4Mwled+lqwiavPfNYVY9lI4h/n
vsPSFM3NPZnwYoz1403wfd2W4ey2R5Eq1l+FtANx/f1RNmKR3rwCodsCH/Ez/MJNsARjdeeFdAa7
PmcYEWjoPa8zO5HUju/d+uxfbHPRbHF8cfVUuYM5J1hLIokKErYOZXD5uZtBA+tfY9tGu8fVP1ic
pVIOvRejUaH8CwK/bn0QNiDLiZ2ftRW8Fo4kKNBAptp1eFLFW4vEcgDILOsta0BeLL+yC6sIpmwz
REfZrOyJ0ptys2gxtFStI7gWWBHRsBZn6qbcPO731GQAf3gkYZUSa/yA/PxyC7QKItRSV3y/DB18
iJEeenXiqABosXLxtPw/tzSwlvdrDn4WuXcKXAZyqpVxj1xV02jJUPkMLY5fGJ6c/rci88tylt67
L3vlkfqI115hZ+t6SQ/8WFGBMJwtOYgaBnGU6knU6Su6Jub2AF/orWATheSKHRZAfFzcOB70tqUw
2hu/hAecJbDOF/BeRoV3NhhK0A3qHgs3lTmufvy9jD5sFwp5rWBBnU8dP8JOntjEGmo377kVzfKV
bsT6p9hqVBnxuVXw56vp0ziV0rVa8c47MSU/akp4OK62OKNgPZkOF0U2jLqbrd9LNMRxkIiK4O8/
JPh6YxU3+TWnOYYpr/KV8M4e3MarTZCaiJ9RK7z8e2vzSr0N4WTRhv8pnDYy1JbX0WkSrc2kXqGI
32Rvw/G0KqCuyhcvqo8v0lgu/kVYqZeFJp74QhNKhadHDHkdA0DYIlXNLj/6TCZTdkzbnwKK4S5Z
hnwGnFCDDhDd3KPSmA/dR3dMm+U0yLjDyn51uaB5u6gDuIuDf8Q42dGJB1ArGUtElE1AKCDmfe/P
/EDFQ/ZBO7LuMp0clngB58S71PnnksBPd0Ygy9ktBFByS4O6qH+ieX9dHjz2ymbwrxe9LrEK/lJt
f5IsQhum8a7vPem/EroFN5qjog00yTaKW1oMbzOlaf3eg/Axi/6BNm9P3E5rWKRUDAuckVVuDHUx
uRq8CpTLKbGG91EHVXQfiihf4uScpEAbxVG4fSGr8x5w6jJuJvoawUuyfWPhBWCHJNY6JHRKekz/
/I9hOe+6louKbmR+mjDo8nwUbTe9+qv1//sRKuvKHaCpxUFI85xx4RkUQvA4x6M+Q7oPIXsvb+xR
10PorbK4QtVVu/20Q38joNuSdgJywyZrlz2Y+gfo98D0Iztt033POg+GB5pxx9xbO5N4At4+xHnx
bzTyUNowO2VDsUXerZHLRqcg0N0u82zKvxhhrT5o3wYQDhHFhBJqHhWw/qyOr4mI7OA7ARmMfU7O
UQr/pwRFoDM2VzT8hCFQ/AlDlUZyezA9frJMOqEnGC9zn/Mi8juibY2BH05f4BUFWL16/QHR9iLo
NvKXOfWaPeCL1l3trReUGjgreUmOtXxnPvHi+q8Q5KiVUoGe1cO/n1z822CoYELBSDNFoXqIFWAc
nPLshC4wIKdlVnF63VgkClJInGv8KYJaiYK2HODHMDmnU3HbZO4gQ/EDByc55eXJRE43aaYXoOdh
a2Fm7L+Q2IcdmQRdW8Vceqh6z+B9iGfkIJSWXyYDij0xanbhcSZ4RoNY7/xgVAhusvjpcwoxBH8X
QPwRWQEYQTXWQfGR2OAXMYMhFGRN3/YUmH5X3P7uryfxATvImnnSG6NcCOrBSPeg28GcSbbslIBK
HrwyA4oVQcawgP9RvFT0DivqXxbXbetywAvE/s1Ft/Uv5UwHCvuwbugVHkaxTgR+QAqr2O3EL128
v4s8ua5c0T/EqMg3J7o8ctP+Dkc8j90Pf1rC85aX+CcM/65vRdi+Qx5rFEJl2rn199R3qrYDJa/v
2A+2InQFBQKSZPlOT6PdA5c5bH/Tr3tXLoJTj/U1UspzuyfX1AiK8nV2PtXj6U4WJOooYgnxPwQL
MM11a1G1wQePe8k0cPaBRUe1MudjAcUeembG6Cx+mLoswGXwZJxNnJ8x66DxYGkp8Ne4ZcFQYdzG
mU9mVe5ofCfW3f4loxaDtL5UTGzQYAIaC42szofa6Mn+Ir1hvYhqrgy5lVEkiIdsh6XNhV/Aq85p
vR7cGQeTZCY6sYGMqbLQYr46nPGvy2KWBEgv51I643Oj87xK567ryw7GKiTqqlwZS/jcVtunx21M
x5wVrKZkB6beysyH7drwaR+6VXePjLZqLv3tNPo4qyd32Fpb/apPbAl+m95rP8VL8ycZgsNny9QF
SdC27DTc7ZIycpF3fZihKP5b4LY71u4M8hYXdl/853C45uzxOYxNJN9lU52W8D+wwlNo3cY8NKFg
PYUwsuZhDhnJj95xWKacc/sgEizyZSMyJcOJebEXhP0RUGJMEpdyBY85x6HrSbrZeKD/0kq6vkS2
xxZJRx0Wyo7dunlOsnCNl3ZShZKQ9pUiheHYlmwAK36PgMavY7/Ax2xK1N1+kLybB4NKGQGonz7N
RIXuLflvEl7xgDjcZAo548i3ny3x0nHawVevtLrbIBo+EgqWu4MqoAqiEB/feMEZgT34voabSuye
t6I5cElhhXLJ4KSvg7IyOzctln7xZRV2hwV0r/da0HCr9L9Cuq74SPPALyO7Geq9fb4l8qvVsfFw
SPPBtngfgo45rnfnXgnno89uoktjau0g2mV9NfijyIbCmymGN0lSxYbModxc3ZSLz3Ix7W0xk6+A
dmDlr3yoZxGAgOzn5FiiKiAaj28Itov1yN2rL76d/bPr3E6WM5jIhWP3H5KYYQCEX50PP59ZllFv
VL68hOeKV7Yx8kWH3akUgs7QV+N6c3OPQ86f+dbFBJfeQ80HAam6NXq+IF72cLVxPorHjMHQGCNG
gPm5gUYnFjcWJ0Lgx0nH/b8ku1qNJPB0erqrYDfAb3DABhEBhMkrYJ5lFKv99cFgoWIl28u4UEa8
BVMmqFOmmjNiVWmoGwJncD3MSglodAm/qx1YEYHk/UN+mpB/3RDUsM9hsM2AGrMX4ZM1Fe7Ls5By
a/qgbxEEIQvhqccTMCShz2jLomM4AGng3mgpBIX34NLfOOpDHOuLZVoP6NbF6lJYxS5qjTXgz934
mhHtBepYbOBSizPnsjJa6jL+tkEY7tV0OwtEGSLfJ5FzD8U3AxjAnvjA9UxTObdHWsOHi1NgmC1D
cxmjMunemskX43CYAxkqH4Y1V7DyxGAVhAy101XJhwHHrR2hpB6pKY7Vl5bWWtZxz9GjAqTS3XJJ
3qoIIBsPq2oLP2UwiitvTKe659D+cX5L9BiANFk3plYweV505pI6/x+VHjHj7lqVsQy5T7KC0DiA
9QIdjQmO4BK8RDpenQF6oWfAsYLoygt5pCKTiGHxc0etpFj3jOaWt+cptsyS/XtLm7cN7L1HJvR4
wBnmVqLGUwwLl6506mTEuncL9iFhacNRDNXa7QT1ulMmkW32BaKNsV8FVBKbcpG12vEcPd4Qr+9b
OLtDrC9hRt7+Wv9DEahU/piosbvhegLXYn1DrrnQlPG8s05vuYfj/xNN+3x/fDW3YvDPURDqMaPW
4d6Xv6xKlzLxbcHKAQsg8jQ5bBmXyByCt4IQrrFjtP5gF0inzv+U4BHw4ScEojtpdBR35bC4hDX6
JLgVJwkghsjiQ+pRPBSo8iodMwiTvb3ceZJtbmLKALzCvlGFiI4UU+m6XbB6NP8VGixS5UIIklpA
mXwop2V3VBXLYGcLVMwSLisoaKXZwJKyuJKVH9eBZAqsQS+hXWpFoKC6ElSwH3egjYOhbuMoZULl
bKHzsmdpdQrt7xAPOoER8KXXEcCYoAuMxcXYECZl0rFoLwzYumcF/oZ2Ap0B7EdbfewH7bvTbCRe
Gvs6vpuus7g5g4YbsdzqGUlYRSA5KCMSrGJPImpk5BFnw2I1GnskZjKi/SM3mNIMqy88Q7jrMnzj
2F86nKmj8qF0mItM6Figd1XnSjzqJc1AHfgIXp7ZvFdM0lVTc+HhhHMPbwchO4nX7ZDtSE6IxJ6n
BpiNSyvABbuAZhlSvP3eQNl0yO1OZ8cZM4v23RpIgsSQNGIrEokImuVcHgjWyZBkDa9OmMmOGhiX
WLubSALZW8nHwHidfDPuB5htq3jpTmYJUUOL8LAwRqCmpo0VJC3NX+kaFi3dL2nCQ1dJeDMijy3J
Z5wm19vmxNMYvDuKTtRhoH6WXz0v7tiVj5uFlLflgJsLJvEmwxj9oaJaUk0XnSlQQzxROkZ6f/Lq
GceLES2II2VROH9qAGkrD9Ai/OYrgHQaNoDnxb4wP2vajys9r/qNT/hGjE95u4/V0uYeVotYL1zF
L24nhNCsxIZvyYRTyp7vlkPxHNuZkXFLuqklrdC2/hVyY66k5Ql1xSenhUdyRN9B2TUEtPMDxKWc
CbeuSganrAyGPqhe8XesVZFgVdJPoo2va3+QHgzBGp57u228NmD1sNQNWPec4+EmeIPPVrstbqB8
UsYeH8rQR+1QiIYcKubCwdiIeTCjtCtx06wH3H9b3sM26IIYmzRwOr/lhQbAwKEMsP+q9lJYnQHH
1WeHz/+3zu8+2xuk1iA3dTU51QlRi3aN+QPgp9ehpsk+qfy86vBbYirZ0ZenOAxrkXFT23qsW6sz
fJil8LLGiUIsYKTb94Bcpk1XCaacqUph2oxUqVXzTiBW15+UVCLpxAa/sSxOzYAQcMroVNCwveH3
cvKfQntSbXW01AQ1Nhwc+1+kcllqfnej6UpE0vLxT5MAHbNaJR2mojKxRZObjOPoPFDIgCD0eB0x
c+hrfqFuRTzBRexvSNOEFx2FIUi211peWukekqaQ417PUenz67J0RswL7exRJ0B5Ob3Zwk/yZeZ8
HvSTBiMPEygf8KRcctpaWqU5SLKo8guU0uY80OmmXK4g9jVbmyi74JQOC40jKmm/1r5WNEM5FAJS
b7B0PF3q4Q6g25lO7Q1BEJj2bDsCihQC/cULD5PWsECWQm/B2jgWY8P8CBDTd1kX/kO0KVs5j8Vb
A7E+/0TzJu6WsgLDdqq1gjzCFH6MT6V857ic5So35+IscIjY6C4j+V/XjlSgnIM1349MZyh8Mdvl
QkcWHjmx5Lx7jUhypvNTm24WjMKG+LtUtDhaCfq3+N/v+PsU9rpLMbeA7ORGSVcRhC4OegNLgxL3
A5047aBht/L/6p5xABDNBN5XYTgvX88mIqzrBQyUBcp7euw/RZD+P3PHakuUBFiWEj2BZ8Iifrz3
la4olA4btYTOOWBgxkkJNIlgWV9E4oHvRV/JXoks0Ms2OQd0cmAyOhMk3PZuoaoP7HUEGL3dT3A7
FdrsGMKBynFZGd9ob6i5ENv8V4o0vl/Pi+kwKVxkqNSlJIsY63HnrMGWUyi4amZ5CIvWGxqfAij9
2cYV9Vcm9pnpLiRiKa+6HoN02on5vnVCJchWcFw6k+bmUnq9ZIuPINGUsFGL9iY2FxjvITDB4DXa
4s3OANtOYvki58xdSGIg/S1VY1g6l8m69djc4+20GzG4g/u1OrzzM+xrE/tGk/CpBNyKuPTn0GTa
UpMtGSyAw6wRxUQ6gpOY9ogbpvnfK40fhJm+45n5j5+Aeh4GHzJw2iZ0sgvbmJxHU1lW/EkyXn8i
2vhEVRaYWGgWjICasfh/vo0EQoxBOIP/LH5gJ8UVsIkPSC1fJ7aKD+wv4E2iUi63Q6U7+hL/0dfP
tTkVmKUNoMvoiXcF5ZzV78ZHcS7w5f7JQWT+u9urcyGI2d2I6ZtdG4M4Io/ou0Zqjzs7himBTwoB
2QUw3qHez/kzTwTCaneWdc1k76U75nhXEPC5E3JClHx3F1S+O2wy6Te3USMfaZOik/FsHA9PUk9Y
LciK8cWZdaPXKQaMS+D456VhLij7+mIU9gv5Ulgn7jfDSPN0Xw3CLCnO1SeWnCR3T4zJyxUXyMec
ChcHE3n+O3UYa7aFvPWs01uLbykOavxdltnBZ4XGHYoCFvm8Ho0wA+tiZl+6mKtqoBl0iTRLqqx0
T4aQP5W9SDnSDrBOHaAeWZgeg1eGBKVM5wh807rq3OYNL+0NOdpQA238vBFjG0uxYDfcnGhNpitt
tRIDWCIyhix8YgRowdLdIZaTI4aoxfAUWvSJAGaqonp/mrsMMRYO+AyR+tBMFf9psm341xCXM3za
KpiMi6gr/RSaC4HNLf5KXFpxti20YMwqaer3OJq126wcy5t21DdCze2n43lQOVLIPCCweO+jSmtH
oNEyP1dd4RZk09yiWolGg9kKt/3j3RfBST4e7qwViAdyPxfZOP5wutqd2BrO0U3w8LSmNQvLmGVT
9iVFTRgOpfXsjzzWYgMrbNNIpTIbaSWgspbxsPi1SgrO4/j2OBIB0qb61gyIUVu7uIIdhppujRJX
dphi7uVilAF9g3QUWXGXE569fiWmCZoatJIpIYxpfQR4MkpInnV+4SMJg7YgEhrO5v3YDWjmO/+V
I05O1yG9HRpDDY+Xj8LQHkL8Inb4SYzKLNQSbeLOPl4meJ2Nexj8T2a9phJEkUXp3g78e4Szwhhm
A4Uz/PtIWTiOjRYqKAKFckcl0ObrVV6bZ5aENnhtoDQY8FS7DECwOuswmmI3iuLPHpDLfn8gZXRK
SecEv/mw83nIr/mdajwfsY5s1EcUM2MB2MbOvBupeYRhBF3k0P97pTjyjB9cPqPLclZyCcYU3YFm
TdCFE6GTfdI0S4hPYw1hvtfEz07qyo8Vo3AME7Kvmu2nEoUV8jChhvvJSD0tdA4f2KXt8QcRBOJe
mpI0qT99quOZor0WEQ/Tn4fz20ejsXfeyh1W3Rfe1kcuJ1dVtrggG71i1rQnIfAX1JjIBmjfw7/G
7ZHhNF10O9Pfl4+GhHBOPqKX3j9YrESkTRpOHIXiXkjTx4nupLfdvgxa/LTkg0Qw1Pq/XCUOEOjn
ranhWv0C/5asDUSTOw+1YAT3aXiMroKikkbcg1ofeEh++Zx0NyVp2CAGpuQG75yU++qobsivwgp0
MU0AztJCxBlasbWDDwRNJPsSHCWUUqsHuMdZ4LSCjUgYHSDHZsi/N1vsq91h5GbRuxJ5o/QBTzgw
Jv3Rd7Ah0e0ciFFW7bN/dqZjo5ORrFSnJBYYNTcGQM2jxS19MRIvxD6nnCXsFzPRASQRUlY5Q8wc
9F8XIEEqaSdt5BIY6CbNql92OizTLMQRtpjp9HhLPDo8AqU7wje0YGJSS2ERQ+Q21TKaTOqg+Veu
K1tiyL4iMIFuV3l+sdBKdqiNhhGKYH0jBEm3a3ieRmSeQkPh5rXB1Ui8/tcbbRdmbKwsaZKdTGXR
3CKbjJY282UblnVnPWdejDx/gnfzMpdCI+DeZx7eqAfPaJeeXNNrBOASJXh0ry4qWHZimEr0LKXq
9p9bzKZpGrCRanPFX419y8TtP6Mxxu/7CdTcR48MmBV7vYZfgD9/sgJ9bU8X6fb4FsdHtF4jQ5HQ
T1Ka0NJs1InoGzt68ktl8kjEkirUHBJuYLGYWajrYGGYd0E5hViyJDaB8eAdSu4YwXPL7GJns1M2
4jY3fyhuCh525NmABQgRdtTnRMyj4VTMArpLij5TPZzdH+i9TCruCw6ATV5iQMwA0sPxjN18vkR7
oxmd60co7MtDRcIWnCMnktV8nOcaTtg02MgZWbeiAtQmbBmbF0h+Uz1DGRTNcly2UUXKNK7eWpzG
KwUcRrboxvQ8iTLpMYZtGH/UGHQZ3oyd9yb6MxXvCdVMom9AV9mmqGdgHzkyLn1Z9FrKk3Bc7Xo3
8lnPQq0aRFxSZdMM6eLiCcDHr+I3R7K3Tn9qyYpWNA6MqafYlpZBoACggQlw2YYuDcSrZNuMb0iJ
he5/RFqFCwn4BqvJVhSKXzIkCYy+m/sZ9TVbNgiUQNX79waWzI7qm/zoAXpYdrLS13jp7cSFrYn6
ZlRpqorAbVkzEAJRf1k9R0BpUFoGezMSc4UvH6qNDQkcNVhA+Qu+f9vTUt/fr+5T3xfRVxaHrSuM
GEtJ7d2g2Z9hOw+rhpRgVzFV7y8APHhpcHS6kF6qkBxtTrKBVYFy0OEhbBJj+x6IAJdWoYhLe7V9
LYKmTTlcO/kqPQAAH7RtmIfcXrx6ahDiAJjY43v/Y2wGluf5QMbCnjKGRTsPvUQRisophTKiioO3
AFIPK3gkXkuUtgpVG3F7N6tfSUgoEFkkKbqsfBre1RNCp/DibD+69unnvll6Kskme3wFrN4pY1kN
OtzT6OGfVs+cENic1Bl4J2VWhFAkkkL4gbWHvLEL/P8oNykjvzbSu3F0mmjhA9fv8WnuFI/gUFCu
1L/W64lIqlUwlOtMGM1O/Ki1yLfP6bbT8ZuS4vtebvUHeiZgp0LaiMA8B63eaorBVAGvKIiBMgPZ
hBPRxZGQxKMCAskMa3eeB2OGfR3lcubxrIwnMMxEiBZULdICQvL9HyiEMMy5EGph3+rICq98z1uj
UeabGT0mbsy+FTQCQXYxjCBvdQljYgbzhSEH0NWuc7dZwL5DO9eFmcFrCK45FhxfgLBiZEa7Rll5
fPl7XvquM8OPsGm0tYC1qOavJVSDOW6s67z2HlqZfjF75Rz3SWUHs7QlIgzfOEUqdYZ/7E5xCamz
aFtd5a2aSjOgakSuA0mzeXFYLVrFo2xXGTQ/kdLMriTWhjJwLHUU0UHWyrlD30ZM8LWHiZ/lBV78
UVc1eyMfvJtEzIMuzYH2W9lGi7VstJC7TAXqLUQ4hHHreAN52eOy5WYKNK/kqGL2U4bWv+udjRlC
n8H/uBHUlZgnyNeJRmbFU6JD32t3FTBDHH/BQ7heEQ3G+jTX5NgTRGM94a+acoMetGYn+27Y6xD3
teQhnZvyOf6+UwEiimnq8D6S+ySyXMCJz16KSatHCbO59x9351bGh+hpCmalQd2SlIS5kWcuJuoU
QwbSFRLkQgJqTFpIU+A1A1iutfdk7UDU+deiOaEP1xy74AR0M8Mh2PSLvlHMoMGJRuTqQFs24zcG
SaiHEaV6+ZMXb20ExEYfd0iqle5U2lf/Au+xOkOGoj7+qhr2Y9yvUqliYploSGapM7i2M++VCzGe
Fxm5JlZFOSRu2qk4XPDE1rWh9vgFM0dmsLgesder4dcJSTSiNRofbNo1jhAFg1xIzbEy8HGP/iKT
OA7VdWKSliVeSD8qm9ncuALHbWRDeguOv2r2+x8596GNcL6e40joLv7cCRsyu4NedvBUx+ZPMvDw
5PAEUqh4WHfZVv5RlNRKtOZUcP1mlDdFmNGXPe3gM6adaCjqDe45L2Y96vlRPeAvlPVakMMg0U1z
DW4DhO7rhXB/627DSm9hfUUd0ne2tvJOACposrPYKs8FZgFXSKpEa66qzTx3tN6cD3nCu9RneTqD
zDMPf/Ntlko11rAlgnrFF0nKZhpQo8FdpLtvihMUqFdeS6/+BfA27eWTMQrvQ53xfk2YRJu4g14r
4eZHndoNQd67C5G453oPpCJLKqMlZSOzE/s+Uz0xNOb6pXdfwuFSJjyS27hF05DSJKSPDp4rUrEp
VqPbsctGisMWBLxpC5oQHtdYiOdPridzjLwT+TROq6FHycxYO5aqToPHXiuFShrPIsmEvXSm0ROP
0foI04wJNeU/llCDbHu0ZPOtMxpfpCFvRXW76MvUcLMl+1vpPifeMKqObLG0WTMIjDGJCA34xeYS
oNJKPvzrm7kXVCwB0MjKc9162vElXUDETuDZGM7Y+E5KsVzg7MiLn88lNKCmQqoTTg6CjSXM29Cp
kxpjNHJR3Zs7oxCnOgNyZfLpq6NZ6pPYchTkQHU0+lAWOyiuiLOL375vKpYpIF1OmUdeG5TdWlYR
GJZCl9f3MPCQb2U9KdObmFErdbORXvHZ3bvJSXD+lAwGawX/vDiLl/+SW/Upyor7ZZC06xbkUxUC
GRv0NVt4NIElynZs/vEL6hydJfp8Wx6QtrwH948ZJCItlciItUTD9HP/KrN9apEkHZVJfD5r1Yrn
7m1iVWScyDw+gysgH9jl4fDVK3pOf2bWqSaPm3r2y62SFvmlBZtNHCeX9SOxNq5bjzqAVUfKvkIL
Zu7mfK6UkmkYigbmKKvCnJW0NZsTMlzjtqCBHUGeYwtSBzZ4J/5mTar0HLQVlBE3VNdeSc38cZ11
MfN1Qr5BPa+/g8JFw5qJq7fEGvCRbRc3QqiDY1kORn1o4spRdtd6zTX4J9R6WCyYuxQt9shLbJ3a
mdpf4jA39r5NDbXpMHSIaPeP43gUtMXhpWP/jXCzkaQSNMvCPkch7di7/dbOJUDw1LIQsgx5gMLA
yZCeY8QRTWTva7KoKXIt6f3PU55KCGYYiqKvAmP6fArmNFQeuxbfawYJsQOaI7wUXXa2EnIDtQJl
YmHRCtQuf55UjJ6V4ybczzbSQLJBILGZ5iD4ZlXSQEoXVrCNuI4PYVsyO79V28W5qJ7VW1Vd5Ebq
HgPlcTFVNFzIc4gIA6tCQtE3c2a9L27s/fes1lLTUd6f/FVGTwzoSTkNql3j9AtYhgCQ/zikg0ic
JjZ6Jq9jXMYKraXtdBphHMURBy5XP59ZStIBe+u+SQzrhinG3IFjlSHIIcp7HaIo3rXa1TV/nspv
jNEGIMiFui559CoCFPx+vGXupEU9OsQNYFIST9bccZ5/rpSJyJUMwmgCZMBatchW9qliN77lGg0q
HJxTLwMfE6enWFU/WlUfjfSGGZTKURfbwaZ0ZVicwow7eDw2aNxhvEocUzYcmZGE+l+Fq0Mogajk
uP3LiK/Whl8+x4lORFdW9CwMXG/879w9jynXm6MiQ8T40jhG3049ZzGeeGCaxX6MDlgalkLaNs/2
F0x2jVDufeFHCPFkWyGn50Niz/ecGLb06quyr+6C+Ij3TYe7Ayd+zpEUZEHkN74W3X8QlJeJsrrk
UWOUPcZ21E3sEC1Iidy+d4sGzMFed0xHpjhJytDXsdZ6+lX7AKcqCsBCEDwR0JlK//nIZh8PReNl
5zhKcoYzUOnlrUEPzK8WkOnDYuGmf/p7K58utGeMP5BaVojaNT0Nx2S+4ZVQn1Z3i0h4vGyDgX/E
TZ+mQR4aOXxbguDZgXUNqGuii3EL9kDWavKxdbjnmDfxtExDRXyOcEJaW7F4T+jTwV/VSUBpP2x9
0TJvcFSjcE2fQrLfotMFJPtcg0Uoi9lmZMorOhtj/gTzF8ZhmUBn0/0jHzaa3BqkwqyZweqY75YR
1FyDX2DbR2prdfmDAEZ6gqatPayWQA2gAsnUv6cN8YlnCW99hNWhx/WiJiC7W6en0nXeS6cJ2QMc
vcd0XvcxfzUhPv5q3p4hgjk0JXr4cGuZASUnolNUSnZLYS0QCPZey2ZcFw8eqM20oxbC7cwOjcXt
QjGwH7WI2z5hYZBudCL9kTavte8ylFrzyVr8anEUAzRgdyOKQ0z+CBoDrhQGb6L+ImZ0sIFJsRNE
lHsMtBtkF6ezAn0llmeNgiy50XWqlR9m9wKwYH6mh570F0LxDU8aP01s0f5uMqoh4PPymmoGLfBJ
41GNAMvKRiInMXJtdHTFGyn1Do2aAentvvuzwQrViO4Fzb/R5LvruqJd7juUSCsgoJyXNsv7XRay
lUNQv2Vjh70unjwH8+khpB9zb9rqex96vWA9fL6c54ReLAyl6OtVoOSq1bUGeNBqMJd6JBk2NElp
qVQTN8/ECGEPsu6+I5DRFDbHozKpQtZXSClAuXJE6m8tS83bSfOsnClibowQ2dRFsb3C3n4/vZum
rApkHrPsrsMPkojL6p8aveb8Ne7cN7yb5aHBt5hugi5n4nRMWeFbr6QTRdZjllKfBff4oa6OMJH9
QcjA6KWACUu03OHkXSJYniIXz3FvWnLjoeSIVp4vqPpaash7buwOY6mN2tTvOpEj9J0eyKuIJ11d
6NY/P352dQwz3kfDBDEehyT9Dyjr4Fe/8nRJM6pkd94c4/6P29EQHaDG0lPkaMfBPwCRCu1q3rXc
bbdGPpQYIDt+ev0hwdji3ZkYxA5v875vm9vRmmXx8ULUftXaPFVsFcIR2bHh1jJCoB6XyapPBL9t
OCMrMGBJ5bYBdL6YHFtaGkDLos3d/mC96FC2Nm3jreKZN34z02/cnVwezEdvZiaVh+RYIPlYqfku
0Je3IanyjUlqWk5urHA4E+ZAx0o3AhHdX5Gh2OSM29UIU8s6csaPIAoVt00H9xCp1CqInP9HkuIK
7COE6GTb2Co7kARj3ay9STbwuh5VwlXEeq1MxgC5LbMFPAzprKKV5+WsS9a0quZ/Xibp/VGbC8LE
stPsy519SRebBWhjOjDW0Hl1U1sw6ugkcZs/VGw11RJnq4eMEuOEgHlw8JbzdTl04si5aKKYPVMd
mODTtKbk5EEog/7uZY77y4uZ+3IqgubIBIM7oKbVtNGt5OASAFgIZhxLe20/6RPelLmLbkSjHeGi
vdXAskxW+U/iVTzyi2qistWszJGTYfGKlF1sv3zF5fW8nRj3ZcWusUIFgGyljRzW6q07Kfdtz82p
FEA/PuNSHGTU/ptg0jzg6wotj8S73tAhQMf8pZPmLdINhG8N/hcrr8Xtp1sARvyjmBMtC0LFF1kE
YfSnGdijX0jGVPwHAepBcZQxBhR1VgHwtnu+7bTGi4gTVnzS+HsnZrIQd4HlXtKp5jggU8hFVSFY
0CKHUx1G/Od0V2ZeQJpM0ILViimWqFY/kIVqFEyYOv8K+pAsPzFPy8ERUvND6fnGUQ4GibUwGTYH
GmYnJcCLtFjDrEqSNoar7cnh+X+atMe8WJ61utHRcZ3MMGZYSmRK3hUzbZxACipUpf8ijORnK6qC
kCy6ZuIorAq6sTzwwdFByCqGSeMe0ou+TdE7IN228Le9OJIA7RUjOtgHltO/eTCw3FJVglfK6iTh
jJGiorrj+6YDUS3Tir2OqfllsTFndIxmT9UBVkgk5Nhmui2ICJthjD9slgg2OlTuDgdEF0ZSkhft
PKDd8KJEL6x+qIYeYvfmZThmRh61vQXjMisZkLLb5ZYpUaH8h0SeZxIWcasoOtOyVsfHwwwljYfy
8Z1ziBCFfEGstgtLDrHc6KOPUTOQ0uZwpcfTkeyUYekwXGEgGEqbC1M0MYwQiPA5PLQ2OR6s/Ax6
2TX73t2LLPBJlwI6sC3+aheWD095m4j7LxRzWCF6Zl1a6Se6W5zBC1BwKSBdCxBKMLUxtXHRERiJ
5j7bLnnarcEog+VrJFUO8i8nkAD2mJYhimfESYDxo993Gk4HKR5WStPi8K43PMU7A4ouZie9wsms
qO0RBjtmV63hCdu9fPW0MXctUbaCyhheirL+ZKM8ExLCtpnjvcKatFaP4UiJfAjFs9Bv1c0+YARt
ZMFWK/T6gdI27c0d/RnV6wZ5XcbL1OyZ3qf+c98aCAezyOKFI5j6BUYRCL8x3aLVMc4AAXGMC4AM
ISv+iGuEiFzUCv2FDAd+bEVFfWDu/w5dAoQ5Q21roI5ko1yrHims+AWLy/wM0/a5GHxwAIhpenmW
oxXj0OrA3GV43Njh5sxiRicrMOqBEaxWXzVp0tve+5X5WEqT4BiE2NGb2ZSTdKirqRcPmHWhMjU3
MfowaQVTkM4orejHpQrzCYcwlTFKVh6U78Zy/utQ9g3s5lb6vkj6Az3HdULzkKuf2PCMJLy7B6Y+
L9v+5Ct4fPmlkUkiu4JEEegfyxX33lhBnRIbSi2YuDoFPkNlNXjmMY0Cc5lnUz2Qsyg4vUCooiOr
sXsi27M2Uv37T3IDnT/0xlzs3/z3F4F4KzSdD/bFuUcITG8eYD4oDocJfzMGvhWWtmq3IEzuLmfD
qniYnqScTuGk3/wcIotMBUcfLf7aoBqEr5xm3hXSD/hAUhzFHDPQ9kVooWCJ0/MteWdnhlCfScF6
EWkodY6xVKhb7THChyxQJoeZhGLglcSCSnQV7puk77SNEl35vmeh0Ow6VzpAfq42wtXOL0iwld7s
pC3yUxcFAlKZBQSH9igMDjscmxZozpQ2inkiik3aAiOrMVleeCkP/LbZlmlrbm4gAkwjdmh7Ej8x
VIcOnQpu89H5tW5GEEM18pqSoHqtGBSaRuhcgDtGaItIgCklfipaKpiPTEyrGqKD54yXynHf/76J
zz+JX+f4YpYEUnSx3qKZKTNhGp6OTflIiPQQUIZE7xxSNQJXhuEzs6Vvji8Mqfhlq+4Lv4JDbn6q
1L8ijaknmVQ7fLpCnCM5+gQmfQtFS6aTH2OZ/avjkN9LJ8iRmFIPCo3CSQJCy6gkCMrTcr2TsbEp
vKv6HmrfUbItg0HM/caUHd4/+kQAq3oCEKPmNYubUmNEErAqrqiw03JTOJOs9LWcujuiyzBSgMVZ
C4FszszmF+tnIixUL7jyPDjigMN0wx+sPUDK/YJ7XjpoEcSyrYjbpu6EcdKWq+Li4tssEEFN6p6Z
3rNzOqvphSBp+K6imbe3ovQl9iakgHqxzXCOyKI7vWQ1lNGTPoesBzykghGFwqxYlKXhmjTmvhlO
r/va7GIhaeFYzjgwzhHBTm7S0nKkpsOHmkfHR6gjW8DlPXxJ+e0xkQTqHWZomFEYwUaBOJtKaWVe
2e38XzgMwhZjf7ZEAxvcszxaTxhC/knFh6Rl2BDobNLN+IFDgfyy5kKh1fJCHsdSKDamGWwxjH1s
KNC3i2lGpgoRgLKsWVRk+ILv+SX0gGkfEClPQuDysQALFOhUvpLzBJGo/pVYn4hAvt6VbeZCkR4C
fFJapxLwjA1UrQNcYU940A7VCmy5NSJAmdskJ85zWsgv2GCX46SZOobZnLVFYNFHDzg1nEfKjqGi
4uiEKefWvTNF0aJ41ab28QjFVsZHtqjZFhUqgk0DJgynXRwqtLZf1nYLocd+O2YjSaa383aPnaks
ace0ZTLjHkdOEp5OsWlJDBTkaXvaTVAe10biSnkjOICPaHFvLkNNNBfaNPP5khz1HSVSt9vlWyeq
Hol5uUOsqJLr2Lz4Uz+bodIcY3WCDgLHCw2lZ11bUzvTJMgP7WPL+BFx/+ZZH+XmUYuSfTU44L2O
C8eTvgll71K2OrDY5C33+foeiuvjQSzsalOW10HGNZC/cQxPqVzuuj6TUGlen7Cumglf+0qHdMtR
siAvP8cunHtmOsowURoMy2wIPrFMeLMa1hnYTwJMNoO6aKE4kMvjwLNu9FROOzVgZ3NUZzIHyFaT
t9QjM3i6n14wavkSDYx9RlAFmK53Oge4XU9tW04H58VBlzeviMkN56tYr9lIgrnUqZqGq4nucKQl
bGeQ4zmuM4snC5Mzod2UthgOF+l+mWfNmqU20Sb85u9wN8n8W1Xil5uTefhnYni9ylkzQtgQIuFw
bsnWtcmfSgKEFWgeiP0H3r3bs3KFDKKparh0gKiXKfw4JoTV5+fhIn8s/TFLhNdUYi55PX9reDvP
sgikWbDw0ymHca+Xhi9RET0AmvEHRgctGLcOnXIdzDd0bwScC/+7TfxaJU00DBiZh+8WHPpJtMB5
w03u34oLAjhVVVvdu/qSL+7X4PPONqmgKY/xiYD9PQbY08HG8yffrYkYKIrGHBAmX6XmWPwtmZyq
oXU16Rhqll4Lprl3+HyHjOmqwTdxDU1e7D1VC+y3OvcqJwfhu/0MM7xe1nVke0fxU4bOasbKlhrK
4Pm8SYPqIH/nXfysGFmaCF3KuKAzJ1/xC2ZkTP3gM+4tYCLr2i24zy+atRHy1ZVZk5P1gnF6eLaI
tlYxzrwkZJBEZbQraHnT8p4p0NAAAmaJRUIsVU0TRQUPFYIETkDpnAphf9fMTyZR+9d1YTeoZ660
zJmxhBuE4cMMOwC/FURsrccdSzguHOOxLFSnj/XWfe0i3Xp6xEcip7vZXuHG+GxENxnZL2VESGPG
99sHNhXUsMHVnkLjpKsklUEnkAVDw+skmiaSPOeHcEAQ+WQwxxjFX8fItrJuQ1uER2drieWPIcXf
DWwjQLL5cmjlnKEme1QF1O/UfNUcKTxU6nGztU0vkQlaR5SikTIz+muUhdTWq1QwNfD0iGrMbx8u
zlTYGvYPDFstNpMYi7U6fPIVIhascJdN3B45ncGY15ppErBlHHxkecrFzvio+zgitRe4bl9Ve/aF
ZJcjdyLudWqcTqiJWWReih5wWsaBLedVImns8jmLa6pOULHH/z9IwrSx8nwN1et61u7CiJtNsDY9
oZkviIDVYohpHd2HJbjQO/uCWXc7xm821HGuubjgviEHE0v50J4J+g0IaDcYUPPDg+TSALQTH6M9
aRk85GKpBhPXKYTWzwa1fv7rL+tJU+zLcap6GFUKufkA4pj6BTa7rdpMqfeNJwOaO9ukBQ+5UuwL
L7z2113yrPnfdfKL/OoQiFkdK4PZsC26AmX8+Bx9L18PLf/rPN2UaXWmSZ8qNAbluB5J6toqS/pi
WlwPSALHGT2lqdPdlfmqPhVwggATCRuq4ikz/UBtnz3sLE1RpDGDKcUiSIkshVx2D4CDiQvwYZAd
5olZXYhSZLPxR5oE9Vxf9pEZRtQQ9PxFEguH6sed3CtfANcadejMwA38WyBfixDsT2ejl1VXh3aa
LiiQr7Vexap5tUCQWYdxkU4uhL+0AASOqprbEEi9xWqTHLORbknguTOPdUh0hPyBfcZaLYKswuh2
1/ZpfqHs25kjpq7GBLdUUtHl7OiRxW9RMa3PZkfvC4GzVL5n1ShBL7ODw0ofArusFOiw/ejkCH0h
eQfEiYPKRnpYSER8elURtb4fWy76uXQ0bfKdMhtmoOSb5RF4Lma1rVXLotvrfdRID97azaQgLvWX
PhTH/lCSP10o/dVG8Y0AsAx6xR7mVHdlXayFWrIjO/TeWAZgG7+aMxgKymGhQSfUJ4at8B4ebTq7
3CF5zWSpczWvaeOiQN5tryl9gL4ACys3Rh6l6bpGVcBM1LhH2hHnmQa7MFciqhM5Gz+7ZHG2jJYz
xk4FmmThpVXMlZ/dbiW4OTu1s786Z8/qWGEsd0ctKkWpdPa1JAPA/EZIyjQdNHbWoVn6pr62SCMG
Nxdqof19yp4cd+RwCQJMdsHen7Vm21ZVacvnlFnXjzQsDYWaxywFfQnp5B1hk007v8jDpS6IO2KV
O4jZ4ujUz2fUW09OuAurx7PwGAm/iKKQd/55vrnvgtaR4939I1J44jl0t1mCM0mbt+bPhREzrug/
OZUZet8k1xUSPPyTxMXrbpaAaXwVwBCCRfloPuLaEW+kBCRrX2yr8peBfNVqBbBXwvK4mAmLJYYC
MXlAul+T0oe1xJY8YxK/vl1RROb2lHUgPSNxS2Ge28MT3euGmgs382jpYPqL6jBCTXKEOzfg5+rm
EPpJHlYJXNlJxRAPjIEtBcp5emooMc/BTt+qVGFaSstmG2yETNGl/WjXeehcNx+rTGRe0qWJXtqC
9ApP2x46GNtUHk/KJVIPoFWMusl++Q46+5j81tf+9OmpFEscTk6yMKLF3IdnU5DeUMUlzM6g5+9B
NTdKruKWMYoLryT0H6b2mAEVjDFfTC/lJRbm2dbQTRJjInXpAA0kv9AJ11Z3vtCtAl4rIPKxxblB
EB5ucanQkVwPVuA+5QQKVEeOpkRZejMXuZuZuQ/XajqlJoRgFtZ4xHHbVFHAUhc8J4zY1vyROxu5
1Es9BBji0xNeZnmZr5WOoUmkbBsd8MpgyTR6rbxcBzrA1VyfV0IbmxUDbzbzNtoOb9YE0Sjr+vMx
2nT/SFJghn9qBNTx+BU2GWAezYyQLytv7H1obPGpiWnimuYyhWkO0U8X8C8ICfE52BZFgG6XWyyB
++gXh9J3/siq15Kwsb5qVnT7ZeEPEs9XEUrISjRlaLDeACDnVH0NrcI4LsUecUh8Ig27OP4VSpqO
GOYTEDjFO5LYnoQ1IxG43RSwbstMHBMoDRl6HB4aO4KtRxKsUFG+CDV5gvlJSWHOw94+Mt6LQt1t
OdmmIp6SdOhx45fuJRLJITfRWO6HqBwteqIbHlpxTi01O2PdeQ0W8ebmhugKWKj3MjnNuSi2bO5M
r6IwcRexdQNonptRpiqiPPNrrQ6MxO1QiqsCtJVE2qm2yMAV3bvTL7iqyz2thDOImV5iZwb8OBmX
x+7A1OwRX+9NDv4mR1Rh1SRODHJxy0MY0UnyeaCdjKFdQfuBQmUAz2QebV88liASclRTEES9ZBFE
JVf+psTWsodrATdznEdkRfNoCMyMPYCOGD56nkfTgH8hkZ+FlO8My+U2nr/IcifYIVKmTKZqyVnw
y4FtSjcyDh/AUEl3Ofbh1uq1uLqK6vh9PaxET4hkzqusZEpg8TjaipML1ghtPzOqlmFfl20gMCDb
wYfTu1JAxSGgpQwBPMfAGwztnx0CwYUm0i1G258IsPlbngHezlThzwFzzTRQPkwPO8tEkZxYP+R7
SeYJzs1PhAT8tcLBTXIfR/0PRMUwpIedbSwotzAgNy/QMwTwz+jS4HJtysjN/XXrxkWlpomT+Ah8
8ATsa/H1Jhkt8DhLwf3Aydil9CI+0xQybzr3HNFaG1qJDAEuvuHnZbDbBCRr3vI6MtJJczQKT8Vy
QtBgeAU468inkdyMo9El4edh81F2WmWzGi4EVdxJ/7pFS7E9YMRZ+SrmuYzNBzYAwtS7XSvCEgkw
lFpqF4s3FxK1XnVGfVcjNHd5TbGwllOHlQs90FkaJgY3cLRNGTEFgJg9r/s5PJDx5r0eYLLDBvt/
O8hRejbDN/5MJUmCVb2GZ2TToYQHIPvGxn9xPUzJBQEiS6SiOSqtCn6nMiFl9lDHL0C9ybtniZmc
9bkm7mEHaU+ZNitw+FUfrl/+3y4YDmHVPKFRFh7F9QRzqRPGx6ns91Q24IydEq1M65PuE6ue2vYq
iLZ6qCwuQzz7lPI3Qp4ofHXqI/3uiuwmk4IUu2CCEvNVfL1wOlYVhOYPpztDhHeB7EDd0YZTfxqO
2fm6vy+f+CQlQwNklegxL7gVjPd3U10zEbkhkxksUFleW1jgMFliEdDtOzxktFIXLwEa/J5jH87L
3rRdelI8mNRbO6mbeVTaLRcoocU1QtIN+ctIeQnj8Wy9C+IkqKfaLcCkJvcFtYSyFDHpT6z7DHl4
bOzTJMqb1tViaElNDhbEN6QjVI9+1uAoUjp/HQ2YOujy1dLF4S3Y9g6QJaTIeSEPidD4GOwrHd1E
P2Xqdpf4sY4zSkVMyiAiu/utFMkhxiEga/cmbo8JpiatufaPeJDUrSjBW4WJY8NgClE8E4nnFR3z
x5fNu7DmpccnYoCF7rU/gwu4VZUQIE5svdDzbp9s1PCByCwr2CxkijOsABaWI/T0dNvI45BkCt8l
j9qfW+GYZvDt+NikLKgCCFb/PcUFVwdDU+GNvsizOSU/R6cB6QBvplJmgwAHZ7KWdmNp4LutdROS
SFgECjvg5LltBQIgHBBSCo3nndZteJLge3llBw7hKqeeOuLYlQ47LStxvHfA/egIxNnsOkYLMxID
ogGuWo1pKupZnr6cczt+2w4LG6qeEE/lM9RpIGvIpeAbUOkyLSWSuabC0w3Q5IzTEqt3K+NtWjwy
/ksma4xrBiDQ6xKsewnrmbpQEVJdsfOJhULNreF+B5IW80JhN6smISmPGZ3j1cJepktNHPntgv8C
7QvvctXxO1AFtdjrX4MOU7Bj/uchlPbJpD8IjK6pyLD7+xfu285Sy46qnvFpqVx17JwbONcfEBVi
xMkJzAi9ud+Sho8uDmmlxxk4fqg87+6Casuo38W/RbL54NDPz577rz+qZ72TPySnKcmD3XZtBLmv
/8wTsjV9pytqyIIXFFdJeBsapRd+xBtQmUzH3rz1MbbiZEMQDOBpwGFX+zWYIKyqIIJLkI5NbyIh
Eb9yWR1nKtubXkGGhzcpScVtdjR5IiY+k83+dUeWxhVB7BadKqx4opZfhl/kP00qHXiv7MxajU9n
wB+cTOmUnxjAKFErlJuT7v/8p26ixMkhuUWvVHSVPN6BgaXA8w0ja3gwErsdf6TWPzVk4r7KLeJU
pMS1XcdJXcpUNKUI1Kc5rqoSY48bkc+Q/oBtGX00S/Wy8uIzAl+vMflHmANlNe8xKxtoGw/gqqpm
n2FVBHo2+ufaQQK3YpltrGnfmVv+3PJ257qqLmKUyTmENJKO+6V0kVMOzlM3Xruushz9jXBY7TLL
uQ3UnPwp4W6bLrcBrwaDAsQwyVbhH5F2oflUFYn+gzkaUz4vGKPOGmAHdd5otwW+WDVUbGuWxAeg
rZ1Rzh14cLu+L26+qBBLyIYzaPLHQUQwYTkoMKrjyX0o+pupYnvHYZoeVK3SFVeBC+hacvMjypyQ
qXtwsVBG+z+ILECx4NnHlw+UZeCf9FS/RxRvOS8UoYFKNC1yhqq8hWHwtk36qg2SqQU+w0BjID1S
1/KCO8aa7dl/BLtrHZ9Ykvj3A4lCK2E3qP4RT//NXlNM/N8XSVm0kKLM1OcxKxKD+WwGyN8NA4Yv
DbQZRq/6mr4YUnp4/mZfoPx5g6I5sUxbBrVdt4E5vTYlR08VSVp3lwQ2EeRAjYEsyblJzizMrwme
myqVhs/o8lT/p4W6TO8n8KmOWh3ldcBq5ZrOYBiccIanqLTimXoJsiLgNCpDGDccLqxXxCcZVk8Y
twGRBl7xTAvTov43ucejvBrTMZaPJnimkzE+v8p+8Qu4srYMF3e/tschnrdVYOORcxSajb/0tEVu
cnVVY3jGxdjhGVt5ACPBxXEgMdzJ+9uAxLyYJBVo4PvdI6CEhXWm5UeTCiwvFG0xy8M7LRo8X9Hz
3WKyaW1j5GPgSOjScoaWii7jeNVf3Wl3iYxV7CD4RrMbDGIDHQSZVcdOx6kd4bxaWCmdiqIh0BjZ
4/CwtdbEUkPLtSiT+bJq8wjQ3xqIYnmLkETBw/VTNnaaHoKFyYKeNSROR2fTe70uhznHW+6rzDvU
kJ/iaBS5wP/dR0j6iD0YhGRiF/7afFFHAxSzUYbfj3MzDzlcegIgEWfsQvn0dSRbNBGlUJYXhqjz
2Ez4huh/wkRI/zEVjQd/RT7sVmM3AZPZnN0ahXZGkM2j/6nr+niQRVdl/v3QP99Ra4SLPHPgCnRH
GKaUG+KHG74I0XZmpauy9jA5Vw60RaqwVL/CnNnxuEbSw/oRJbxtIpMB2HvbEoi+xY7xZSaHrGxD
9ypjnfo4kKTZg6pLJlaYkW0ItzxsvwJFKVZBk7cMvjiu4bFz0nBGaiNsKDdZu+O7UcHDmdpp+teD
3Iz5s8VqY2BbmhnuRpjKBCrS3/j7IxwB4WJgBFku6ikk4qZZsOrC5n5Q9Ds9EPKd5xM0tJyLukVA
0YF7GkqoIUsXRJ28ihjykpXg2UztJEWTOUHq8ycJVL//BtoqCrc915v0Z1q15ZRcnvwtoYYnXr3N
+j4WgoNUSp7Z10iG9TJkZZZdzoDHoCA8pLx/7LDBShosFuTu3WlyLke9lSaBEvgBdKhC1C+lL+eH
M2DPTOh+fDVjSk/12HC2vYMMD3i450BA7UR6p5rSqvrY/4eyE6kdT22Rm3PiDDaxUzdoQHx3JkDJ
wkp+jD9vIyqSfaS1wA5qMjbYsAw7Z9Dg2bJZ6moYjyy4vmCJkO+EZYth37yNVcVwfYeXLc7lVw/i
xfMm6aQH1biIFmmZOycTQG03pHlCSLXb16vwEl8nBWcVPG+nFm+ybbllqDKBKRoFjuRwVo4w/Moy
Jqx+eDuOiJVz/r6XNq93Q2sWSbsUusWBORaECQW2rVTiqOtLmFLYtCCAfbEPj8r/YmOG+6S1U+ae
8Lu+JNZ4VRitGdkQYujvj+Hbv5tqZm4/1ODo7feuuCWbW4fqWXybdLNQrfOKKqDc87Fd3MyTPHPr
Kg+iWl20Ox6nxvIJX1ztQdSlwYg90fL7+vYYL2tFpn6DrWSuVWvEV4vi32ts7x1WVG6pQNs+RMrd
gbjhEV7uuOT6a2JkGNWOHnKaubNwoChGV5Rb3Ti82WilnzIQi8yl2u5PdtGc5H2YncFHdnqTuqy2
Mcqk4Lbe8hEAnrA/rkHa5Tf/oLlQnFsCNBgaJ2FhgAzcjJQEgWucSzjGmxd94ALqvbO/0cXCgnHh
5ucJa3fQyFJLeUFF5mW6dZwdW0D4pu8BxTKudXxJDudH9HMVwTqhgi6pX2MnKZhIzAEapoL8kT1A
IYk6fP8TDP/TJ0ObIU4HBKrVPsAIcyALn3tiBFAeo/4NMXTzJofGU04JbKKQPihZjlZ2hjoe7hNi
zeXdGfAliDIv53lxdHG9Zxjo247gspdRQ33dl5dAZkJUMnABvEKc9eIn5Pqq48JQOK4pNdoytA53
3qzPaX14/Mod13PlXmb41TV6uZwLt5SdwKglifbzvZMv2FxTsqOWmDDgZyWAMrher25vaLk6Oo2S
lR80C/vH9vb4YuW5Mjf7BqJHAmuAmQieqzHu9PshONpe3g3Eb6hcJ1ljeDDn8PbOmZgRwe16fjgw
LTO567vGuQRjQ+AWSbi4Z1Cso2j05I7f8d+lNbthjjnJSoDvGBp95guBV842kedYYy4XHU/H9jSo
Gdhg0Hcytrh9YvF6Jlmou3A2KqdEx9t3XLUykxhlyNUBWv24gIL9pq+vtfIykUxyJR5UkcsyLl8q
G8FJ6MohFRGrfn9eQvTnL3f9Yf9eEZNG9x9Iam/KOyWhUW3RjjXcFDWfdhx2ckUbjlnxFmX27dkf
qdUzqCgZsc3yWMijx513hh0rSGr3N0feA/y7oY7HHDltDQpObdAIsCsCZCKNOCwwNBgVk0//tf6n
FjaBA5l+kZVqPlCBaSgOhwy/2Ee/aEkqzrtySr/xrEWdRrm05VAXxNOvk3fXYF3NQrJ1thgAEJSh
/CVCS/MfgwOET7pBowdn+/WhF4kCIRNQ7W3DA2m3+IFBERW77gdFt/1YXhLa5bhO9ZY4u5CzBq+N
chxTW2vGH/A0ORdA1C/fB2ozjrmShejI6Pu+bFiFcQLvzg27kFfhM3fuEJKqhZCSRXUO+DRiOHGI
pvsYRxDC19vmixgFFc1aH8dNmuSKqQCAV5mE9hnU7pXt2jpUc+NnSS6Lsn20whmYUN5AJ4lOE5xY
q0Gd0LJrmMz3GzGJL5bDf2f87vTz1VVqCoQfm9kcYlo50czRVOObuDHHAHkDOxSOZiI8Hdp5Og3S
162qGvaYJRwtoCRmuUTUew3SMDCbyYZPeeM8Mwl9Dy+xeDUiezr60zsTc81GHRAg2x/MDGenB1vR
0HZ2msPeZ7uaBv1jJKIOEomvjlfJopRMKFJcSV5Rm8KWA+858yu2Zcjec3Du1teDVbYuJ4bWamwv
zvoHVgNKZqwE6ACX+2zAiVOGax5isQ46EMT+se4c6e64qDFGuT1nJUCLODWVdq6/ONqy0TbQrSiM
WDgR0qGTm7rMy0i0rZfiBTH6L0iWWi718YOIJkai0G7Ayi0Mmln3qJhv8raTzuFqasCOQIBrHMYM
WylwfzaqgUdXk+acxlLWp8ZryWFIdDW2sdHw2Rxuu01MkWOZp4tOcfzEPiVAQPUw3o+b5cURLStF
s5Rpdw4t7CgmyJ8j7gE+6hbKfSZFAiiN+s/2G/mrMZp80OEJiaA19zk27Cx2yQIW5Z9WfZuhQlb8
U5h1TYH7Qf5a84L02tZ2Ha/xJNRdsXju5a4fuMHvxHJLddRtkCIb1pK49Iro5tUNALJIz6IJzeUi
KWJ8XQaYfv66QY9QDxaxIO+PR8yDlPKxmY+iJC8JPPnCnUALDgq4fviY+KaYlrBBSbnw37gykJ+W
UGrMXm7KZO1b9ydcOom+DgthasqYGxrJ4Ozf5d+OR5aatUrGuCsSq06Om3rYVJkUgUiUfJB3PJaq
SjCkoqMEax5fv9GesKMuqNEXOf8FAz/CsOm4DJ7sM1kcNsPJ4aoQCO7cAp/Hd5CUoj+nqcOfXQqJ
AKV8NWq0XRbFiaaIyu3fjkFRlm6VNm+fBbk0Rlb9Wdt89ANOuWHR2kEWJZIQCgRd/Hz+pfqU5ms4
iSrxgGejC44Qhbo+PJRU9k6rdJD6uvOuny/BQD8VHuBeIQYAa4GFpIIOBax1Pq1iwfBzKrCvnJwL
k9vwmVRm1t2pKU73mFF8Lq0DM6hAFI9loHl3mpV7qWDxZPFMDVqRtvFuHI+kl2I7M+R/Uh/GPUXz
A/9Ck1ANIdwY4WzhAyB/XfqgzzKXRelSgRdhTEw1bieHD284jtEO1Hn5VqxgDNgetpVEvBcyuGLy
m5i/IlHV0EeOVW7yCcWedyKy2Jq/mIDqjtXvqKK/IDUiQpK2/mDepndNSNGfp7SdJ/YnPoYC1ziu
ssf5rcdNCJSrANhKb8sg6vUoPIkzPYWUSeEECUKBrDh23DfqCtlZp9oB9ERgm7UJb1uSX4+rcpqZ
PI9+l7ypUTS2/tHyYALqOWRnlIDh9DzDP/ajrbDAHaVovEx1UeN1YMtsRgdXM3UG7iz2WfGx5DTA
yn06orJx4NRbeQ3LKLksb4cUl7ZZIHuAxDJGoHaMoFS5RHpTySaEHjOQNNhto/Tqke3056+48TR3
0/rC1QWxpW66VdCfwdl+a5cJbN9Uxw9uSjC0eV8i9IF+jk6F+A8ewSrycy/OtFhtBuJ7rvNCpMLJ
EvZFBRs/+5grhsdEqLgbYYyNspEO23k8Te1a2NS5jSNq5ctt5dNesqhRPVuAC956L4sm1NkpowHG
ZxhaXhayvTidgqSBY4eO7MEnZB8jwFxHtKPoZOtrzpgF971JsF09HXaqojiHSNOZaFKIFC8XU4AD
h5JXSBGOtEnmV+7CJvqqLBrwuXsUgrfsJFAbIN3FHApd83+ExlFtNIPfzFRDHucrVWlb84yBnvLu
kdRbZA7OYd9oyhcRPl8pBT+cHBMl+DiQ3gbm6WK31b60aFQB0avNmp1T9IDP9r4mtR011atNM7HW
xfJPCJf8YDzElj6TPihpYzTzAJfn/knKk5xt3J5/LLm9ktmEdTAVsoRHIzX63Q1z+QUP922WbVKq
a87YZS2LnwShoKx2nKdfssxtGad3gdfR//bI7M0m0XMgdm93vHw+ur8ocCD2afxoRcFbWNK3U/RK
Kp8xjTX+2noCHsoKo4tN0QZorG8HH585GzHG52NzOM0GxoxV51EuYXzb4F3OaG+sUJhSfe4mjcWH
4Qkrv666NvTQh8wiImywJCKDI+YeZBkQjyJbCcmm7/DLQLPYbKEw8edw3aByDZmiIawv4RFcTEFz
rSMZhddpklgPO3/GZNy42HNlCrvTqeL3mh6Rrv3jpFbVwWWgrneYLLzh+f7eekH+L6bHNWOTfJiN
eQeHlJ2cW4ue/++ZJdSoJ8y132WFIUpf7FdmYTgwILdbJp5+/iJAxwZEN1rY/CRMgYr9BqHaqecu
7tFAjHF/ExhYQQj/zRAxqb4p+jhxIYP/CHanAdQGY8pPFLsDcTjntX2kSJOAGQl7OUUBcqERCKH/
b0v6VJjBaQH6G7SdOcV2bnnkzzEt/Iu+XyO79o/LL3Rpjm9TzMt375HvpxIq/BaY3/mWtKdF7See
RxStrKpfcoajO3wfoLGaOAK2/FOPL9p0AUwchvrcExC0cBcVtQoolVwDaQF7wqxSq9c8OLtjymHr
PeZnf8jGBb6JQD31q8mPaCO/w/vudxzUFBLXlX/PflIYz08XatMim+RXmE735pEedSrhDrW9dRhk
WIVfnYzdZBjstvkjt2AU7J9UHfNY/lUbfRzTYBHXiFw0ZLy5IFAA70OMm7dCciZFQglefmc+Dpat
yGX+OD1Kyb3t98hjYpO90/7Amw4ieoJeGKCuqM8gfQUlQZpcu/+FGBLG76blZ0eftfV+cGFq+Jvo
eF1mxiI7oAStVaQZBW+KA6MJF9ggBXpTqGsD7X+yYwsQhDMuUF2oCDO4JOaVXD5XcDxRsKuO7C+D
vXKhymkveXVg7RZyyirr+eLJhMaJTquBmE1GmguezU1taBonp6lBW+Rjy5un4t8C43mBZCcDV496
PBAxdQRMcKheQrgHEyUirgJ1sTQVc/y5Yg5zvTJDgiM45n5BGzsbRaNWCa0ULqE4Piy8ZmFMbtfz
Nzokiefs+shcw2F94kYFSicz9mG/JMQ3kAJ0FVarBi86TKTWalkSpKvAcLMSD0ztnqUbL0aB32s7
sCc+5Ma2OMEYm68Fphoed6VK8MXaoET4J4dmnrBBikh4ZBHIw/S4VVh5z4eRSdL0RbnVOw/Z78zS
Yay+rb6FXOLplJFtoXHF2alf5x1/HvVWpe7/O8fT62IDQ7UdxkWqi6kp8ouviXIQXmjwNpxC0L4J
JlLGEYf4jhyYXpywZd7LC5nZuSK2DBKXL1k1gncj6QRdlLPtDXEOwIW+eENzSocdbS6/a8oLOw1l
geMFTfaT3dQo/0BKfKYncWcKY0VNiDiKBCGT0K5luSJfJ2NecSEu4e8q82STeF8M7tcOqyE83hXp
U2Wr9VEHbC2dy7G3h0WcnAcn8t/1+YLOrFEkZeeyNGpmAzvOa1900wP4Z4oHB0dMZ9+jGpGZcze/
Q0ZPSjNJBscvO28pCFz7AL7zSchEt3gbMYHsAKOxKium++DrubR543F2PzjRESy8NIPYAqpoDdZu
VvsN38EtJzwfJRIjtVh7rM/hPgeTdmpaoLzCNX0wmylhJvEdTrGARpZ3IB/sONX0k8brgDhldG3O
94K/ydi1Rvgp2YCeuQTtA/OD6SEBK2LMD91PQqB+Onc0U5sGwXR4x5GlaZHQjfi8mR8rDH0ap6bV
k2YOx8uP/d31Q0Oarpq1m948bz00sStbUpSHo+D4x1TEpPfHPeNnLPTfZNDgBSmL3zC8pJlGk91I
PPI+jIwShpSckk2tRrb+0FDxqMM/ImNsMDuoztRRSZpF1NaiXGn0AHqzipH55mEoXEPAJGyk4PCy
gQeQ7CNWxTnIM642CJXcfcK5ap59MXdN2xQvrfY+yp8B3hrOg5CnI1YBoa/6Pu1MG/l8uRACEz4p
xlFgYSEbDb1kM68PJ0XGFgDna1cU8KHEJplLCmJdZWf8Hh+JjrCB8MhYX9U3Joji6UFS+HLablvj
wT5lYifxkB+cCGWNXzCj/Szr1e74f8vFlfcz7J/4HBR23OjMluXcnFkqmPJjYQSpAWUQgNN0k01u
4L0u+BYXXkOeadYpSitSuE9RJmvVDO7nHhMiLZnDla+yOYir/8SQns4xuPa988yFl55HDSmXmexn
2NTpLTeRQZNmWCdBxUUV2kpDy8AqRKG5AVaTE/Ail0n73Vb1pOyANrBNppegKMUnB9xaC88ZOa+O
CxHVnUDfHg7C8Or4/h6C222ZGIbTuWWpbLd/m3WoidyfUGH0F3xnQSdikXTaq6ZMrXy5lRsB5ESz
vgfnWVeMHpxSqjCHgxo3//AYlXtwEWbWckNjXNtZcIyziQLKbzL7dYYXdkiI0M/c0kWVTHSJORYU
DHoRdwUTbXkFe8IraxPqewMja54Ej1BwAMIJo8RJlhqBK1sFP4dgwNVbFzU3gdb38cXdWuKzC1fH
Jk4NuvzEcRTM3fUQX7DpSBA+Bs5JnmwYSNU/XcKGnN2a0bah9UBPde9EXnLkjrNaYactFYU0CIdG
vQ1KMPvod/051WzbgVj+G6vbIugd1CoJy8g/Tvltp3V2++DNlfZirsASwS2DQj/QbAlcIwv13Jho
wzg5O/KlvcY2L2N6ao+pX9bAmR0S5gYSAxF90qZSlbYOTkJnH2FhPKblN9T1wkG0q5AKbp+dRhg/
Pk+LP+XoIQoYcUnZVci+uzpEIEoHLtbchM6hlBCKPkX73t2RxPGN3X4wo1ivgwOZVvC1mMx1HV1e
kFksJbhWM1hn2e0hdUCrK7jlsHWUj/Qek1pqUxOKfehg2bHI7rVLZvIDuw/Vrp0UK6nL5IDUWxtU
j26FOzEGAi4lQWGCxocWNd1Th7byVf09sdp+VOx/5r5sATOABxnhfRAgwryRx0tlkkYycsxpQD3j
c8iWsf7XZ4IHcq2DI/ZrJHeUwQyWlqjT6vqlCQ9/JsuxR8Z/n1ljC2ZBQ8Hl/DxVKEuGj7wR7PEm
Cj7pw3Adt4Jl4nXPhOQ4pHAM/f/B/WtmW3z1B7LYr6RfzcGBaHI1Ru52q/AjIGlqJ5cTAtWPoMT+
NmoOgsjhAEgmPCeTC7Wb/ZrXQPcLSXur4AR9MjTuFi/MwB/bMp4kCG1xdwhjVtK/cihY2MXgkdEH
+Q9+FENX2EoUFvLrCW1QHcuPhQPxORx5cuOulBCBu3RQNOcGBiAYaDUPgWRSbxhrEtv9ColLYUqH
+nM0IC4wcO7K8VWxlpoF4IY8Y2gS5uWhAXt45tQAOL6uhSKeX1p3wcRMzUwRxW8aXe19Rr+6qMku
MrTdrsP7mX4Nl+8eDTWcneSEukgmhyOlYNkL9tQCkwfnID1fS5yQxmrqnnAkCD19iLVz3VBUsRqO
4ozUrrHeSBlwG9Jf0iPpJNYjhDlLCvl0v9F4uEJkdf5JJo9PvzJgzBMwqRAHWbs0DAMJP+qybnRq
35qopO4R7c5C22uPbh36gLDjEIcZ9NZF6ilO4iJ2XBRCX4c9Msr3ue94V4Mr8L8NBMxNtuckgeJv
HZ4HAup06nNF4BfQ7aTUWyyRy1cc2WbRc6DPF2XDVWBrOr6G1uXG2XCdAwCdumXX8VLZo7stLUpD
5V79gqe3VKRGS8KKFNV2G5FPvRo6NwlX7TBum/0YcGec9NxuNGpFuR22sroz8DD87UVDYP6AEni8
rJbholQrTq05lUHoPOVUBg6zPpZTPFB7WHgrctYoyLaUbt+QXW0cnnFfrb7uMBpg7lDn2j+Zvp1c
HhiRzzfvB3oS49Ky3NTlTwxi1vLRMQL6RFrJ/TLDGw/0jM9nNFITtAmDtkoh+TfnAyV0Ax0Xlr87
wnJi/OykwseWEEEC22d2iP/Cf50Cdo4YTC8J4ZADB0pXbZHzyrN99OVBz01yXh6MX2d/Knyhq2YY
4iIBWz8rkRERXB962YveeUErpECvXZsNLfQIpusVXuJeCDwtZ2laBv9DgconDujJAda5cG1jqX1U
MfScIniYgbBsjpJImGPXWwx7d3BmKLfStTQYK4sZTkxDyuF77iqsngSL/TZyag2xaeHerIoTZiHm
Lpv+pVxIIS84Rx1dISIf3nuZii2lc0/6YZeIQ/9gHf2+1H9bUs4zQEmnt1hPbA4n0agnJ5hdwLxu
zDdbz6RWOfEUfm2aZFFocKg6wwa3USDmT7hH6g28V4wG1hW9Cv9zB/j+sPlrHrpmtuC3cG4oAbVP
NYajWAS8KwgFkE+U0wKA7ViQx51TfeHprVdU2in+yra4mqB1kpND/Mn5je5/Rwdko/MPncCiqKTh
T23vfPtmalX5EIWLZZUAllf96ZNJPaVjqxZXdtf4RvEB3Tmod3glTEh/SrPwg7F/0vcto4XcwDdj
NecKTbKA+cYjZZ0FJB+GV4Dlh9Uw1STaRij7MFzRwcThDPFzucF0RguCfFHrMclI1NwymlrlSMlr
+WvZ6nu980Oi4V79R7yzzWhbTyE3UZ4pXSaPVOAocID0aK1lHlonnkSvAIwqLXOyYEVDfsxiWALc
BGD7B9YmktLV6BzN/selYgj8gz0l6h10aM7kDwOQr+f6WWAj+Px++XvVhWuT2Pvs3MwVg0TOjvMA
LHRGZ+A12pii9LnXfnouXK4BTxGRASCpujQWKM4UnbXlJXAuch4hdIQreb1Tg9WqeBMo6P4eIv6n
ur8i4xGF9iyq5c83fL51v2AlAteohY7ZqKkgCWXAUx9nUWimLsLrqf0GUKeW3kaKiyOA8hgkSJJE
W9n1sZrzubqVQfNKMifHvZI976tLXoIKQ4HZPP2LMHGC7DYlHlTXci4TX9Mervqp8MSfi4BXN/oc
9furWHz6zpHFmHgqROy10x4C7pPsZTM4+IyjdlXQ8t01QooYxnBmUDn02EYf0glRnP4zGpSTDepY
JPpNPuG4OcOw3WOaEpMPnHDe4AkxivK8YqST2TAXSmdxV/9JkPy+XMv9SNg+zpNUkXcVv2/ujghU
Opw892LZgS0297g0+EB4mqGRxnWgG0P/D2NRS2qndjTJ9o57CPcB/Y3S9+nw5kv0Si3jZ8tAgTQQ
w/o86hc8/PjnGytifTKK+4nmkRxU6MMxspEStajLXHHh64T0kGtGCdI+JjrYS1LhI19nYE0FLIB3
+XvSj32TQ6BotgaAMLSsYPD+bTvGI1R/a8n+OmYIRommsHZ1RADFJs3w8ShwE7Q5gwLarWxfWj1k
NEqBUJJIRtWGWxTJ/yuAZ9B+L1VAHciGLmy7bk8qW6bkkNDXI7sKoQOflBeOqP03m94ZYckSazIl
h/hhbIic1zXaQfK6Kvb01fPsZxv0S0YNLzyb510XySkLTIwFPb3PfOT38TTgKkT66OTvVGBx35VU
LoFcU7uKXqUgCjSSkt2AXZUZI64BN305abuCo4DwNrwgxU2eHB58E1mVnw/iGsMR1A/5czbziBgu
ZpOEavjfDHW3hH7+PlDfxtCfDvtZY7tk7tATMqZw1TsQ3vV5QpKS3nj7JCCsRPLKh0ceb4EXXkDq
Z9Aoane/NRJj6dMRb4k6GPggnqZvTp8HsxDnG1otw7Y+Mx6dAOUUHGHk6k9rUPzoxIy5oE3IUDpC
QfjgrVA+q7lu02oTbJXiWqex5fZAdJteEtccHDfoD+9zFTEP3EPOvNUv9UAWYpZz2L2OkBpaxvl1
Hp2GcNkirNUTwJFBDynUVaMcpUDNC3Kx/Hk8wymEEuZFoV5PDf9zTC0mxWwN/OtcFDDFUI5SiLL9
uEqwMuFAnO+M5ua/uM6+qX/YyI29ZRYks+NeW/oUKpJDUoRrGk8e/Ab3kJHtN2KAiEB+fvSNbE86
ZWvn/iWkh5feP4rMbPseV2Jy4+qOO29Ctj5/ltmdaSYXyt4lk7/r5luJ5pBmgZzIjToiMzGFDZzW
xq4IVn9+yalM2uH6pTvpVU3+l1c9Iw0wA02BTMlCq5F2Q4XiDmqkdehkTJnIT2D4QZ+LIlyxgcM2
se3Xk6BufpIf5HbJDjoJBU1mwNXwHKHzEvPInuV5GAVtjlnNLbdGxa/tVnwC1yT/eGWUfelXaHG0
ho19JdSBM+U0uAjV1wlbmXgxqKbHuDXI9KR973hMel5NTRDyKXydjGV392s8Ng/VOGkuxu9fDlwj
CagV7THkj8ziCGYTvTi4jlXy8ma8x3yDi0QgzSvjllvYmdGA3A+4zl/SaQGlLtfwZnmdEefqjFo4
g4kjzBT3VhY/eJ5d6ObW7na9iuh4mz2Dl88kOdxiiR8SOGRL1o+p2YGsUkxgxsoiq0JrNCgsBdg3
t78Eouue3ui9X+rVWi/1sPZhsgMAj39tYlHUrG/hhBG/tuxIaXV6daDQ+YbDLr6+FqJ3+jhhz0Tw
fJdUxo30yNSuriY9La2w39Dxzyd7QFPrTtKAcNIj4I4oe2rvNoGM691yAsH5SK2tSQhi3GNe1H84
8e31iHcwX64mDvzBohDl8LMlYNGG+j/zQ74iKRP9txs6ViGPqk/6lFr13kvJr6m3Dr6hUz/deie2
OHDfPe6rsAZfZCP32pwF9leGfla9/1luEYANWvwfjEcF3f4h/wWON+UCogg+dn3hmUApJt3onkCo
gAvSqn6DLnnXxeU2vQOU1mWBrX5iGQ5X/l59t7damvIEcv/t6hUDKHIozsWYo0JoFd6CRxpCDyiv
Bc9dm0vMRkJ54aBZbfMrPkJENgnbg/DAKy6dPtjxF1OfN/jvO2RigTGP2Ik3cJN4GeIi1bVQk48j
lPrepmcHbsciv54KuxLCHHj9xQVuKiVsHHA4jN9pDH0LZFRMSZpkfQvlNuHxe+8SqL8KOL1E+3Ok
fEKm581srcRCNYfQs/f+eTdyeacY5opMMZ/sliOCFKqHhe/IHcpCisimf9SkAB0FTXDSewfULCoQ
9dCfrOvHyaDn9G5+MF1ZJfg99nQjVMxxpOaAHSAUC6cKoqjKETjAVZa/MZhsJCpkmuY4p80X9lm9
Fbk7JFUXdf6T4sgboXAO7ddHGLdqD+OtCGuBo14UDpT6q/s+REPYUVlkwjlYeBiFFSOouDnAUlmU
XLBMEPHWj1l31ij08egdEnbtFZl6ErIw/bZkVKm1NIeZRL/GCfcwbGI2ttgoV59xVb/cnnkQt98l
XMKIN8ouQUU+sKxxoDaHqhh6N7Dm78vxjCkinULWCkTp/xfTWke+ZGOT8VgTGORuSRXtMG7xadQP
s0IaSsgGQbJN9l3VuvSmmYSPL4RFyAtZiHokjKfZWfJ/vCInApiUIQfbx9qwDzzOcO8FfT2+KkS+
5woNDI8nXZAL+le2SrvOjV0ZwJ2PtPcLdVsu9iJqe43fm7DUJ1FmMBeIdgUmN7fDoNRYe4haplNX
Rvh46ebWE05nv8B1NizNoo+XvuhkjIPiKx08kDdVL6+aTJ3QdLK3/pphl/7TU194AOG447opjmpY
uDgZrxTYAtZPcRv4xmW3fWsVVyelbuekUXQZrzOlk3bLUP1jkKAr6L0HAYz3O+Vw+7WHtUAkVVpi
y076gGaMyVTJyCAg/VbROYKYcRNJA+bPiigtUkoUBO6a6clR2llruSvdLIsQhsaOz4/skZ5dPZKL
kR0tz9zzVRw9vaK1x1a/7/W7/7Ty2oSPYjq7mHghqVIpmgXSkZ6DYPSna+XbYkZ3TlZF8I2Z8w+b
S8rgh8Gwy5DtaQxKBR73IfXyuaxGyN2tsRuI5sltZNRQQ8VKxvrT8w4+6dEHr/3lKLjYkD801ruu
quNSh5C4xHkFrOo7Xd3/yiEiPhn14q8Ra+91bay8EJ9dt+ectvnwL4elkbf2bZv5ROC6wMBjAZA8
x8c7+qAj3YBwpiTAIhMt7dStJOYBg5djZYyeumtktdnyo3ZusyV1ceVKSvrk+mWpQKLRlE/lnTqY
h+Xpuuk4yZQAORlRLRZ2yIzULmrNOAaIaLBg+Xg/rUDOOSPoSReg2RRFM2YBsQN7JM/MNexSIaJS
spDj8cmqzHc3bXn09LtXE1p4Nq7PXRUBKhOAAuI1pcnLoDxjdXyVYcpsCvxl8g2wrXikKDtVjBgU
2veODYBo+7zqg4Tj50NuB/A4MNgT4KZY/zvNfAL84OW9ygjJEHzhNqpaMMOuykzVljLzNIzcCs5a
1jdmCV6cW3VRefsJ8aem3Hj2X8qom1uJGaof6GkS/GqtSi705J2S9rCwY5jnQTQUrHZuXZhio7Q6
IZAeWyfwWUU/4QTKuL2TSUsSntMI+qga8hdqN3qNL8uaC9+H2JFDBlp2J4Q0/mZKOKGmE8mqUX/N
qcJCKplUNTITS6yeEoMEFe7PLmFi5uDZvIGh4s5uXUkB/v3xjr8hsmUiV+8f/FW6P8ygQWtRo9zx
F16Bn3lAeTcsYOkyrE/1q/EOHZRaTm3L2ikvgdSJD8NUk1x2MQjoZjbshG2JP4Zc5YbDkMwJEowU
HheSqKGfzSusfnHGmjEUPMnkWM4jBmXvX3D1/JqEMGvMgUEFwdXs1bJk9ffGJPJ9iMdEkworwnQ5
TYjGR1vzS0lClx/muwTIW5d6Z9Yv3OcNHG6TIN7SOd1vNbqEYghh0xTu7PlAyg2k/RI2MSNEwF3P
riVCATMd3lrMThVqd/HHdIWALD0N8Pb9vZGgbaiZrM23rsbdiyRu/jd91VnsA1R2qjavvynsXY8S
9l0EGcirIPniR2MEnl/mb6aUBadlgQ8ERNvanN0x/Emg/R5P6RS3PwoufyrC6oyAS6ZnOsl/LXYE
yyqt3On3HaWXc0CBY7r3X//sIfFJV9Qf0qySWCwGrZD9SO2ZVITZcf7Ob0hndnIisczp8/5ztBc6
2+PupsrHpW0TSIoInnj1kVLFil9+5RzSWcHfUh/pfbalObAouJCA4rDpt+d6+lkde7rz4XkQisVB
U8HXyEnnUuKyPPCoE1QhMRAozAe0m2YyHg9zTgl6zH6ICOU8RgxUGSYTnOh7sYro2JKkAJ+Z5MD1
Wx6SIU9aBzjkQJIGyOcwA5dCuJFnNUhxzbyzQFbnTfQxaTM/VxiNtijhtCaS/aa9eKHTVyDkeMjA
aETnb6DF+9tgz7sCiQBk6TzQqzGy5HM1Ou2ftorXkn8ZhsoORVoPAFIMF1q7jkL1cKMHQsB+lEAw
rbFpKO3J+MrgghorqoxtfTVw1XXgLuS0RtHAMizg4UYqGk0iHtoMXFWEsjEV0Bh+HW6tKJyxuhJ1
61aw/jdoGxV86H3RVtIEn6P090lLfanK9qPu+YWYUV0cAajH/tBx368MdCrN+YM4si2UBuUg98ql
pjRr7DXga7m2DtKCvGx+e9tmxqdiGhglDcADsLv37gVSPNevVzEOYLi1Ny2Y9AoH+2HlN+bgMNes
+Yd2dztoIhlvpXHLu86t0uL0bLEZPvqPSyMFZtPGInruEI8Gxavv59o3a9cyjGhm5irHdGV0KRe0
zCbceOljCui1OJcKrMJd/hgAcvTNAxEl4hzj1HXXfl//joXYntAf4TFqG/y6/twmwLjKt1hfARJJ
31YN6VF5J7sZIVu4Socu2oPtZs6/kuH9dzzbGWf2ctPihHvCnHZtuqWBClyz/l4lPwaQAETOt4KW
rbgZlp/25tURfK0300RnAz4W14cJFgd/vQmsqzw9om8sZ0VJpp+yt1yH86FxbcN6U1OPgdIU+41c
ijnsvTmuuVW/SjjORWDUxCcdRLyibH7lIs1SH/O/dVAWbutwnxG8jgLnDVvEdCc2jCZRQzJSYuLS
kpCsw0Z2LnkdO2M+DTSi0+91qXcWqZDhTqz2iDZhb73PsDoBLPyRQyVU1L538Y8xwVFZcM9fJrQ6
1dOcHAzrKdpbMXYXEsR5aEAThpYqazx+VpoBAsDmB5JhVxRGmjGUYZ+iI9wyoRR1LDETpWEN5p71
5rlWMhj2dRZEiT/APHdDOX+8JbOsfdZLDQskrhxmYX14fMAV8o48xB3lYblzJSSm8SNfnnn+2QEu
ILyZY2d1YpO+GPH8g7+y611P16K0lNBHV5N4NToR1qtwG2Z6PQexFFFhOWZHyKCe9br9XtgpjbyB
ydRwH+Jt1hHAfTv7G/pMFZhftRqlG6UTOFHarJXM+0otv5jgWAhBkoButIfvAA2OWOU5KWB9LxAC
MP19O00OFhVHUEM2kiikfRC5zd4pklA9Wvcxyz2IoEa5MxWUgTefQGmfaFuk105lM6of4NalU+gL
Ir9QSybI7Fr6QfuDh6/joLfiYfhCGbPtciguyy5NgTvRcbpEXk2MmYAX9UcR6NXY3O7vbqJ0IB+z
fFIHckjDMgfcGsj+ixvH6eciEsQYPcYUEbHwQmdBgBa1XGS3xEFZjYU+gKdf0Keh38NI9gvuP3lb
EC9t9DUevMo6MccFRFjkn8meJKrtpkcG+xmeu/YMlBc6Nk+xNToQiyNJjHcKmBs0BQmAtUuHS4Pw
OVKqSuF6IfJWsDeROaMbd3AIuGFAZIjIBraSXHsP4xmiOXyHr9XSXRjA0qu7EJVqXtCHacQ18SUY
mRmr8dXmPvDwqDzLZpmex73kTKKf2lEB5u3Ybl2Svb8rGEaYxZBWGkJWT4U6ea0ZGmX8atCbQbmY
O5ulAlsfZt1zmEulRK+W3xZuB6B/4r31WurWuE1NS30OX+KWnKACZXAeS77d18i2YEMfXy6agW6W
qdeneynrvGfz18ZyhuystPuDNRyl//U9nuOB184UAAEQMwdDj5VqlfaVYgrSTXgefRWBtCWHJK6J
7x8cUsz8+sOt1/SRpoPyugJXl1NUWjf0Yd0+YtFmkTn8Cl2xfUZT0aJh1F0Pbq3CtKctbbP3+Zbr
ndltdEHzrAY30uQ33ecL9bZSdWJ3k10RgcbMQuYYeUKOt6LwiysWop6qLn9nmfj/5KlFNefqCIfW
4ARPYC5ZoJ7HXn8LOFoycHtORVIerMUCSJ+M7jji/tv8d4q8jVXpKHkYLNdzBaBpGN6vKD6C9qAY
cgkyRpgAuFZLXiDGVF32dKL+mXcvzQPW8Hrk0E+iKEMcXIwLYZGr5AQ34fTlOHoL+LUi+Ws8FjXE
RXgyU+Ikl1uHWw7VS7GLFDRJDm71lupJRURoPGfhkNggKofJ0JcQBhVdg5ZZ7zUC8ioQFCPTXtmW
qHBz2jlRYsFhhYMSCiNdGJBQieue34/1lYbIRApiyLRXf4BESIgJ3X+QfBhiGfMr4ykFyQJAYsLl
FmMe3WZ+Ausw0YjF0ZwKx3KJ2TGU1u0Q8e1xUgg0HQQ4d99Bz/w1B9kvykCiy0AqNSVM1iB2VEk/
ZfIOnT9Sy2HrLLR/2og8fPmpiQa7ONg9pINM1eTDhtBh1sGN5ePpQSGG9C1CqPWriWZ1nfc2Iy8s
YFQ4i8gYJpi2apsfHnIFN/mgnl32OwUAj7BsPjMTIxI8+S7N5vgJcgSclxlDQUE6hbjn1vp/eOpv
mNycEQ0CYGA6Y1+4hMKksIRxaDoZtbWicK2MOq6pihPHD2uCe8yAjYKrBn5lv/rdxz/T1M4k1STX
FKOemLuq2A/qa7y8uPIsZcDkiBE0QdFhcTJ3kjNPuCiENJHDiALy59JxlpjwzFmG1HSKXD/rXAHP
SEMfsDTECnM5oyrsAaGi/hLG1Xn725klsPmdABDoE5Cv0CjIwXqTbGxOIhCO2zNBcAISBRL1oKr0
MZgwyHdl4wnzAZoL95ed58Ho1DV4Ks0OhLFBRxvIAzZID6nVMaEn1/LzOuxXIJ/usLPVABDFdQjE
rwVWs3HcH3GRZjWl5LJY7dLPVTWM5fhJMuGwQEIFz8fGoAiPkmpue+pwvDxcyucTjhwyAmfjgR2C
RG/qE8xIzoBROWMbh42ET6aMJTgQo2xXMB2GF4hMVfUZj901pIYodKsb6EGIN1ichLvS7AlToVDE
AB3gX+zaZEDGEvFB2TjDJACPD0XqRLrTY/MZQe/tb1BKDiYLl/MvFDbSfyUH0t/an7yqffC6CBfP
eJw2ofdXNbXnzoQagqsGaBLp11N8NXVXHgBtYzRiNP1cYp95UkOWhldTbpfpwdiQgkL5Iqq8lRAt
65B7/aIBh+oiVDJ3bHESh1A6NjW8x0SSCTTBdNlVJwPtkmym1jomcnUVF4JNeKh+83jKjFaHcA3S
qsQPJfz70cweYHwxouaAsNDc/qdy5G0o3TzKueLwAs5DFLZ4M3RhkJ/eTTMmkN3B5IlLEpg1K9Tz
TLdxKJtXOSymyUSatLBLCMSlNdCvd8vsdr+0isWkUMKB7II4wwbIP3UViGIchji6rOxwOz60nP20
Ec9wN0VXXttVuywWw1raq7WrLhrir2nD6aHnJ2qgALulBjOhc67UXsXDWRS7jFsjCDqRW8J7YGUV
fpR8F+6b7Vm9JFVE8FqyT2LdQtxkuGtZxEbzGfbheucuOkapMQYwdxLaQLQJ+XWemdwnpt1MeHMn
Zth/su1o/ld9lBgI8GH5syBUV/8jLf+fdKemH2aOn8LVmoCgtXo1mBscaBiwVs5cPWGjdI2QGNXZ
U4cQpuBxu4PbXHbAHb9Ez6feizvuAOSmTGyDyirexdZ8CFTPxqVpUBb+yNzdWiId2C0X0obP9PbE
uLimxqJjxrreF+1sVlV5jnK2Xm0aPyjQv4aI2j5cHexoxjzSp3KeXy1Re8+2sgdOD744Ny7eqTUv
vnps90AmL23O3nQbi/RQtCZ9WGMy079rmL5qWJvR+yBbEoPz0pBWMkR9YGtSpCCtvvQ+/i1+MoAL
wFcXcbURvJbtGJuHMmXaGoRcI9Sfl25tDeIsrJ/7OC/a1HyZyfgo+fRjsTTk1UvYcrK/thOoDOlc
5WOHHzD9u8OwDpRgKx3Ojj0hYyvWBXs6AeZ/VmV4wEjMy1gG+b3m1HpsMAn8QPstjvH9uviNh49B
fToG/a5s7ZvLprtDid8Mr1LdMf0dqczBdYvRAMAxCvpIDLN+siF9uhh2Z1VkACjIiUutCR0M5HQK
KSa5Bt0VPTczMQ+reEs3sDv7rGzjtFXlftoH6tU+CnO47PYvUiAOIprpHtFibr7j+6hUN05aSXEY
LQt7x8NeGBD+Tj/G0LeKBApPzEaBIqcKYRS5+vKxnuHCJx9rSGaAGtzuJ3GvVXRif45SAI3d7RsR
9mvlRQi1ESqfvNY05bdMe9o3AcdAFmaB1wDX1uMYQKe7+yOf2NNPRsanOEVQTZF5zX6ECflLx0pS
PLzJIJs6dF5aGBmu+qtSYGZdfEyTVZMl1izNzrTpTTxKPAhaj1bmWkydtfVPwrq7nL3Vs3kvOG/A
puAV2oqcbmL0AyhOV8a/uMRLfmmBOHzJKgU4dojCnB05eDWOkz1JS7XXfzU2XMwu4xGu2Hm1wGV8
IkyFIkjSR8B2nnHcgygbK1KqALQsCHg2Z3s043ZhPqJtPsktjh10NdzwIAgJY9Kx+lz4AhRLxxRd
8z8LPpqdNOGmj/yT5DeJKkheamaLdSCbUCC/d4dz8hTGJQrrlUux2F/Q2nCMTvwWG2F6BFC2chCO
XdEWw+WIgZnsgaQd4XCt9dfaTNqC9chLHHPxhd+DBVtehYV1YyviNTaT49qv3X2vUv4K1vlUGqE2
z8eQdjktAsjbbnD8kw8AZroPLAz0w5CvxeNeSGMr+SNKaLZ0X3e+M0YmkCkJlOWPStDFaKZxOqjL
CQkZZFXWoIqMIQGuz4pIVFon3xD3FBml8ons3IIao2L21zkKv+s7oDz6Idh9kcYaNxB5hHYuhR7/
hMXD8P+AGhjZDQKECqoz3wsYzkXGrrdJ8uS/cuWXfhOB/esH0kduLn8UfLWhq2V6VhLcwte1bZEj
RpeIzRLY7rX/4pLhHOw1de9+JylmIFEGTvf5O/X6boWKbkDxgLDGs66+n1lcIuyr4qRWzY3RUvP1
teAdf5uZhE6E7t1FRzq6FeWNnOcGdOUitNKYpbtgIBulP0IEixISkrEZTx4gyomaj3gGC7vaFdat
hCjit6lRMIOmmz975/Smnw73EkkD57IEV+q0ylEkv15j8Vrd7ulsO6wHm7d2bDa5sI5UlKOcvlkV
0GqHkKjcHZoXlqGEGYfexW1DWnCKyU1aGkyulJr/EV2ACJFWwxlAgNrffX4saX2M4A9KqsAb7s/l
IkeDTckkavswIh4MKaJ9kUROgWpB4LCwCOle+0xwsW/Xjq4WsYQzs12o/D4FAP/SCmUD4i1oDnxR
eqfm+cEUOJqkTIjCVQ7CDsRbObq4z0GbF7FxPVUgMf/BPGGml0tpy8n/L5hXn0aUQ5xphu9wk0Go
AOYrcR/L9S7yOAXrwtGMgFbMzgm7VQtxmsvfMRx4LXsPiyLC4BIvMKyCB4kq6BQIw04cAU/B95YO
t6cAn39CmpkXDJ7j8hWokXCe8J7jN+bWTO/bcXnotelOffzggIh3wHklbtNthVxMWx/JV2WI4Mva
tiQ2OPn2PqBx+R1YfZLBfsZxwJ7A8d2aPhLEq5yCmbvXSG/sr/U68atho27tDQc7X1HZItxj0Hkl
q7cOnPpK0blBhRyq1NR8ewZ5Hufbhl6GAjlfsOroOHMXLTlz3/27UU0D3opCTYCs4EtEyEvwAdIY
kpMMr6JguWw/aF22WAqZNhvRuobGDUfXRb/hOGxGH1LW5WWcmzO8EQ6/UEY0bt3YzXk9wbiBOAIP
8NZI1u6NqoeqIYbIbTNfQ8eEx/d1NIF4ZGfHWvEktanw7KGLfaevYL1c5WBNyrGzaD7zPIOqmGYi
TlE2tZ/7DLsIgkEzgwUakx9WWGpQzeB+NvcVStoiayobZoEAYYTy8BsidexKpFWTOw7MQZqtomw9
nJ4KdOTv9BOVzVBvJo7J7AsLxJF3NYb57g+w/wq/ustDseugNu9oEG1MAM2cZ6IZDoRCC/9b9Thy
KDRJJiFC8V7B6t/+LsYkdXWE0y+CU1EaeCUcoWLPU8SKdbzqGaOUDv4Ee9k7cX4PHV+mlbze9TNE
N+1VPQwt1WuuITXPaSC1Cx2jWG+WgI/bQ5cwCMVDtiHagInKetUmQCkbRgDpC9AaSRbFlE7VCefy
CYDzFfiYk0a+K0s4S4kJvMv+FfPvkQWHHeTlb5DNAoKF90p2FDfA+TOZQbyjUfrnwzVDc4lUtYwh
E8W1ZaGk0dyBAx9StOL1ubCrigSoDrjqqGAdtl4JSHPLGSWIi6WKfDgD3TZC7JQPSx5or6XPUU+C
MbNm9mRSWvP4y4QwxUdsVVmomr+osO/5WrZkQj6Z0OOBw2LFu/27iwbAeQ9DYYPOWnIl1bwr4kXE
Nyx9aUML67ooBQqGv2bfezObvVT4YY2KB9uu/pI7Y2wX6FZc8WBTJ+oS+g5Zqr/YaCoB0RYK8HyP
DSToSeAOdyBWZAD4eILaVYnmZjGFw9C0kZ4plqlfu6euOViUiyVxOQRIPkgOjgNDpTNc/vr0bXiM
ISNlnaLvRnj//WXTVOTAZuFjxNQb/BApWwUKJCEG5kQxZkflnE2NDzuH6XPSo137X8q0EjERmiyF
iBqut9r+tJdcbLVBhOTWb9oZZoe98o0kdmmqKwInoi9vopmvGFBQDOH6WNKEMJWLH8sXX9JCO4T2
IZHE+4agRV1zXdg9EhoukkmOiKv/Ch2LL+qXjDQjYMQjLSQY5DsuxerkqGOTWFTmYjC/XOLUQ5LT
AqirXcqO/ZlUMDmxxIilN1S3dkIQosuBj6CbT5d6k51Lssbzc6X009RPpe2M/RcEs30PMowsN70g
Ft3jhiZOQO1rOvyKFi4xxhYmrfPv2UUv7LBbv94kqT+8zBgwQr28gcgy7wm2mZytbhlEEzNfRYof
98c3utSsXkRvVSNT8HMn0KHuYii6184LocBr7rlmmpwvW+iVv/W/qM7JzmKyh3HrIg4aGi2SZ9Ft
JcT+q//TKNoMfYArHNdip+y8BmXsCwbV3hmIv0JJ/uTTgdaVKYmGGlhN+FI/U0DtMZ7VQat/T/2i
w9RZ1ZsjKwOv/0I58j7d5C5B8xvB+dtT21RL2bn483BV1d/J0BNq8SeldEhtJl2QuiqEEMuyn/S3
imt5oU4BTvuA8WLI+oyN44dHreL8y5f9LE90Sp9nRbl3tapJKii+4EbSFnTGGtPfBwf4NY7FKKZp
25HSbR1fgkO5emr49f5/VHUPJUy9qb2YpBR0zrqwhcBFggM3lo1YrK1LOTFPMDxFx6W34uZP56pR
n/ettBFv+BOvPKLKRDKgDu5nq/POkRBdk1PMD8xcA/hUHp86XNjI+4aSLIXKcgdNQRtr5T/zOmNp
BzXDY0OBUWHnusg4A24jHntC1RptnhGqn+KTTtCGNcKovUG8hQI8dRbgZ8fTaEueKjKIe1UpVWKO
X46yIVmQCQ1Z7R6y8uB9GlUwGukuAKTpSxT9qV0cOLNMJUYopM+di/7G5Yy9g1uoKAkPNzvFcML/
C3CLlYvYriIRw5gZjw4jL6UgK8XjzurGTAEfQ62deRIFQNMSUski2/UIVJ8D238H/EtAr0eAC9b9
oBZ9IA2GTgnpEMXH6Z/90NKu1zIgROoM1WTFEntpHHPeKWRHZ8ig/+pch0z3JDoAKeJRAqYF6+aT
0ybw7zFmoVEMKNxavfp5kEwdvG4xdQudA5iyvEygyYrsjDrXKePhWhfoYjjvNYA0EdKBM71MRwm1
/I3/sjCV5NRsismNXMnw4XqtepznWHula3qcKro9VlRKCoZRkiGCHnhpHRldpeyxf4aNC8CnjliR
wMNrM8zWNRC1s1J0VQ5DpY5SUbOWN8Is2gOg8GyaUNiD4KxBA7XIp/hKZtJDwC5po8FkgA6Yu8gW
j01w9WyXFPAPz+FnovJqzQphFidRb1BK/f7Scr3WaBxSFFJY+RU5trJKDYu4APqXq0Pjzqg964Ce
sZmbYoLxrhNuafGI1Bw1PVVl/+lxarrs8NfYrTrk1Ocx/fQBZOtSrGhgms+k+M98IIEJ4eJfTYjK
WzQtVEtwqKS07Ei8dTY1JnNhbvlEDoBXOw+dMDkTaKTSRG0pNASFgq6gU0aVAe4aFfw0NdxS6aqi
1G5pko5Qh+9V4IQJvJu3FUAtfpzeEF27x0J6N339TeD/RRq8ftFGF4/by7F2GN2rxMNqjZEBzCUT
bK1eoh0C9zM0GIPXT7IbbyWUwARap1rFlyvXOj0FIbG0ht2H7xfJ6uosSAzjBV/iQiDaBpKq6zBc
HBCu3Bhe9y5bJOPTruSmMB3rz6Br0XPs+osVu2QK6HCXR8aRhsj+GuNM7c9WeeDehuJNRSdY5PkT
sLUqCWDGumUyam2NZzwXRS6CWg5YK6oZHZufKP54J0TdJk5fkTjVo5mz6VU1FApngz/OBzatBY1n
1qHS54hBx0F51v4zrSnQSKZbvdpDK55lw6Owlsvo6fa1vnAj1M59or3AXbgiKjYtgg5x0StKHFnV
qE8oPrbOZzUhpYxhnfCoIHPiriaBlsOUi7G/PsDId9oEi9sAgY2cdKQ3ARaXW3MM/b43SLl9PGkH
DAkexklONKgRmqWfO/gg/dns1PdNONPpFn2Q39xqKhpdKxt93yqrAObjpVxrd2U+SdSinVe0iKyd
CX/5tTWWmHqhaOkZkecWMfZRh08HbZw0Q6mS7nMKYfwbKYaTZ7mjJb3t49KQfe7bMhs7z1PabxWI
yfszLHlR4GFW8bHmcpUuoYYHpvzIYcsCYviWUy1hMzKb9mUVFp7ZBdFOzBMiVZXjzm4ve+4Ntgp8
P5eU9r3T1Csay3L2Bvlvfi8fYZntorxHUE5vQ3bt9w5YPHHgYL/zN7g7xxpqZ4xLuApopShiwDH7
kwXgn1xkhCi26H3fwxQJMaeBL3cyxesVqj3S6KgK9F2eAi/cjfCf9mygNdhalLjvaW678xOn+/DC
M50xWQcXNbq9PxAf3VZpOkqCFj6DvRsoaENPtnbu6OG3IpXahbq52cnvucrsXgmw1W/m++twO5hT
yyRg3qKezuhBBgCYUkl4DpQSO/1BguEu5kWW8YUvQTNBsUS/qa/UkkuGrg/Xr/hVbnvH3Py7YtZ4
wQ+GFXtUVVWJNRZrgO2h3mvZYBgpEa2lfY9AFUVkflk2JdOfEXSf/Jhs19qstgJ/+EdhRVtZnk4o
uHG9OinhukngTD8N3HLHxb+g4vD3hcAJtxXbMvsxk7hfOhmXMNDijEpYXd19jubjmDYnDiBqATQ1
+hdq/MwVeuFojlPqDUzLaryjOog7VASkZrzHvDX60q6gX8UD5MGgitYltw/LtVyDvydQh9Sqtx4y
Gx9shVNhHXenZizkz7N/Ckt+5oSwa2RdOlOb06Ylra9MtTsOjbGaf/vFJ8azuR4GbmlU2ZLutwSu
7T0g+nCuCfQ0U/jAPt712x1QJQBTT1v5q4xOEdhqzaJw7tMvRdrjZ3ZBIo85JaSBQrtgeUgWSDbF
7jXrZAP2QjdRbNoROG9khq5FLV+73Da1N6Np+dn0TVu8ZRVv0Zwhv6Tq052U7VqGM/iAOGaHvSgk
3r4lw0/yiEwoiAwG8uJ8feJnzTRIY0zp8qsp9SUHVyftttXl1//ys/RQxtIUj61VmHJiF13pXyg5
rXZTCAl/vVhSAxgk26IRsT7ePjCaFetr8tEQNRCThKkZppBJj559rpudPC/rDVo5Z2UBwFVA8M1y
2c1cfFhVFm3dLbWyh2ebSixMFdcwQt/D5vhlpKgAYR3+vFsba6EOxqbJYJYfcIxnwilv/WoVHLgG
eSuGjlGl2AMxoaIN0dDoucFwnWNE/q1muqCNTPspMahzY7CfB/uVl18kqj2tV2mX1DBTFsMLSfrw
dVJGIn4U3d5S6pFHHksWsoI6HbwBWjm1cW6bbGAe8r7vEe5zGLfbjNT/diBq+gGCXmIVmXkRH0dl
u2CHm3Hsj2c5gNWBnzg2/jgSDI7o28LMz49nGxe5IoZDwFoxlcsfGKO1WkzWcJiBo1ljOJJLvcty
4DSzhzzgEOYz4SjK6brU75HsJNxIkPxHh1LJuE8fvRYOINT1GIlyG9H/nilAB+wgjMeN82Z3LSI1
+x6neSCXiguTakHaxHu2/xSgD4QeftbwPNTMvVMNnlr/UXlpqC9awVnDbewh3VBbvLI6qODW217o
SMWPmyhCVLqfOjexayUv03ZNBiX0A4VYK0zpwXZPP/UVHsElYB26G6vOz8/q7yBTkvQ3rP/TXibE
qQ10oM/pWWY57pMZfZkj7dDDjIdxXdXLnK05kKW5ywno5v+2DLiMjmBQZN9MyzfYzIZzgXmcMGUp
50u/gWoz3c9XNKwjToClXupyf3HZQaQddCzatMEDVupuP9OaB0EI+0WYYZo/5KmqF1O3Sg0p3cKu
9MFicosCqgICkPQy+rfopscNNveQ8p8YfN1vXcwv3JZbLdESFJYe/8Ezt+jox3ZIA94r/GT43JmL
+PdYaJmgrUA8vsnJbNuxnpuABUHCZxseTURhM9ZMHqA6jYudW6BOziMVXYLcRIjgsnrICV08pmCd
XmxEaX551V9WUeJfXDV4FJ0JrPG3m9S/GfYIEVzqCwGaYvBa1o9tJpqJPG3pQ+TNcIOgDSR+Uoyo
52Tt1WFEsWJ1TEXjX9gEXuBqyjzh0Rrn51eW6/gsKrrwAZnuyns8eAUQYuDe9XWd6j+x0x91GLe8
yELsCoUzfCR8CcyvG0MOx621y+BlL60MbQlAPjFYZbiXy0vyeRiGV1fOxrodyh1sKiQuPiIZRu/G
6FXJy9Vfqsg7jjFyU/nI06x5bZGMquW+obNqVP3o0jtqOE2jeIPX+o3WaNpTeKptiYYvE0gZC+Ww
1aMlPSWtKcEPTj2SpHbHa6G6JXjUwG7+YRNge0cvW6DYEIM1rDWtlszhSQEShlkpvf1CP1SKGYKG
+pkrEqjl6fLzmYhoRaShL8NAuFKyMIjOOPCy+GG5bG6FgyalhWpI2beHz0zzAlXPXuFEQkxaLf/f
Au5heqUfLgt44wQHRjSV6roBgQxQNb/JNjf9sw94z9Bm3JhQKFLVPHosCng98U6HrbvqPFELKply
IxjhufD1cRQhMDLW2+SLEia7K+TAma4Hg818NmYvQnt8lrLGwC4+WGOly45WbYLqi3savmm8nqAJ
vQ0BjCFIntVSsKKajm2F3rvT83vGjNEtSlbooBTEa5ty7qa7RQFjk5hX/oUzCLLvkZAV2N9B2i88
9mfz7GzMfZr3mRbjldXQGfbQEOkUayl5W/HDRiJEEDz235s7AZNzuvIBRsRPtP04AeAp4H7Y9ThN
cfAvKQ11w2vlEAGtRYkUfOEZ/JI9uDkZmbiVugteV3rgD6XgZLG+ivTmfzDNRlEP30BqasW3lrSj
F99kA8mAuxXtIpAZn1e1K1MMJGyUF1pF2WBjmUpQ8px5/wfqTyQ5pzU+aa7sC/LFxsQl9cKuRRp/
V6hC5nMgwi9Z1yNISpmsj6m9u2JBf+ppvkPolvNNiweybCe59HBHmCKYBM3XiwlIPRnEVWeFjdJb
oFGY1Vs3nvN8X4UIdKaNFqBg2pQjBAy4GQ2uHiZ/9T5g2jeBzftqB/4WfMLNqOKSgEoPhp80p4UD
TaCIP3HN/yJ7WaSyiB7QoSGl3qgjZjJ2uXhoKM3+fXAZ1rLIfIOWyFrgMqgVzGYh32+FyFvf7odK
FNERePuEvH08j5mmrdrtU+D1gfBkDmut/rgCoeqP+bHsrYi2cCNakx8RKoEZuYhi2HfuIRABnpDS
jl+r9eFuDTS5sjKobL75tq0NYvM49IhsvAG//WG/PJk71v3zFrD8NTP3wB+dyDxraEDL4T3iuGKP
VD5zmMAANi/alb2iIxbWVR4GkkyZellR8Fw3emQckpNhTF0nao15GxfR2O5aVO5Bveu7WPX+QBjN
ujtXBhNmftni3eAWp66QG9cMhedSMdT9lXAWlJfNcFzEaYT3hmDN1PX4VVDv8hmLV6h2zcqKri+Y
+oj+aMq15eOfUxdEkdVsDM4osUI0Z0FfBNh7rk/XsIeutXsG/eP+KWQLieQQ3zBm+xB4ZGadp8iQ
NaD9f1TceByJEc2hIFl9lAPa0yA/Hcm/TrvSI+dywjHzUV/LeFsWdXGMsJypwEryn06ioS1HUjZK
pJnKEzWyvuCmHrXsCphHKq2QBDKUPrsEmzJktwXzyeSUxI35mZJTVRHhyAl91sgiyjRjvkk9v8Gm
KC74+qDcgYHe7KUBwK/3eos2f0PJKBjM1bCs1LhZ5r4Wl2EdSNorAdpwiAqGDvb33/x0ox79r/R4
91rxyAgda1BBSY4XnzkfW2A5txCDLYGVjF/w/k+/OT+q8I5Y2mjazN8a50g2a6YQku8osOLUPG22
sLnWCtNffmZ6tSPqXjKqs9w38BvsHco335TvWFW7PUL82USW/TjCMRyXK6uhd4LiyyOttVxeIesJ
7KfRVCSOqD6vzc1Cec1b6iYvZbEnyd/m4wuxw53H8C+0tNkhdV26PT/dC3dqlZ/KuuMNqVrwm78Q
DtxYangxaHbYthUhqcTgqlyigL+nLmelz7j0EVgtHTRjVceDyKn1WCiVnNmx1V2+xkeuLpSpqOzl
LbO8gzN9V4DlonmzzLq0yRWUPnvPUUy0prJ1WGfz96Hwi0hImh3ui8hhPzRJDvDM3Nl52sZuraw3
Zkns4mNd3RWvqY+JXjaAcyjCJsB5yg9c/y85KXRNJ47r+Pk2+vjS2KF3CdFAoY5EHYgk75JwmHz5
vIeZO084gcs6VxVXT6a+a40vGCSdalSEm6LluAUEfCHxu5bM+g6SFFt98uJ/9oEZHnMtFxFB853r
xylqfUAK2QRfVKTYd/x8FORTqVb+7aIsDQ/DYziFuGw/2BWr0+JbyHtqs2gghKa+hkglQXpzvxPv
P3vpcKyWZ3ofO4vhQA2ltFvPkPsOKO+ZqFvymW6JmKyyMhbM+FvTSJXxyBJ6RmSAoZqoENUXM5ev
BNC7BPAFn4b5+Ow3t75dbHqEFiQ7Xa5M6hjszR2+SbrbA75XUXwTu7AoLR7oIT/4lUy8EJufZGqw
zKxJOhvOA3LNkA59AilsqkBZv/yb8EPzewyriRqWzAHRogVURjJrqHuQuDfHuttZAFPDBxac0yqa
UuxVid0MK0x2O53vFESOQg8bpdi5vqGb4H+sAnsw1FxesXhP7gy8rkBsC0YMhe7kyFriooHKSi2f
sKiyn5ukAIbmpKl58bK7wmwn/N5d5tL0wbd5OCTZDKJsOZnOFWq/LkmC9T+d/Eg9iFyO+tUzUiHU
pZjlEMgxFZPmSn1G6z5wG3OqytEVbk/0PJswJKSrF2G4vuPaTItwdqJkGUqHvsQ7yLkPNxU84SNR
zIqbVBBznV+1TcG112Vp+B8W/t30PbttVD5B7LYWHpUmVzPPXDhlMSFGVO6AyyCTRCfYAyVrflw7
JFrWoCW42JBV9DHUqoYsAdNz9ucnANDrQYKb7gVXuNrmqxk69Q7nJRuce4tDijrySAq6yKtkuASz
Yl/y6ZrP/6UVZyUw2l1eWERWwwFkkD/cL8y+V1Lhi0hWdmr3lkLYEkWwYaV8xO1TSe7d7AjyQFIo
kvrQrJb8CRHCAAvFy6eJZw9I7RFPviR7Yrc/SGlQnj21mrZjbqRWILoPAztlqClY7IDJjit4S3T6
5AqdF8XGJyIWSLHW1e6LHtGXUxHoBKAOVeZY8t2bn8Cv8NKOrZ5zrAH7PAdCzQ2JjlpQ/XwcwyJ/
mUVnaqp/ioO4TWjS8+2QztG2yOGHqAltCkQA/ZxUHpUxnCrSHGfb6Fs9NieP/Ca2OW5kwGsgpu9+
fIzy3fPt+Of6SJ+0cG1YsxwNy5kmx2rZSBAWq3iqP36jE/HMXzrKIiEPHYLKhYxVwMXLCXyKOC2E
8nFPGliKIUcqvhaXloiEV1OTjyq3Qx+9EGysJpzuDgHQrO5CNopXj2VWjQ+efmeqGSZaye2CxJ90
ZoXQokaR9xxkWgWS8+DHt+XS367QFIq5DuBtHiwtmukY2whc2ax1cbq9cC9SEhQ9u8GgwPhEMnHw
JMKEd4PGjrgAk1+qFvWqsDJIp/i70HGKa56PylFGPOsKxkfAeulfK4di/ZVgGYVnYiWsYpeyUKUQ
rLOmnra3bubU3nrwLbJnpz4faaTcIJL3Mg/btgspTxJhpe9jm+uJexKV2+zg/2B9eChunzlo/WJX
2HHMJg04DWCkpq4XXbd3QIIxHqxrddt5Ci2H6vL2UEFfUFTo5FNSUbPZ4lxaLh/+AUytkQv91b1A
I/LZO9llLSctnyKfiPOyNOl8cFsWqdEFLyGCs/2hg8HPRd4yLlbqyYjgdx72nyTO6wMHKnBWE76+
rVUXA95ST4NWtLieCyK3iAdVe0XPiIyLmfA9kRQIujiA2rOXRgIN0y1TY3vQ6liMYhXzrnd8WDEQ
CQwInWRf+a6dH1YhtfIUh9OlOSAfnBxSNmYpe0VrTNXlozvtkoDMYRmTNxVM/R/U8vC2vm9Etinb
pnQLz1tTGnc8XQ9AfYem2lmDw0EXQx0V6SBUJx5soG3BXxgXDnd69l3ik8kFsaa5tSty363Vz4oE
9AswjimpLbBkF9tg9fFt0HGSSY0dEdETn/yjb0R4drICMg4Oi8rf1wuHFI28g8LePnXbj8k7vufn
Q7q9RUpIrqWMEO3MT+QteRAl2wxZjEOSFQG+iOHwlMvBAbZa67q0Ps3235HMggg6c8MupJY80szx
eo8tC46zWA4oOROLthGdrQPC/0R4JrIE74r1U6TxkyYAmTSWQ+IR16RJ0nTuGwQK7zd9N0NJJG9y
qWm3S+c4sMApwvN4o4yzeMQGfM2qKHyzhwahZCOvgpC5vxK3Jg/5Okt+JjfvjU9OInz4X0CoK68C
MERSLbQBtlmsVD0Kq/Zkrv3xzjxK0XMD2CdTZ1xPx4p4t48zX3vLz6m0NpqQqpHcyzPGYQGwyu99
T7VWMdUB+56dxMGq11rX8tGzW0zreP+h3f/2Hq7rA6aOi7g5ezlLnDbu9sR6+s9yUgP6R2QQ7+gQ
biHuXnchnBPyHa6oPk3m5tq4C8bcejtAUs1N8OsTTLKUDwSEVniL7cIdC58SQG89z+aysyHjMzw0
P06F2RnIVRpsYlvHpK8/j/Yj0l9Q71XK3rFHizKVM3oL6azUCSyU6xi25GGYjTbPipNZC6ncLT1y
N90i/PidIwOR0xXORot+2ZNmn36I8zRlN3V+mo0EvXoVfEiPj9Rq/yFYKElwU68JWAQH3Uvb2xPi
ZGnfTznRzt2IibcAsdM8sxfQNdK1k/Dr5p4SCwi1YacyTbKgpDz+zpCxC7nByv2IfMD0l9aYL1lg
v+uWUrbBhCvz4Kv2S68bGVQI+8OymFiWv3VC8I2MT+79hxhWrL1WHEU71n6sbd9/oIlKk6LHKgC1
30gM9j2vg233JTj/gBXrJ7nAZagwa2rC4rmRcEoM1O/73DU527i1Nt0/S9RPHsftcLqGM37g5uVl
jpxMjk7rQAuxEsPnZIzLDQreziXsmLNE4FSh8JA0l2dhQY38WuiaXzaMjQWg0rSW/PayskY4rq/8
2oYjN8yMAXVEIuVw8ZlO257PGQdforJmsNHslReUqp8uYfMJOu58oYFh2zyTNbPdxoWyI+1MMnbs
sVv0sytCldYZps4BbOn06STBiTtbK+JtotK/hTyzsFmnPixlR0HAtSa45ijvPLrqkRyi3fmicIAy
gVpACBmtudLkcmYUkXvadU3r3CNeN1yAaDYmTFrvRc+lRMKAAGaf+jsnRRfNob0qZR/RLkWgkF3B
SUYK+R1QCcD0U8w5YskSPDLS+3eFS8bVdJZMCdIY3bLZg9ubGsotKbi3sYx+7Cr/GV3InROcDVVb
2dBDXdQIr1lIpU0SWfetKcq2tiiJUWl5lspDYSB5VuCAxf6/x1b+N789eUvjL7PbG0x55M+Gzeq0
PupQy3IZY0eg6pNxcxgWdnOSfvu04+ljrpxDPP2PMUPg0OU6yhx7ONEKkiBBh5UohiZdp7CahVxn
oA+iD0T6hu2rUwkVX4xwPZE8MRspVfIgswixm27IgIRaDsS5eI7z+xWPKX2SfRbAKv0K3byWkbiD
XQc8HSNDncJTKhPlGllZvBJREalpW5L0Cinw6ZjBR1CVk05Y6csAHrD6s+kGZ/b6JA1q/xXLdZCD
iYEVNOJbGv7iNUVeS5fmJnGkl+kJ/WgPmiPSFto5fInjIRPHUJr8Hf1ExGO7pzb1TBHCD8uFoKy5
tyCCiyqZqc9Pf3gO8uKmPGmj8KXUOkFC7d9aFuvOoU/k2bKwtbxR/Vqyoi4AVyUEc8CaOgYq17Rz
EPKx0ZDawwzJIZaX+VpcvYFKJA5asALaMB483t5zJRu8RtD+Xcx+tzAaiCkAQA/PEc3J1XZG8JZ0
xkQ3MbB9a3fig9zz2x7rwkpF88UgQlpliKUQOv9Pgke9XhaeANtasrE5bbgTGueN+UYbYYPsvYuR
WVWp53JwsQgPZKLanYrJM70oGn7MB12JO0kGUUzmsLbbCkxb7zePQgJGKqP1DM5FrqpY48gpzmsD
XLrCVSsxGjRv7ISO3NkO+AhGeiB6QfsdwHYvC93rNldUj+5BnXKLz8SuGFEAyLzQojV57cfLO5I2
4VbDOV2z+0yIgJ3J3FfFZdZBpVUNL59mR81GlREDKs43Ra/JmTr0yeiNLWVAPy9TM73VRoQ8ECBC
jwf1bw3W8M19QFaPld2oUZqUEiiUTfQzVwAxJffWhvb1zIVljfC7Ist5nMckvopPHjFbHeM+GNTL
rBLKpZGb5WgtO6Dwqn8bEEBfFrwpV3KWnU5lo0GpC1Hj55xgqhWzjOddBPkpBwssuxOtwJqRwP9+
56qNTzMMxZ4ztiTdHQQ/7R1pGWIYKgbwXcV8ULlcJ1OVhPH3QBQdv9jAGWaO3uxrEpNQS8xuv8kF
ZkNAvgE5jOSamVV6Cl39jLjk0GE7oyEv556wYzyFYu6Jp9lXPpE4Y/QT+iNh33QgUBGZ8UmGVtg0
GVUrbl1qi6UhgiPtC8YTQsbqRVw9EWYtEnM2QBuHkGtCLM+WHN6g7g/OTqe+OpAJIOu4sU86mvsb
r0vSq2EzFLUOFpsFrHwP84ASKdFRw5RpxhgrevG8VT+LfVYjcinDL1HjCKvQj6bqmFgkzPXmqkKb
rGXqQD/C7rq0sevI1CtQRvL4JTvqGem3btZDfafW8yvsn8Qh8YMUjYKbIf+3RQh7hyA84rpjTBgW
/wQa9UOiPmVf1ezM6llOa2X0XtW1V3GBvTTUlDUlNA1VX/0dnUsiuvdA4n46jO/WwiaPBlT4Q/MX
9bAayWDbqViDC5F2F1j8iD1gyh8WTo6MiQ9EPbfW/fSQ0xm9XMwSSOzAUqAEnkfluu5AIeT9wAVK
aO6CUYv617y8VAGlf32BhCoWH6T4z7/Oq8w2lsc6Gt4A+HMN5+zb429i9nh4PiexPnm/qMBQFGxW
ZfxiXeIOOCiUR8Xa47mGljC2lCufSbZbhus8IOjCCMPgVVV6lBt1g0Tm5coc3Mii7JjavGw6sojG
Oh+Sa4y/2xw4zycybI6E/1ymwAhWBXhy5RpPClogrdV5SfuK0q2GlyEsgGeRIGHPfnTqcr6PN7EE
pvzsvDIZrVSHFDVMa/OeAcJK6Aegyugsftgawk73l+kol7JG6kKyUIinzFggga28rEWYYUXfI6nX
LD/OC4d5LkatKG8GrBloaasyyIuN/N1oi1yxGFsqkx7NyKKKujPyqsJzH1u7TywQPdrQQ5gd2EVc
YAyEjMeok1jPCtBGJzq39h8b5jQnkOdzymSC82aZjQFuG1zJpFna3kT4NSMWfjiykZv05gSS6M81
QhbSeX8kDSMBskTWxAJv2EgaZqItdQ9FKd+fi14ant9SC0ZeoUmLlkd7kVXVOKnzpwQlh1M5BoKW
2/b7PaL76/6Zdsfl/E6TODmcrT1mmVAHBOTZBOzmlygVSSSke+PgvDoKpzlHnLpZO7GmKX0EIUmY
7/2xeG+ctOWy/7Ak/nu07pGpPI1o9hUsOEQgusjBa49Eq5YejvXrjmwIUoabvUNzVYFj9cFDwgwQ
x+Ndo+KOUatA+T/m00VZlD62zXQF3vZVm9XMEL/erE1WaX0GzFpEdmgauNFy2cDAFcKPERyM1U+c
AYMW4BEQlkV0qvRUej4zFwC8KRXaadZd0c1fj38o1h87VMIJoIfnUY59qH3tSmUiOZIp4qvMLn00
xS+nI9Wy1VTpRQwnf0LFyY9rEm66CZ3iXDdx6iA/wPWXXy7YRDfGekZ8A/udgydOG/pTzFG2T4CK
qRUnRhf/nOOaG7xKNYgmDJa+gcEOyil40xmZZYUmJjSnd/4R2StlRN+pqUZ28Jj5OaGOR7Uc5hNO
rqOQUTXnRnW4tXoEDOINTn0dbG/2uFbDIb655RLSQCqQUPAnNLY118cZYO/ArY/dHfWhnEkqhZN3
TtIv8gbd7j2R1eUf09VnUMY2SrfM0TImBsPUgp5YG/7tn7C+kmYVOmmNklSXW+wQ7xkEui6crpFL
pGGyWetmKh4ZF4QBsLkPTQrO456WmlfYFDEj1BMqpInI+qczrJQr39OT5vnJ00ZKlDxUsYkt4Lcf
pESRFRXoGVoZMQkliu2P68YMSiYDe1ZI2ciE/r9tkMvyc0qsLb7nrU3vw3pfS+Ccpw6Kepw7J6+0
MFus2WPwtlGgYstvIz4r9RvS2+72jcISL76RHFC0Cm2eHYEpZRK2owZl3irzLzQp/w1/QDVNEApu
TziW1q88MDYRC/vWVg/DcUywijzKg7xt7E2+KTJM1zS2ZKURAcFEbixHKt5EBpaRT2UFJNMhf0Y9
G5+vPh2YY1XpVM5wevGZILI48Q2YEJQ47QZl6ZGqaedBouuziHPRUf7yNx1TU3kVDgTPgrBez5ty
ONJg5GdaMwUFNp4tqqPy8jO6IuYvVcxOFytecjPY46fehw3jr14YSA8NwDEbr1znHzi8PX8OrjdL
xg67zH3lfiWj2gHqAtyp2YfXoQ0+ZmdIHHYN7yVCRluR2POJo0OC3DVaLnMceJ2BLbOOkdDXVlki
bv3b7z0KnwgpvIBko8smhZdVwAlN0odc9/AbpXZR0IfyDRFRaNqIIj9UauGwIyRVVo5ORqos1CHZ
LThlCgBPUhR9LuXMW9vviFdzFp/I2/eoRAz+WfBHCG3yvYf4Kb7tBZ5uF65l15ziTcwNNEynzGgk
NGowpAmunOXWcmCyiPdatzWnaNlZnqB2/NB59z1sNQXKetio6r6qLonETDlEDDvBW6oAyT2NxYjU
bpuLcX2yieVZ9BkIX+mHRP0Fmrf46HUNG1YooUdetI8s/c32H9X2jQZJ9yMIPWG9ChcnKzXmXNhf
X9BKTDVa8+d6O3+qntpfba6UJMhi8noDXOaTe2BNq7qCUOjCMYEk7mvYjKoH1oFlEqP4w60TdRQx
UjYQl7QnVRuHQTi55jdfYd/jPIHADfyzCknMurgbG1m9AHux1gwwAZVYgApQ3OXH+Gd5bw1gWHkx
a6aInG+agQAHLMaAazpUCBSzLAg/0auX1QpgEJNdqcA20BM0ORq06kH1uM0uw2GTnNXDrrZqdbrj
RmY/c7p3LgqB2pW8K2WE6Y25mR2gn1Jvf6smdjjwZTLdQoxvMEguxfDZrnnzpbDZGSbyisL0Qs8E
Qj+cSZp7fqmGwE37RxXC02joWHcbYfuCs79zITAacES3frEfMnawRpb2IKIgmVPmr4gX7SShRW+L
kPoIE3bHEMIKaH3e0jV6DTQ48WkkNvtTKuk2cVatlazIqZ/vAar5xxr1wNAf9QaAnx2hGXRS0Iip
Vl+y0H6ITU3PtYDHkLx+oslWj5ZE7A11g91FiDKes4w+SFbFaWxLdMteUIRTnIU2+i1M1beGaAkj
kTtLqj5WAW/rQXP3f1CMLfKn+MQgiSdrwgOOIoXxW+wI9Gh7H/GP3D3rS+nI1QNGWg/Jf8d2pajo
64OQxz/Hj6/rxJt+crmQo7bsrFRNDRNqnz9V6zuyp7Eb+gd0PmYRL+zN8VK0NvR4TenyRKUSzmhT
BugiI1/T1723suPyrIbwG1Yq6RvwjZq1ZCSV3kVp0l+UHq2P4tTteSmMT/6ylsrdyT2Zqv8d2f2H
j0rLgWzgkvuvKKx5/orjf5OjC7jp7Caf8AtVJG1JKixtXuMRPcozABatFnPL/MFeYQCjJQrd3uOx
as30ERejEeHH/pOLEdYCLaTJa3iI3uqOfZ7LetkTmAeuqrY5A0p6HAGh8yx/OrViXNMW2Ub8GBoS
fOsfVGPoPJ/zbwxaFGdvPMycq11XqrMCJOudg3sJv3WaI8J7StYYKksT+aUtzXY1UQhNZTNAmRiD
3fhfMM58kAZa9i2TCx6aPKoOSd0nQ7SjMaPOw7Lq0ELAcH3XUbzFPAf7/9m9CRcuI34ThldEpImZ
Gm1nhWnLp/MNlUs6iw6S/0KwCh0vUew4AEKPgtQ/DIfLY/C/U5IXdVnTgIb/Ov8b/S93Ij3JIQvu
Jyv9vP5tOIvf/R/CfW34KV8m18POoqDWhi8xB0TicDgiJW6Wgi7w6OKTy1SY94Fa8gmmdugL1hAd
39NlTrncFKqBJ73W9SnW9rTSCeHMy7gxIJfDmi0gaG/CFOKaU35oYJEHzzLIeKoY9ynNWQh+/3UX
+imcgB/zcRL2924HDQ+5MyuCyJkgS++vV3SgtwKT6YJSK+xEPoxNyxGFf6cIxKbkf8s05ImkEGCt
jiv49wt4D6aUE9s80nGIaTDNF4bjML2r/EPygjYQKGAOW9IsCg2X2mjrAkkGtW8so9qlx5w6ey7N
Gx85OFzxMEt54XyocYRP3Mz7yNKEFeSjsrymMqII5xJOZ1FVpLPhiE72rHPDaI3Gwk+qcsr3Dwbb
OroDY71fnHAgazD84Rdo41PM6opggzewL+guFp4D3F+Oskz2Z4pj/dXmFBiC3/oLEHsqav2Wdes6
7NyMyn8E/GYB4eXxB24WvNK7Z+FzVl2X8sx9a9G5g7ccC3Bw6blTkAHQL1w62MMjGs2nvJ7XLvcT
3Rf6LWFLhis5CespCaDI6GaIzlPdgNCZggkKHubfRYiobBzLGkMEH2TMCsdgUYYQ7r3RFliKbLtA
Lpw7P5HtyqM58fyE5t2KCFJNjsHomd9WbyohhlesudlolNWWMYys++kV6f1eav57KJUwbblBBX8i
tBAtWIaI0ehAKgaQmkrfTDX6bz5DWV4Yc+Ne8Wg4ycyaSkpDWEYo3Jh+7TyxJRaQOwk8+u9cpNP2
4ipEu0dTByN8FWQeTJETNisRgUhcMe/FwldjJMWkS7zlEsT7JacEiz0S+w8Z/ofruwdO48qsICSJ
FX8mM2FJVka7pR7oQy9onfL3wP9QzaBgTMO+F6j1YxKEwTB1qwRj8bnnsvhTYk2yMAvl+05R/eHg
miGNmILlhgHnjSbPL224XZ8c6AkHlA+tUfJTidunjce9gzV8e1GtVMkH8Wl60e9Hfw3RjVSTkvfn
1lmGusyTEbmzyk9Sn7ANmx/8PMQPQ8xrmHUiMLWRQNQ4iktLwn1aPkfvRXU50oSLFhOxkcYb1pQA
Q8DuDhGrwcBdpnD02troYPLNHV8cDrR2W9VUj8V1hiqvq3mIlGP5Kx2k901KpWNCn1tVG96o0//h
AQM7mhi8GuslWe0i71zXybZ9tlGfddHm6/1Ig62At1nTGcre30H0gEhqFds/m9jmy4dKA/I/Yftx
oHK7uroQSXYO2mXNAMEdBqPTUbGIbP/zDGGQH5NHkaBopVoLXgnJRZtWD57AzXNCjDP4WehblyCe
iIgMgQlVouKcQw5lYqBUqSn68nQN0CZOxaUggqVdsd6iIAdObZbCmggXvDUE/62cu4pwgwaSgYoN
8Qv2sDiU2NpjXdc4NVTljr7ufCJb5BMHhxGrsaONidItg5z5aDigKtYjiwnDegdW4+dBc43RhcL9
kWPMzN5YIcjx5FHlzIpgaNDVO1HH6Pb+qmcms04K7Zt+2ut0MD/3u73FRwDQJp1BAvSZo8HQdDEi
leNCD0AKA+wT50TV0EhD2SaJsi+oMqP5Kpq7obdh4v654/1xyMIfjnuDtIGatOx8VM+/tmbFvpzJ
y7RwEjUiVMssPJ72t9FYb6IMweic92mPXufe8ZQVQlvlMQFy6iKRsHJEApBGnsKbZEYXbHbyRNXg
ibFJCCaDfVGCgrLfoNAaszC6TSHlZUgfopa/pCQF2XAEiez47vVVPpjC/BlT2TL7CuyAc/mmf9Qk
SzYpHIL3MGHljkYRjZpO23tTBBN/VRNDpNSszWslm72yQKjgnDsnmdVGr/Ubmuf3L5Gv9LlRdNwz
ClSgbDdTS+3FK5adByBqESYNcBDQZJlUnVsXAlzesO2IagbY1wzLYo7tbQLII+jdgLd1PSOatGsJ
BI3flZfC4PrzFTZd/eh840+cL9gie3aX8tgz/dmd2YWUlxeMeDvdtnkfXgKeX5v3ZDJ3qwAjOL/+
GYabAtO7CrBQcFc0kPaaYDmH92q7P+8LH9OGsEexFtAPZ25luzsYPOLbSayZObxmebQJocJcZGOQ
7cQO8qMov4d+WexVI1+PprRAsDvodeTjXJE5RLISc0poloo7isdXxtQDmD1K0HH4BURzEyF8wNyk
YC5wS8Tzd6wkOQTM6EeoI3Z4PwxNNNNqFDquKLy4KpkgKYjMYSIHIJvyTA7+X/1b9i1cAIKK6MLn
Ye++qfOFTaKWdyjii9E0SmRuNxFZlKTXHEK5KyxGbrdvBKHci/4onXLp09J1EvJfogoIwffF/xcT
GD5+l7tb0F+Yor5vccgu4l6HGASnT6jf1P9Rkhs57CvQPhLCRc/rUvrDIpmAzFiv9XdRr3AaiPU+
MotEDruXfa5mls8LyQ/+Wc6QhY3XqAXTWwDKEV2TgKFljE5J1H5sBUz6kBsvKu4L6C+kSxZHchzp
URMLjWWPezg+elYsUyqZHzsYJxlZoe1iUF5lxyske4xqIgfZ0qgZ4L5y2sIgDIruL13SXeS47IX6
LrO0Pkh30ghxBhWMEx/EtM39TJZ/45mFLu2abDhHvlU9s1ffcWNspOyWhnL86rSncPeBsTKiiENq
z6XItWSfTq0wuIJPz4GLHlCdLzSGUBN8hsr+2ZUt3rX+6W8gQzmqoA+G1qEaxBdTmda9fQt0ptWy
5IuxbQXoAoHyfs1HRYp1OH6ELNE0DMg6x9WF1iiIdzexeUefbsXiajK6FPU8NY1kIzu+sX141fxn
rYKKGkEd2m+pVjMIIQfOPSCmFwSw9z2aVIvjbXx76ohe0L5hGIAHw8j1q3CMPb9rV3h9XIsJ8XXv
+0dYkOV3Zf1xfLMcJPOkSdb6jP+bYZPLV8wAw4uWz+pluWgkW6dSus0J0NySPalYX4nWg04ZeXgK
j+TTFc+Jato043uJNqmea4HYSJyJhFVDvh8EdwBkHf7A6i0pSbkBs0mffGe0AYcaAHP7ikrEqlx7
wLEYwk3VJHITV/J8W9driOoT5mpwXf3KM2NwnRQgbAQjtsJ+y8SUZsFCC7FgFzU+WLbfBj5kQJLX
G3QL95K1Vh6BR5SngYZtJcoBhdXzt5ruEfMV65VGro3JpfxdFDNn3Sbgs12DWbokM+LG1VtjEQjt
y/hyxxweClFDRrlx0DBBsBUZctnOnkb5GgxiLbp2vIRpXIVFAjUgYNfAMLJl35Z9j+alZOiVyCu/
+Ea61GYRaxNteM+GLT/MHNPoo9Z4fJUYD59vkthEF01+R+nn4gDlKzouKFYqjzRjDoALSYHo+MCf
YTQ6vsFsMe2cvuUAHx0a5OzDRrxl+p7xyLdmFJnEW/bQHKBeejr/ThFymT0CFizrpiEL/iGISdxw
3ieqGyFaS4713b1etnj53fyvquDnxj/zyPkZqdnrB18bHaKPzjcUc+bz6LfkzEnCYwp3FNSDClu/
0UmUa5G2UFsU4MrEWBSHrcNtFRsjLs8R+arnmM5FUZPG/ImDWmxVWVgvCKrHuA6K5yvG+IOsZja8
BImwNqz3kugqc8R37OmUBZO4Z5iFG2hfsTN7lA14XZNnHXCoD3LkJC4lXMeNRF8GnFObC/DmNb3O
zvHQPdj/4bHF+3NTMajb8HLOKhYVGRNlCksvoyQfmEb2utw1K2aFCnFG/Hf/Kaf4fXjYvBBZbO+f
0OftiWDZMDQoQJyvKcwRE2mBFc8YggAKBNLw/ckz3v0DCssDP5noiKcpb64hn50kJ6ZdV5QlpRxK
kCQnsQlLOefE5FkBcGan/egAa+UIK3dsyL6i9TA6yQ9q1vu/o15tJ57ou0KXRIkvTDVPUMaqbrdM
mqDvlxWVKYF7D4rsKJZ/24/9gsXMpFxlu7g5Pg0eS7cSTlz8Q8k3UswDtbnVFNUC1qW7KDoicOfn
NhiB2XumGVoD/Nr/XFS4j+S3PfOIZSdUZ3zRHLGgZ5crys5Q/VnR1NTY36jdxnjhlrKssXequ456
xRfGbYWUpcJvOMMkjjh5LIAjNVXsDwriXdS2jvW3bgfgagQa/T6FPs/0UcFZjqrtIgcjW1lFHjMr
a0dizC0aoNQjKT6vBjn4oHGr1iumb5Bof1ytjb2G6YtdBAuWHatbO4MWBHBfgiozKSbQoySMF4C9
wLyltLR/y6AeH/4BTnb9D9OF5QVexWYBxe+rhHz7Ex6XFEOdZxUvr67wDBHqm3I+n8EjVYDu0mxc
wbT3tFP3P7rrLDAQFZ+Xnp7ECYSyRAnJcYjY5Oax1qUWum1yGPABCt5+D8UnzWd9Y5F8tfjt6x/7
7ZAkMzVyd4J3npemrKTrnzi59KEahYj4D9VnbmJt5ugnLgm1bzG36xKwNtjKxcg7vLCewIgdDDiJ
MZsQ2p9YpFi1Qf6fq2VDw4ObEsDSwQkO2KN2fk+b0vQ6zSa9qCtutkatRwpDI6TcKU0qRmanj2gV
8sLWNhgnSOg9nlFjuWxyEndneUNuEkCXIdaZR97YJrTthNYwlubD+iTWSygf1LXypsu6JrdZSWfT
/VBe9zkEDNQo08cYytYSB8h9Qj9asafs643snt1G57KpcONd1Wzg8Kgwrz3X3+MfXxY8tZEnGLQN
Oei4M/YtLrK4GKKFw4qlevj5k4rqhbX50eLEA5MqovdcIgEk8QpnBGPHon6oMINiCXEZ17LzLm6G
aWkgY33x31MRAmpxYU/vTNmxFiv7Hwjt8cq42R+hqnqNK9JWdyOUvGL19WvmFh5jpnRmbjAWB7K4
DomDLEmscY6+OfV1tW3BSjFp7upzUnMGkm0/ug7jPqseCvCD1/049Vb+WLNuFcFd6rq4986DIf6U
onzOSznU7W6WEYRLgsdjMJku9IF7zquXe51bYbhSmqfAchhLvHOxiE+ngNbYArpDTtIVH7HMgBld
jBGMrjKkVLSko002KfnYjo4tXCsuBJNQtWJHJv4GGy6Yvit7lXn55iUk9gjXv56PcsdcwhQyAMGo
NWFDTE4K7i+BIeJhicOOAFX/92+6XUENnXgaqOqXYlRW+bQONtITU1SiqX2CwKIeaj3ldz5leFZ6
nbPxEGVKWl8N1CD+xWjbN6FZA6T+ASJaHXi2IfdWnOLCZuoUV4DcyHYONwm9MMvUIF7nilxYg+8w
b/LXJ5qvXzGhh3Ktg4v7HsSKf64O7yMJI7rQlIh0dwy0GIsMQvnXbsMH+kpQ8Y6+l54MNNYNyUhe
nxhDpOTHjzb1sw4agdoMl5WbYXxYkX3bmRgf0kmqeZ2oA2JEligJipWYGORyLh//12+dcQrUEXKV
ttjablZPbpVVfrB44BN6ougrVudf9W/Kib4H90MtB+kJptNfavqRlb63wZYFVfccJdBxvldesTNG
qXMHD1eX0H1nEVAR1pGyt8JKfm6TrTUIr7GjOM4XdFH4D5IFCh3gBgYsQnjKLH8kpBLzQfJ08TU7
TKSMeSI29WgUPYxLvTvfOKGjrFzIJMzVj8+FH/7EZFFAdybb1CwtdJqV6HaCyEBJ+BhVWD6nCXKo
iq6dezH9tnOu4ArynfDE14P6jFQIsQ5HNe0e+1JeKKXL2q8K/GbCt65HukniPd5Ys542z21sUg5j
AEwf9/mTD0Q0dfuB6VgONKTwJfdam8QhiQb+mSAIpu33oHlBGVgP3ATAG2PFwc3p0DbBkAL6U+Ow
eNnwl/F8xHyY6mB1BoxcGWmA6PJQx+eZuVMJeN5fn7Gr1xZLl+I3+hCiJah9UYTiX5lNrwUBF/5D
armIvYYDhU5lmMLc1uSGKfJGdqICJXR+gb6xRMouLESiEs54w2xHARR1VrSO3XtmqmXDIPrwlbbH
RajxaxIveRb6hJhTt+cdfv+NBuNKg1dsXTKbYybRNzsfpzh1ofvHSSAICKCywwEc/CRjlwlfc/dQ
0jlMsJ7NUCc8Zb5LSVs5NB/p3Q6wmJKLkMH0zwe2R2PJ47Ok9L/wsK/gZNUW+MxQ0go//RCCJUDO
AcW7nF+FxvjD7Mj8Ld+aF771r3saKzHq1ltolPJSmsmDXoQnbT1cAY5ME4U9flrCu5x0whXb2rRO
Jjl9tNSqdkQKJCu5q3d2AqE7PZADq4zb6TWuBZ6NZIoC/ui7LMyt+/mGjsNSkPaS7V0E88NlzE2w
YpdFWVkN9nNRxNf0X6PLEyXYuCAk6rds3x2KzgLMQrLd+cfJ5ybU+t+H0j8/8wrcy9QALyoKGDi8
BSdChkvwvrZ+G/uifOfkOmBVpLyQZHGIE4CNDG4wXWsVzS6UTglUnFI9kGToRrvRdqu0VeultkX+
JVjjjn32VgmPPyA2AaJpx3+KEoVfw1VK4TSPE23pJDIET6xa3lwtJzq7G7uHHDRFeWCyLme0cLdW
twE7lAXqqHwf29Sa70bRV1J9EmSt7ES3vcTTP6mT1eckilgdVxqEasbNZB8Uv52vy/t2lYyABQYA
vGRI63qPnv6tNKoRk2oKw9huR0VFrZOGyeJbLSgeIM2Qi4UCHCnYjRInMsAEVL1Lc3NRLn/2er9c
55oMavlA+k+ox408AFJ/olGjp6W88f3NJd1jsKR8s9+yT/5pkO80dw2+xj/qAFuR04Ip5ErxUBo7
pGzIzeQ5zgGLzcX7b6rg9oJdw4VdntpCWOS8lIDfGgNKeax5OqMa/FPVuzZewOKlL9BMtLO8jeQJ
jRDFuL+bwXred8mr+7DlyaGGJePGI9jLKl5p7KBsQOQO4NJZGIluIKyxC20AcQIhYc8GHfqd2VRa
8F1uagZJxAFkWRSFT3Ca5gHyOp2COBg2FcGWdOE8dN6W3pr1pZnF8UJZvmzqcSmKr2ab3QKvly5x
U7XCsYFSivpTiHiO6s1bpaPqMp48DzpLxFj8HU4SE5eLzf9SaPXTlHezHRs1ZavAWPracG3S19kK
KFIf1WlVi2FMiGKPVsQt0bS8i3CUa1+MB9ZO9jEuVNBMx9cZTkVqO0pDH4cvg1dP7t2pUHoR0of5
6hSNZdOADVy2DUS4d+Wkh+XBRFRBjswc8aJU2FTGuYGe0Md1upkxVpxCtN/p4mpFDyRDLBs5AxRt
oJroKxV5vEtktkWVPKc9P9misgMRSR14/2dgexhC/YRKLs+lpr5QFmS+2hftjrOO9Ee9PylBlOUH
PMYPnH11DFD8sVlg04ZfyvY5cnxGM6CuNEbOBheHWbfoScPO/W/wjgxXk8l+2YaSBjpE4KDFqOd2
nlWbJhBpxeoTspPtfWxiLKXWPD/eCfInkGrAeXpZuWWgV5dWsrJK+/6UyeewVtgwgTrRZIfX3icX
I7FcI7OAGYwMYZ96ue/Rn4cHfIoedZ1Lfk5OIceksr8qpDaMGfUBuEyn+4CVjDpWWDR725n1FsKt
g9TBm+gYwpxU4+zaqUTV8z1Y4tPDB84q8UQ5qkNrlxn8TSoURfdBKxa1dxUCwLGAA2Tn4YMmWHjG
YZqAoMrYMhNGW4ghY0Dj0f66wr/jCLO7XcC6No14Ujj+iXn0bYVdJiD1FZZxCeCpAOICqnXDvgzf
wLpSz14RnyAby2aJMPUQtayGSq66SBjViZ2RwStJEVbOJQ8d9lNXJvguJQliDMcBtI8ol7c7+eX8
BqfieQldn75oB0XrKh6BfROAwIspgdPMkcW1V3AjhUF5uSEkiZJBgc+R9U7z0ozb4DtmQcD5T1n0
xwPRr12jRy2Fduwzsk4dg2b6chVKqkad5MZCbnNvv6mdtH7TRFH0yPwGpEeVcsLFUVo2nxu9Ryzn
BBHKatC3z7IQAe+MNFkWCDWHEuuaquXDansckPpoFoPpqKR0Vbu8I/6Z8yipJIIBd+yfnHptPdpk
kL4hEAhz563VGNdsyLmBBfPMm83lmtV6Y7zb4rQroW0yCcaRV0wQZsRIGTrgdI9Evq/kTdxbVM6x
m9+CkVSLjiRuZ9O8lH6vOoru2ga6ryZJElXEbzv3NKUyV6YrBA4/DkF0AQwmTe/gIDi8MLN/kJY7
FusevV4+KCd21fgzJq9Krw2AkiRpuHkqee/Lx6Xq8/84oBQnFSoDI0xQBNVy/8pvpJgw4lE17cuw
uJZtGrquqctvqdZOmdMcY5AhCBlmxNwqiMIbprS57KobuNjncaQomYSHW9HU7ihqHgCUTjvBRHtC
d2boJEP8pEOU+T72hg80+H83gCGysVAv6qX6OhX18fAJAEEe21Mm7p11GK8BY7jDvnRXXwLwTIfZ
D9/0AUOtsc3CYbd1zyNudSqaPshkc80ldies+VNkhgK72NpvQQ4hv3w12HvuAZ44AfQZ1DL0iHO0
S0VG0q8MkKxYt355MWeZ1/IFr35cLRvFRqlfObeMbBIOBvTb7R06dHNoQh+8LynSJ9LNYYFpaK3o
37FQuLY9YS8GPHaXtmgQ0cCWmhe2Lh6zMEYy+Czi/OT1aqwBIOyRj/qh4U8OYvvwf7ZbCzgNqiCz
CkzLerhNliqtIPR/tmnQ9WCTGS08T9e9I0YlrV8iofQqrfGSrnPdKExsmbb1j7bDx46qsHXn6JMM
2Ee2XbR6FX+DrOKEWcGxDJUSAq2KFaKc3If2qOiyo0VZV0TDtvVPzatEWjfu3pzNVlz/oF96AQ8m
CzpoZJX6XmbN/yxx5g000v373lu4oLlv95kv3v8UdprhuI4OM9nb082tXDPfHv3duQ6zo9lyC7py
xUZL6i6Q37V8oexpa29QVRHf8KZdX+rMNWBReb1ZsEdOlz7h/v4tUqDujwHvTNa0YaEPezCmrpkV
e1bcoIz9fqHJreTdtt1Eu57XtRkIO/tdbsTLqVk1Z2VGMmhpmx1exDXm/Z7zGsx0qUgZVmt0AOfN
XoQzQde1EZH2Vc0y5H3x8biObKx0DLEt6JGDaLybOElxD6w65ofNMhlFIlSPcYkQg3cZIPruDoEI
4xgHbeAeARGMj3Ip+x5ALn4F84Eh82H7QlvsDg8RC6IBS9PNY0JD7KTe5KXA4Y3/WiDs0omVzvL3
eixiplXNTR4n9i6Xpx6KZFz2CnzCcbzTs0LS4DDFBQJN68AlRDcm+p02UWjsHucD3GX49nBCGAjG
k45Sh/VFiY6csYD96h7NuOUTiRRTg+jKxScRSPSzu1/D0rM9oGzjqYw8ORn4cSph4V6bOImnxAfL
3IB2bGb8QIK05NM/dcFtIt0v3jhS4cX+YYm4T7w30buzWHDsjOYZ/PosNsr/BRgtk8Qb7YoD5OnV
XacFjclXNwrPKh46de5qLrhiqdRVsnBwDkXMNouRQcq3ROnZyns4UjjrV/gtY3SJWexx64eMyHF/
JQFOu6vwunzkihfqeQatgDrfP2PluCDrjb4U5gyqqP1As7wQubVUA+48aDUy0cnW4MIwJvzRG2sG
XHrVU+szZnuyrZSFHaGUNrMNu0+Q5aq+k7XpyWCISS/NbcVSXXEE+6Z+EsnIU1hBjKxWPGJznWIh
BhVW5P+qxRtUBOtJGXH9F1xi7YYpmxTdeb/zi/nZr6hY3CSjOm1321WCgOzo5pJPTXEKmg6r90Yw
FsJklWw5QT6pG1xrvm+sZ4R8gXXyfqj7lKKMInQ+zJ3e6GPjdk0cT4U/bojYzwzL4lg4EPF4kMoj
9LksIr8uPCEHT9u8sm6yFK/MKKdxE2CC12kYeutEgBp7kFekByV66GlXINrUWF9opDt81EPc4YBm
D35jrmpEsSdSmElDucHpuoCR3vaOxV7b3pl+1rofoWYbIgUL+rdumlwlH1vLy5MDw9nsqMD3guo9
idVZrYI18uQYTlRCjadkvBUHLUCebpUdG8LfbU4+krv7P+zbXjsPSpupzkTTgQknk3RfFK5aXlBV
mPMioQfGq2BvaPExgQCnJP9gl+jPm+hfxS6u5jxw3vCWJO3FagJ2wVh9e0P1589M54ZKfEFOrKFg
4dHNMq0znkmedOlAVbJuodtxr4MuTuDpdWprDyC5SxNmA0/4XCKW5MgC/cXd/AF+b91p49garrp/
MP33i9o9uQOpco7Kv3Fj7WalKfCBWf9Ohn+A0Z87AHh5i/+1sY0ILFU1llzNxPSRpvpQrrbMdxlr
XjhQFNb3Y3cczavFizaITsaAeNv2+1s9TeqnGng/9gTYXRqMPdFRbZnN8HZdArmGJX33OHFvBBJO
QBM7OyrT9e/6C2ibWBPE4rOYl/xCYXRZACGV+Q1/T7R5JSS8TXuXwiES5q5IG7JKsAWzcqmcip0C
l81sgeKFaw9Fej7Eywhc7MUEyja1P84+v/5+VGWyi/oyPKc+G8scp75VKoIiOEQpYYnwg3fg8tcz
XLskzBzeTco8jnCi1UF4LWlmGQ2YuelFHLRTGItOb3AJYZnXxIm/JUmco7yODdqH0T+36TO+7qyB
2LSOPkMFfNDfJNzZkdwEQyIytWg/kxdLd1Xkoj3df2q3xreIbgYeWJU/aYYAMt14S/zROLNZ+Hm4
wxiND1PoXAHgNDEIxkdenUOC0aRRgMHR+Y4bqkDQ7DHqiKFQwnSRY2RyhShohAbMR2F7/Zr5L5sl
kS24RQirHQDb4eRGDy4nP/637IzEvIg7inzxMqZeYvSEfekRNCOliGpuYLjGkmltJpFSiH7ENMS4
jwHUOrOry8kOreOV2jSTe3B5sWyRDC2PgIg3F7gWg+EuOnht7+m11G8DLaQn6/DiSMN0ee0eGT89
4AZBWUHjhgsYEeTSVfLsf/N67tk0aZcFSW5PtycTx2dUDwx9PJOO6Pmajf3EY+2bhb2gOytXl4v7
ZaY4bavkPvLYlg73jRf9OcNaWtiTevX1wCzUioMCItyHimGMGN9Z6db4SqzRifPJXbYyRMZWNprM
7plo3pqurVB4kdd7v5vzuMVFAde8kRIGNP5z33/f6BVYc/XPkA0JpcVvwFxSu4gKaeDU9iPltrGC
PvoViX5pmFw6rjo4v9CYS4m5o+EffWdQ1xnC9DBLZwXohSFOvtGVnJ34Ofzm5B68nmM/58oD/MSL
RtWztUW9uDvzwAp/3ETdmDkUw2Uz8mggwhgMBrjLLPcMwokTxCnEL4Yt1SaA/8IOV1OAtqADW6d1
LJF03dwGos58TVT1I28pRGQj2MvYIZN1xGCy9FvT1CoKMglCvXKrQofYm26S0wtCJk3xv2mX+tLN
yTKnjx2ECn4EYBRmcv6euNXPbiu0ejpRNkulKWErRE8Fiq3smM38d7iLZTShSDl+0saUz88Q5e0V
Z+BZ4pxVq2bTR9mU3PtjbbNz1B5YeakfP0cG5r9GtRG6R8NzG/nFb+B5tFoDR8XJ98YoLWpVsOvp
gwQ0KQ+y/1fnP1D4Zt2zsV0l6z5QKbBa1yxUBHg+1yc/HCjCGquqWVFsbNbPmwM22bx7M7m2y9Mn
0xUF6aoqVAtKNOgShBlCIDe9ymZf9B9J+tR8xwvJEjdH2aQlZsDl3ddfiHJkU2CZdFfB9GnAxZcj
CxETZkVjlvBel5bxDwmuZmcKK5VYM2W4s/DSTqeASw9YS47yQsP0eMMnOOUUgbAwDEM5Ox2Aa74f
EElqPn15YVWoKAlX4yCzB0jd/Z4Vlzqmqh6TDUnY/sfYUa2zNkzKybVrA1ES1coWSa+gKaHPlwR+
aZYpq7HYfOihROTe3rmHqszqB6z1ZQvJ/ZUbYFghHgIWd1/jXR9HmW2hr4a6vqDW3rAN47wGJd4B
B+L9zRjiNzg93y8IeuO1fsRNtzisA0+cnL8fCchRYMTCwaQYAnQiaapQ3NsLbqpc+lrBCPGUkYP8
ZY44Sav5oxznwB3KaE1SZD0CEo4lT7widQoi8NCKDizbImt/o9hhdcyrDZnVzgALx15LvBWXxty4
K2Re+4iy9L6KEI2OT+415i2LuLLEJXCkAYGDhgUVZDvs7khGmWm+2yVzLquWIoHBYCBrQKS6y6ly
JLKGuRjXFn01l4ur7yVGE7xl3ke2IAFILFUtmgj1i8zl0Xq6dU57iVlW0eFF134FpoliH7FJTYTr
vYKjtu/8LcDKVDRZT61ElPdwYqzn1GBc08r2hk4jPad4EH+eYmwrjW0kT4kqWlsZRqzDT3YlEfxL
bSRuttSUeuhfF5cnYGrXyPwtHa4hrwhSvQj1HjcPUCauPZgUL4wkxpcxDM+DcH5m5I73vnX47pDL
RfYhajEWIb/QN4gnD6xg7l9F8SssMSclu1Ls+DjrEYx6Qx+fGfkiaPt8lejDJgH3FUAyJiXhoVdM
p0C3GEdb0nleKN8Pd/5MxZ31STklWDfur134wHWzUwYbRrNEMvk6LHJpkkbFcPoX0KEec5Td09mB
1g9UHWqRIF+eLpnNPFh6KxItsn0tFq00wS9qe6St89GQqfjaJj54Bxkvo9CveVmncw9FGUSJoxd3
N8yvVRs+BblMAXZX1bB1sBciLGUd1RKwooGYACmqomLLWZoVQV7NPHlWDYXvLfRKM4GDjXE9kfOY
gUxKVxk7vUR6nEEc/tGk5HD+dj+eRTqpHWkNLrhzroy0BUpoiaVYJTBdosOi8Y8uI8VIlF13L2aH
51fAZjXdIlZCQhKYqpd+CCQ2jEFHhxY1PrtFDr/sml34nHOgioXqcIhXQ6fZwK9Y+OVqKCR4Tfhx
joxx01B9tPVXXvpYx50utnXavbE/EU/sXBy+on7/SuD/c7q4PyVZ/ASkkohoSidHp4JdobrkGaHe
beVy7Br1f9jLVBPUFeJKaTbTH6zGYLLkXRTeSwIlu1igsFkqAPEkl1WHlSEtRYEyxLXHdMkdY36U
PLlvRzRXTrbYB339nxrnIVQlNZ8jTqvtfwpABPJwdmDBEl3yfeDP8nrZMeTSeDKxvdgX6BUpQ8y2
g/tV8YyxCRmC/UJd8Njgjl5dZpOuAEGj1vMA1y85pyfplgaHSV6ASdmfe/laj4Vb6uA+jlbzkYE5
eaUZYWNjVC1J87MsPVZAL67cEocn4T9xZctI7J+9nM8rnt2kOA0mUJPLF9QUm3QMmmolZ2elR227
8H/uqSUztatCpvCdbEbsSuM5CJ2hlM90ZJmYLacf4Qe9+s2zLUBPwQ116xh+Z+V8zzT0cqANlI1+
LzsQFCuT+eS/izmEFxuEHegyHHWoIHgRmcEyiTrnUQbJCVvgj3dA+qK/vIJP21uhTcqy1AU+QdM0
qzYU9fk2pfbI/JFYwQCimLB5Vq7BbSVoKnCd51Ant3/w106vjIFjTTrhWXdcZQXyfL6BLnIdz10P
Y+zIQmTSOZxtapi5bd6NbCX5oiPn6+sP+8ja8BxETWqgfWFw3PZXHlp/EpubTENI24kmDAqobqik
rzWwKT9W2BNVS1rWC6LdRs6GaSXLNpjEJEiEs1MB8Wt4WLvpCH7C8ExXnU2lU6g78JfPWUwCMbJU
fVpov1JrjJ3W+gE7AWe86uGAdQ+rLWppP/ayD4BNcWxUam1o1SXSH/n6IM+cwEecWIASWcqlQx2s
bbzGWhTyPcrU+s1V3MzMcHjePalDtcYm6Lfz4URDleR/1vBuHYgG9AuY7sPd/vpFjHzlRvMxPmYf
aW+BTRrq4IWpwTOoQua9bgrEwia7iSYAND2XL9zQaU0Gq1WL+y4ifXBTOAQXUXDCLY5Z7SDsCa7i
T3X2DhgO4729b2An5nDDnNUlanETNCumQFgMnSISxDN2yL4Jh9nbGR0pyvhNgX6E1VhAXQEVxnxU
EP/mOoiCbag+/zynnGdLH2/IpCV1p/2C0MVEX5aP1Gq92rA9Tuc70DSKi1Ok/o7DX99ngYjGFLPH
40+/FxpjKxfuOnAYp2Ed12lVF6wI4u6o3nAmxHtWnySBLVn9c2AjyIr6QEP06vifQjaDQRUFPY9r
V/WnBY4NJgycgFyHgMCStGJ95dE/BEW03vbaD89ro1hhdAWmUYcJNPFT1JipObVDyMQd4v9KZykQ
V5x5LTlI9hZxSxxXfBcYdGMSy0woT0fd/zO2ailSxIq9/AOa//JM/lBSmvquDzNwgUQp5S8Km6Lc
AkXhh78XyS0iEgdpTYW8B74HsHhDfhAJHaK6HfYgaT/EBpG/I/7NyKDnkgvzZfqwFYCd0JX9zdAx
C4YTq0pxpYELrkFa+eQkcWTOaM11G0hbZY65I1KLofLED1TU8Cmm2j93bNzTdA8bP1po5F60U9z5
uRwlOVirLvvaXYHNoh6sbKczv3nDthm50jp6O/KJZxXX2AJwfAp1bnQcFSUnUlALDENV4TTxIQNH
k5/2Oh2qBiziaZAmBs1dqgRE+6sVB5ulCCqXx01Hk4pwTc5XXaQ+MpOxDnrSqsLJBOst+CnBJawR
YZm1TMNZ6u6Rn2IeQhpvcksxLRPzAaf/uqFK1k4r9k8ZVDc4CfYVMZSBDWxDnRHRgFaXmiNi4XCr
g+ttBSY9x5XA82cULV96EkHYXRzVUoVDsG1Rgiw3UNilFAf8qqGcfZ0ZbYSOM18JDBnCC8AqGBfQ
a2nMuiEnElI9zXjsxWsckEMtUmvCpk0Z8smkZWWmFOJ1Nm77Xl1uIq3pfnkZhwrgoaBZKKtr7v/X
XxomUIH08a4GWHKzRrHo15z+5wGkG6ULO8NgP/KTAhR5yMSCPXAYiLIyPIghgAa2wvHvD6oJRDv/
b/luzRreW/dNzG+cgGxnun20PcjJspMVjrBffzD9eX9D9xbXj8N5dNoXlYdBFdKCrFBXeyNnILus
b2eZauCNduCW8Rgw7yF7B+ZAWGYO5mcbP/vF1w+JwaTf9chHUFKGi8U51FizpQA575m6ArI0eILy
Xs4mXcQo8UA6o9x30TSCos+aoU9bw6qN+xWOIZnpyDd0KHulTv/dATJ8U4BLvbP/4YUJZnm2176Y
mICXAzGHwvZocY11zriCzUb0mhk2syu1V5s+o7yxfgYGiLTjJmPWK0sDbNG0UOText8mGAe6O45L
0m3oZQYxzcfywTtV//8cf5iTzrFFbpy1MudiGqsROTrU6HxCjxyVGlIhj5xxOTfTj6wGY9hE+clS
UNWh249NTbLsJuM3wt36iSy3ZoJlFZwGFviBUSbQRaLUg2UxQHiikf4VziR3SLV7la4HxZfJnzyj
yBU92pKmBFd7viiHmblZKrfK9yZMZZ9bG5RdEv3vhZQz8WVkIkqpyNHwD+JlOi6Vbv9CZiUjnQDa
Evo8AvWFtiUSQIS65WhWmxPQtW0E/iHJci8Ul3IVSgOUyI0vF3RSM4c9WHCHnutBSIYoG5BmhCZC
8GngLxdDS+w53qPK1qjzUuleydsoYPQ33kYfaDfX/PKTKwRCMeytp3w5ZkI9IFBzcm03//eyTwYM
Y5vosFYq3Z8PyioL1DicPMEg0Jk5mMCsBInVJyBufFGJiYPA2Ujbwg8Bwa2zHoBp5qSiUhGjRPBH
ckELKB+yyxAsRSd7VS9+gs8P1gyXBiWhhNDUA8RFc7nAfhtaNgeUP/kXxWZzDrgQ+sbKQDS62ckm
NIJTLiFFbFfq+mHb4Pu6CtQ+xRhD+UKSOBjetZJZ7oes0/tHpftBzzUaPuIOY0JY+2/eVyR9z7CB
p/bufRWXrx3Y886cQYOGs16E4IfuY35xkjslW0WRw5QfvzcZclSFxnwI752lBW7aHnXsxyZIPCjn
eMnOif8sGOJ70EBE8xd5PdTvx7nFHHLDzEjhHCQye0y+MWx8rjNlrL7E4yjRa1xI6a1iGFCgGI5A
6DXmBTfASUvVwVhap3yALVWbn6Mpxz150WvOPGQkt/f/bNtm8KLnzi0NoShk+p0lTLZxK0o8BYGh
ax1E9Yu7k7WERyprYVFchDrNBqf5mARX3QTu0x6QP2UYe9sHj/p+ENzHUsGFJmGTSSJaSE1ZRaBd
fVKfEDpUHY1FokY8F/d1ZGLmXlGzpM/1vwRtv75f7JInMkGO30p7VY6k80PWvBHRoZgvT/a1vwyP
Q+c6zcshT4SODXtN79O0zFEjj582ghp2McXZXgWSjaEpEKDwnEnFpJpSohKDQgVeC17QdcM58hN3
oMGVk1G0ccRNUrsVcassVcn6bcXUCN6w/UXrqxOA0On7ASVg2RlBbaFhtUp7eWz09hcgxDw5Ade0
jcAYM0DXSHecomxLrCe5kbH3fq/uqSIEB2JebkqIn0Ry9RtW2iCf5Fsg7a0Ml7pzIcRQAhKWQR7E
B0cnrEMlYi/nhRwipS63uo7I0Nd1W+ELxX2i+b6jRq60zxMVfE1poKEJiAOHGFJOpKLsACWZjMv9
8cG/20bTBzswdK3Xc28MkQoRROSQgQUopaNuM6KWGMdIAG4WpX5f4TbNCfOCtTZhSHhnYfQt/vNW
WybrNiEUgVt+wrBNhNN57ko7W1N09Zi96JPE/5xpT2VjXj/0YcUxAptMpEBTkgz44azzGKPWSwqD
lx66AcxePWCjMBVEW6+EHzsb14zYGU1mZcrV64ZHBFcslsqAww5sdWnORf8KtNmub/cl/+twc1r1
j3CA5BINVqrZRz3uOdhS9wfTpEXcgfwmW0nMOqgMMLG7PyX7umWC69quWyVtIrWamjbFOkjKCUAs
oDfk2PpU8N/Y3vbYvxGeLnVY7WdKFCybamtLHhXRJH+uaxBe+rbSUoEcPvNtrQPsKh/JKykrPEgm
cMQUswJS3fvJr/r/K/JoDQYXO1rh+xMw4gdAkdB3hPKOnnJZkLJm1XcqMLxa45a/qay0FZhWOTCN
lwggQ3I2JRPoSg1WAE/cssn9GTJ5kq/gqR7rbj4n9ddOCoUeP6n+D3nW2UiKdH3s0DW6sWzSO9ZW
bwp3oqUMZFgw0xTanwLjcqEwP1scsj+CRRmiIW+h4XlD/n0smBV7zUxDlEbFpxoNttx4sKcxVA/m
jjP2+4NET10f7cXvC8FN0duUoLXsNFdF0crNXkPT5NGL9qRGwoAD8g+kQ9NAYBtaVSqAjAfVp5b7
ylwn9WYwEzJZcgWbUnMYCyFlyy4BPFolmIqT4MTUl36AG6ny6yq3/eJI3vUFT7J2IsrE293ZeUY2
uhbSuErGJ6/gDs9uN+WwOguIDCTZqQXjduXL4awXGkZYx14p/1wX830T3JARREjoe57MScwwsD0A
IaTlBT/0ukfFRgKdc9G+xp0WjZh7C25oq+2Q03emtZ5OQZu6y8++2PDPXiOkf6ahbarTFStA8th4
fLmyKvz1BeRqm5RygvHOFedWicjtYubZ1tzM3FDejhIgxUqvqA/UK7kKWwVaoeIrpvQtMeLa9VV1
gLufRJ8mHFGHC8Gg+73pT+2h8DLYt/248K1StgwniKXvTFgR897ZJQTM+pqF6OcE6B9M9EA969o8
ow8z9YvWfwB3+EkWQnTIp/u6ESbEVidFGXLov6Sl5WyeDdZRsmCh87nqpgwkYM3K2jjBpBHRlkQc
UgFPaxbYx//gxNMtdM/0lj3iTnTzpzm6D+1LfHQ8iYOm9sEKaAbvQo30qP4eGDFv99meT2k3At0L
md1Pkk0f725oIwtDOYmyzIgfruTQttlKQtJs9yMKmIPnz7cHOUPc/z8WMRuJUp0ZKZZgDCtT97BG
BQiH+4GeSTtLDUU+U3lNGRSijo+SZ8OJMYJCfvETJMm30AX5zvUlA6n2fGtdd7XIXgI6kzjUT64Z
G/wJi9sWHhJVSx6iwhw+oB82ZNo0PSnJTCoc+TWQWSmfxFNA5lHp9Pq3PXeRv1uTYe5iYsm8bGv8
dBQ59erxyvnRQto8m3bIqz0ksnQyJ4G95U3GCSCRzaUYlR0lL+UTJGPmOFDndzs/NTWMvyOGc6eJ
/jpVWXs6KPR1eWuInvxUjE8FOZK/AlRBRzf5hKzSPAx7D5C1aVUvqpH/3GoM0fJFXtoVlyhsn0fZ
K0ODebEvzAmGUg6ZPRQEzzrONNQSZQ6DwEcSO//zSIWQJ3JUyW+tS7efez+GwvItlMeGkuf8jjym
cX+w2mUQ5tZOyxplO7L7I95FfqUfBePzlcXtFMO5WWmHfxxXv6S/0q1/R1cJWJlZCDbzHlKgjN/i
aLZvS1eLfDne7coHYOneqtHoEQJUCSI2mjQuvZ1e2KnchZ3O/NWkiBLJpf08cPl1HWyXUOe9v+np
45dapt/fbJamZKb8Myz/coj11cchC8u0hs/OJH0drt1ZB1DvQjhTCFVj76nWgQKQMeIVtSWhJSkI
E0HTS1hu7hstQ2vz1URhvqsTilDmENgKaCpERrDdQDoUbfxAxtoOPue87oBlmASGm+eXZYIaDCbj
FbEcsNH2+L8inuu6qWQsHvk9FUJvnpJQKnCE1RIu8L/1NDopf9Drqjt/xodwYx3PzOYXp+y7ZcMM
kBN53j+0BrVF5XrPGVI7YMVOUSjXVdCrEIEc6qom4PMhe2AnTeUmtz2+dF1x5L/HQyPr1azaBVx5
OCFebChYe/7n8gLp2DVoUPaZAKOxu6hbMH4o3w/qlG6us3UD3qFVFVORHTaWaeuKgQFU/bvGWuHj
P7PrVvm4YhaaXZBui7CgaUFCOU7SN1bUTs/xqxCKvUK7aaHi+KBqxyPnabPIEaYb7dBiWzf+eW0W
+KtZGJsCsVwb5Nggi0nm78pGetwiH61fZfW5kBXr1bmArd6YgPjuBTGbcpjutZEWtsK6iFHtQhPo
fiVj5db4ZktYatnr+s0wRsWLBglRv86yfUXIAMFY/s5TRQ77QcuH0kQgiYvbUx5IdynOpXNVzzrx
cQK7h1dAFlxJebQVysb7uzLxPoFN9yL9MAvwjP8hxXqScee2gZHcSA7nfMxsglEzSbEAt8I1oQ5V
4cus1/0xpuJe9ggXbCyjtdq3wu/sg8k/dEWGtbTuORo3lDqXXpmB1YLKtFO2QaUBpJFdd52MCB+U
PWY4Xf27ESGQz7QIxvQDdlLdfayUF2T+Ne4k3VwWkGlQuZ2dDrDVxQZ/8tINzhlfwdlPrysee2+O
YeaqoJrCYiUU0VaiK/+EqynOYHP34PD3FvjtNAxjXTQcomP0iQX81Ez9C8hF9WrzvlHxqYQVLNQP
2HwlYVh7DgMLG3Us09emoyn7bOwRueQT8mQ+xeJK24siS6PIwj65mKtaeLpe9BZ/fmEZfzGRn5N4
dvF6wyw21roPpySso7IlwehfeIIKZxJhW3QV4T1BF6+1yJS+VoCDipWCAnSOH90tFJxO+3YbYELu
F1T3YWXlpniW8OyrCHWxDruvUmmmD5IwyjuM0PWkzjr3NF6y/QNJTEQS37LXph466Q8jM6IpGIg/
cGneLS1b+ON2YxmcazdfOil2KFWWwVpgw3bExVnZLbxT2lr3hPdIvd5jEeqWCA2Zlo3V/3i0CMwH
JlWSaEc0AmDTTocj8KKePdfbiHjM2TMEpmSRh5ppmKVDPmqAkbO9H29UyDFCJZ4BI/QbXkbF7EFh
dmz/bYbl/q8WMt72A1THAVItSTk/eWV9Ltc5mIorkcRqC4IKW3g/fRykhgTpqrnkYcCxwd8nHrNN
iZEmmAaCrx9qkUddE//OFfOmqI+pBxYaBBRclmOyJ7TIuD4d5wbxIqqHZd+1KCPsUS+juBjiWPC2
yG7cmRhy0wBcwjre+Y64YP9KtIP1BgwJXQ8a9QWd4MrTv7kGGUugtlv7IGduWw/rHJbAP+pCm5T+
4q03dmjJHnhlY645cA8uOox5VVcsawwnnKtlkrkh4fKpHGdqHHJonizStySBCwvrGZYiPs6c+glJ
sIizBfTvdaxOMMgX/gSV8o2q8Wt377IxMIlfcZPI4zE9TYMutwCPysvhNmaeLvJpO8yERkjhfh9F
s7q1hD3XXJvBwIxBHrwtaUoYFTKtjQLzVHt/IUhCIp41Y1I/W8bY1WbvBZ1WzqnWEdzdv0b4F9If
MuIK0hw9wfx7dnTJg7KApLOmR55AwqBZpaiLvF25vM10RQFpPll/xhHMFw+cYHO4YZMNgS99xGar
QKvi+7+z19P9iRankTSW6S7Za8oVysG+9yfFKWorhZQBgXl/7KfHEzWF8H/fgslhzXbLlKfgbZqi
D5sxLu7HQwZRlKivGxZxBftegyEzn71hCiNAmdZE/AfPpsAujSLUgI+qRavXhmbw6GXDc5EOYxwg
8Ag9NtuRouRA2k7zau/a0YFb7Vr4V9EkDySO77FYSWGSJKk12cUfjmEQS1MUtHHqxmT+Zvlz7m2T
nIbBoiE36xBqtNK6iLSJfYJrbVJPjpw6XtQ6XYD19HWoPNnHa2FgYIasQ9jHrxi9reuGJKVK4iX6
RwRQCBvGtQAjL7nko+VGk0Fdpjy5tanvU5rggnxEorhMyrYCBZwv0jfimfY3gRE1e9QJNA/eRwlf
CiHVRLE5/c6I+bgqdop/cuzUEBfuM36/CRSdBkFiBbP9fMkMr2HOpCMm5gBVjQnIfXq4UhnVQhvU
wvMyCsr+MrzMvhAnOm1TBw6Dl4kgIiEZOGfrP+FXWyb7ryKRFJx2mYDueccJm3fF92DS7p36c5y5
iZsVeex8SH+MVDstPTLcRpsvyNP52E7q+4iIF5/ejKrAVwnz3Wl7PaRShHTkxeBZli9wQoNTLe7+
m/0oPcb5VSQefkYKb7obHWddaZuZN9dp7CTcv9UfeR+BDLN5tB5YGL/L4TV6PoxxCVFTKkNXQou4
EczHCCR+4ggNKPmN/T5xo2C/U3jzmlKeORmgL+Ai1SOmkhgR5qKOIhsWw7091F6ugrAzwJxpPagO
P/R/YDWO9sK93XrG97j7qQDtkcwoEa+a8nLaCAnAwdzsF/lKwhHBpUkmeoJ+UP1rkbLrbL5Ea0tC
wTu4ROnelEUyn0LUmG7z47wLT1qoyt4/5opfyBpCexDoLx/l90s9wq7JgmsJKLFVWPPCWLwktVMW
A9txWTNln3Mp9GnQrC6OreGfbz5HqGUD/tna+UTzaEOaH/m4HGtt1119VVKm+UTCHnT/TStJjMD9
2LOn46r7qvsizXXHaVffTpIjshE/pF1xl8tlX3ID6cW4TejcHvumkeA84Qq/SKPhzQ1aIenCLNMN
G5h2eW4jNG3vjegLuMoab/2VTboLGF6LJu36tnayxJDTN5iUiDRFpRNb61cGj6KZf6VPOC3y41ef
+8tcIn9J1PUYzb1HNg3fbLLHxjTzHWiw3gxFReCIhE2mklEDa0i9XUHuMJt+TTNP/pgXdZsAZ5Dq
ix5JbmMkXugkABqhz+OiSoEzOv6vwuIQGTGOup9Ts6+PkribuWQy9qcR4u7k2hDnfopyhxgcqRzC
U6emzYFDGRSh7zYmvJRPB2HWm8E8WlabRYUFL2qV7jn9Ur+zyZ9qyjeVAp35BpAVVs5FyfC3meQN
ov2A2z9/N0eIUcHeMKOC6EsFvFfGqw/Oj1qtafW9OIAQQzKWk7aQ4rmoiFrW1t1U9R5A7H4Cm7gJ
R2KeupZzf5sy/FknGOuh9a2r0cs/xy5VPH8RmzfA7VM7YXk1rR1Hmy6FQUhSq15EIftv5gNxF2lL
Ku3GSiddgK59HDuKEjsEcBp1lxixNckrlXZSJoinzvecQhsU4v4Pgiro5kiOcX6YMPZuXFHG1b1Z
Q54ONujs9Ze0qhP4Tr274Vaj0RXybmAeLz48Qi7LZi/IfxLUTCH/wtOIHFJYUuPxIPDRlqK7cuJk
s5MefKIUKv7h1At9oNZmq399gWgMuG15VKjpER6oBwVQsZQz+0YfEltY+5UjhCFiXfa96DE0ty0l
/Eb2PcCBoEGes1gjQ8dmkYQuH4gDhsfgu/0LKmw8EOT1qMvRoaCvMuHGOiUNKpPKwY2l3vQYeWRD
4FosGFoF2HZo/oqFm8eOOrg8sCt5PECTIX6VE4A1UZJtiImyhUiNilbF9khv38bHeJxdj8lVWGdJ
BV3t/uOJfaHgVuhkSVxi1nwwewCZbOKPmB6IlcS+slaQMznXRUwgdGLIV82H8D/DGRahf+HzenMa
9q1ywwK4soz559YolzHRV0Q4U7XEUgccGzve+zeDlhOGilxHM+/UVTXr27RRIYhK13uiDt2qpYHn
imITWUwvjq3951ZuW8OnzsRQCN+H4yYzVknloC4+Ew6S81klXzuGmOO5eLhzNV1s67hv4JqDyS1z
x28+Oa/3NA4sq63pEmMD60ianWSI78TyPp1Vj18uwT9/1Mm6Jvx7FzODTYIRKxYdTnSbsfnv4xXm
Br7JRS4hHUTyooA5vnpQ3RbSAfIeMQP9n7XVW1bXWl3SreGfT4Te0cr5FE5pW/rKb+VNZYQb75Ee
jMaWpDkITq5P9moQjVjB0VBY4H7VEJ8QB5YZa+RkORVNU0LMo9EPJipdui33ywS2q+jdGhXfvAHS
yXPUEjoUwJJuy3AKDU+HbPEZxLLaIDxRaqjok9Bs2KnMiiZwJ0fr4z0aiEyKaNWgipGaRENBSSZZ
pEWfDLkVNw/Sux1HDbDVBiuG7qmudRhXoVFLSTqPMavC6YWhlQchfLutcO8VecsUqOy2TC0hHhf+
i9aPGvDbqe3J8tKxd9CewgMHLzFi/2rrEJqGdvDKHEPHh6y0cB368SgiwzuelFAORt84zvogZCHV
hAi0igGDWnQMl4YxerVC+2maK2laETn50G3XvmupRIH3DzTlS1B94AOlBt53TqK8ogRayJHcws04
wbi3b7X56ow3tp8945Ihee5HSivw/yW89FwKqQ1kAMFVMD4vhdVbrsf3vmz50Or7FCIBsm7g6X0r
nNLEsLZxYoeOajL9KuyVqnOE/8v3/hDRZOdQCuFhsFBinO3/jUw56O5KMXBveiNDP2jZlu4t0X2/
smJEzhe/Bqfw7Vy7BUCNuJDqtgkdHMbcBtDhuEPVaxi7aIKQgxXROALO0etxPpjJlyTo8thulEJC
iu2W5ijttD5zGy1QamTzJhljRjkds5wPHTAjkjTUoTSzr4EOvMuFqRojVkdv2t4AQWeeXRgA+kE3
qjjIcIfGUagmAEBB7fP4KNfjwefTBvGLCaBjm27a2uShOCr6RznuoFK2jl4gWuYzyJh8hNODEuhj
SX6497EMJJp35VZn2wRgCbdne0gOeBcNSMSriVqgr1sS+i8lq1j2Y0t7P68QprJLzkvmQgHca13X
afZwPr12kzV8y1hWgVLO71xzYiccBlWxnJnbW07bApOmqdzizTgidUIsUEnpkin7DkIfprC+cHf4
6F+59jXuTGCHUK7X4/2B0z79etEGn3oUSYQrMV7ce3ICyA3zgl9lp5UUAEtAekOQZcen1lJGdEQO
l120E01dcof3BIYwUoqa3CkixEe7z8iMB4uRuCRMFaIegToLpDPenreZF1MMCxw08JAnXUw62BXT
+3FlnYb1kS4FfjBTRCXuqnDsgFz3+h+RpTS5PEYxmgg5IyQlsV8ExvLddM8anJF+wWBSNwEhpg2a
Dqk7LfskSJ40254Xqx3go0Z146Eg48cKvNRix1akNAa8BMFvxlJL5b7ZUOUuuR4vcA10US1J/4zX
GMnxhG4Yl1ES7SOtlNQQTGMhPrUt3wnQ3/PqUS+4sQa8XyJIP3HoP83fnOA9PbRJAhBLoPc2FT/Z
dCR6EnonwoZ0xNGHRKcWx2zIkOIT67mgSKHXJNah7MAr2ypFyjD3lotun160VuxloK/wvs0uRNLV
3HwoM9+qx05wJc+wHRz7qtcK7q77uoV37fRUFtkGCUO0+FGdpMr9EM+pYa6DGIFZZhqPIzGfCjdc
rTtqbZqTHNjkokxK/QSCzw2yMsSyHhAeurGFuOPFW9Tw+JZKsP+vLea+unjhJEFFAGX5pkdXNbkj
ZL45E2n4yqEvHXaJhQ+2+PGmsncb2HvDc0Me2R+wnlYEAJtQ0AP51lJmtaZzHl6bWAYgTuNfVSTn
yKfLLvLJEua8rIFSPmDC54pvuH7oM3ZVFYIEZRFBhS7KGSbkavPr2GX2uZOX81ReLQ6EwulZxNxP
tZlM3eRPIxXg8wko3z1YcRka+pKfkvzFual5xae/4OVXSnSVDUtvuuUmxT40tefFv9Nb2Ze8Zm14
dZnn0W4nRjr4XwfIBJ+B2d5d8g+S+ShXU4uW/bzXlmjovywashpgYWFYPc+Fe/oAIDQLjpienlnW
m+SIwEHI/nU+AQZjogLD5+RiMFq0CZoEDWPwKtfvyvVd9VfOvUqHGAbt9+2ly4IfIegBKJDwCLFi
sTS2Q7NUI5wNmV6umSdk6KE9pG0ANIbirBesCS2aQtV4u1LncuXdy6d+jYI+nNdCEN+q6ErZRVSw
15bzEOMdGVAkg5KNi+DILNVVkqesoNZkRDU6XnrKfbZH6D7SZAo/dZVO0ptAmJ23EwLFj3lwvmRg
VPe1nllnZh/ijgwzlMxlpOAE6p9BVJn89njPbfAi4aN3iIUb1YwuCKd+5+0GvdvkQf3fS8m6TuD1
NBUW10u7Ch4yk4/er2a/Ia6cBzEY4kf2JThaJGIELDsQzhPHu14aunwOU7T96t9247yY3MWHQB6m
5IVd+kVCj9mOMUZrwCorZuHDUZQ2/CI8Cw3y3luN2D8r0dJXD28nuRfQmeXmg8zTMjWG0GMEv/qj
5y/ex1AeFFPvKmSxS99x/pecVAsMCc3lUV3KG1tdKNt6eTggm0o4fhtrI5Vf5AVvnUgmmP7N8mOu
7v17qvin0lLbP7khrRUDVuUYTVxdA9Pa7fY5AXyiKuMXmOkPgKvMUjiUoOvrYnm87xmW2ZwGWDIw
LA4xxIwe4OtxVJJTd/230lilI7/8+QInDDQUiHYiqDRc5dd3T81KPpGzO6pgy0Xt2101uwgbFQvB
+VtT9gTkLRLUKQmSIjcJJ7fm7aT6naCFV7BMkYgcylnmuPNh8t/f4xnKL1JN2/7uLYq7jHntmNfK
Z9ZALeFDKnHnTctTpRUr0LxlYdpCQExbnVy8e31oxZpJirkuroMXWqiTBC8fHV0rL25Mkb9/o5AX
ZbwLHB9WpsbJB2/SEG2dBjqskHcJycSznDVrmeOzVJ+lqe/CD/6CcGKO1uL4wHDZg+VGuzJfnGbS
vT3a3hHNUsA+Sx6wTwiN9X4bnstxQSHlG1vv9efnyXsCI8PyUZHPoosF1sb1VMDgV1bBOv65jcjr
AmLA58Ghnolo4VFo3Q5cMfPBsSwLEPAq1c1M/WFte/YpCU0JaN3WQnvC8JOOqmkJRxUsWGT12d9u
TicH3cry9V1szQRaMfmb6//EVgokZiUF3ZNeHQhjtm65Qmo3bQJR0o/FRBMn0swSykVk/8sLP7AD
G80uIrpNsQlGQWZ6dxcN4AmhEGBFtE3QWjjod8U3fO1ekMdcHGVm6C8rtsLmnPegpP+Ot+aFWUgw
xFxpPpV95+n93PbTqyfWdELhGv3c9gneEDi9hzNQLNHca5uMQPNiw5cYwgHTV1syqGgRMRILomTf
l5C0y5LADiXQzr4AAM33xqEKG2hT/ec/5yC1S3FRXpnDw84lh68u9TN7FAadkoIg0xg35MouiO46
oOGQbuvhhNS8JdrnpKwgwSLoz3iFG+fEZaY0sDfzZ8gIpxS7Bxa/5vzaMyJc0+4qSut2QzBgWJ09
eQ4r3Cqpu8/pLgFU9lCm1/jl1SCv4U5feU9fQVEs6tkmvnOSi9ij3F4luz/Hf26tfMQVKFq0IOkb
T/JWvCp1Y+O5e6R9UoQ4d8278glz/Xty88ghfxCQ/u99YiUrZJkOvtO9e/CM6TjVVLdHe8OC3TuY
ib/EBso12JckpvhReys6HwnQ9K5xKM3zoA8/cs666gZZoEZVjF8xebGR8qHRbtnCah5hhWmuiDUM
QTyl4V3qnm5Wl5tIZefJbwVkT1W9xF+7lttxSgWQZNGJuqgIY//KTf3q0JUwzHMizId8IrpYeMhy
OqjjBu5PZz6wwYZaF3X/+daeCL41y4JTK8azXVl/QZo6Uijic0xSDccJAN+c7VfV8nmsuIctqqvA
Jd4NfQwByXrkKtFjZLogT+/3vcEtWfxOk6kfpkCf7SzuMRcQnVJ3qARgtdD53oPkZXh7dPz/ibYd
EZw6EzFXiAtXuxrmGNtDxQTYP9CP6DsjS7TPB9X2JRpiY9C1LzaC8Ki1njJuTdOhU57tXfsH4+ZH
HqzubE+kZ/Ih17nPLc03GVjRwPOuAY1A+L40FnEqMNpDta3V2pAXLw6tftus3ofzYYMO7qEzaqYi
PhEcaAXjenjzg2e6iaCJ0KGogcxxNnKsAZExChZOlvWlA9kdNM2N4aPqRCZXte5MhsCrh3uMsbci
I7FzO6Qk3YBlbr/1mIikCruxCqMt6M0ulu7V2ld7bI8RyGI4MitW2+HhOI4jZ1xSzuZp1E7D1PHp
BE7bf4ke0oS5Pxdc8eN3THybh1USixc1vN5puFCji6LUyfUp6a8l+A0Wy+b1LzIUZXht1l8mT7/m
q7GGUo6sjguUWX/IFAR7Zf+zSJkn+1HFnpzVjbp18LD+4ex+3axZ2ZtOd2GkR0QSIPTNoEKQ3GhP
MPQoUGk9WlJVszyPo1BFNS7s1FoG6p/sUUS1VHLI2HC7O35tAhwaUtb+9iAoEPC+OY/McCoLB7vy
nFdSgiq/epZ1Q/xN13TAHrEl3f9xjwSmCp7JIWbjUfyn2pCakeAio+ZiZzzsGwI0b3rIuyWGGfWR
teV0YOzzKNj6XezoEJHu6Z8cxVQSlxXTUWFEsMqaYXBg0PfL/9ZS9xW8HffOCqAs4x8iVfd1/omv
maLB6U0KaZytuJbPuKOz7XMioahGIm4i6d4u9tnsp6DCSlC6uzLKh6Ekq4AJ9SafBnEVzbEic8zJ
eeJ0ZxX1NfiB0atS6pIzh7/79Z9uojq88XI/jIX92W6j4XU6S+euL1gBYpQ7fmp95r7fDGEryzKg
DTL6brxHUGRyBFMhnZU+MzDq2uWyuCm0Uv3OM1mBFzauCsiPwgRmAoS4lR22F/3mDiSQ92uRI7VZ
CvS9vTDR6XoMj59n0ktDDcHphMWbNrpGpu9PWMvB5EbUUj0xh/oLgnTex4jNDOV+1Nexw+T1MvFR
S6cDIYBlMpMojJ8vYalq5z3X2PYFGcu8W21f+0jShKQoWQpYVFVzoWYYG2j46wIVjhZssYl6ESM1
XJg55I9C5ESx0SIfm9L5+/ipUOc+Ic2m2B5Ry6HkgyrwN1ocypfRxCM39CameIzBB49437JEsLt+
mklr6W1BO6vwItWp+Kpe8fc7c7YwV74f+h8AAZIG8eHI+rucDhOt/GH91pNLx/JRNco3ExXPvrpT
X+wt7SXx8KtipBjOw5SvJnWEJHUTtBC/BB0pQ65wijE36/VnkVvWyZee4hgc9x3P5Gvl7v7WClU3
dPFqQmqSUE5AnL7yWRHbv9YjhVnMKSsOU4fcwnQYFOofKWvcZ9Nx3m37gM0Wy4q8vrP3XAvWY1oM
46lWXDkb7aOc8oshnTtZQjuRcrhkUXRUU6naaqNOuL0YqHcYHqeLL6JDAPo68KETwaIz6W04RiWP
x7yXBz18+FLg4mLDG4f0pVC0fkrxLyVqPzX7BpkmG3nE4mGQE9jvd1SxwqMYCstl3HCC4Iuls4md
KTJ9ort9XcfCeqQVEnS+LdKT9BvudygwrHtfeURl0CzI9k3u5vf+mu4ptb7AQsGBa8OYMIBO83Lu
VJOZR6NoBcn1Kv6aEXe2csVvvAl8PjSWone8CNAq8dUnWKd7F/oUUtbj4UH3X6/Jhbb+RyUcF39z
muQvMT/mfhGDyywPXR2c6CpRDQEPVzoOfMUpys7CQUqtt7RIU7nZOMRaCBJbkgYDWbSC6Z6MDDUN
/QB1Pksq51MS9CXQLvpnpb3zuAUmg3SlShSsNoV27i4LFQPLsIMDusIEEXTdjQMgIMIyH2UxgMnH
HtfbUdCiqFjlItEIFhdowVfR5vUqbLO4v6WC7t1TF4fIaFtzonmJXEQ7EwMiyJEXrjjo6wlJ98h3
URDTGZEGkBzZbIiEbFJ776ZvqnaI0UVRwx8L2y0prYC2eP9YuJJMQe37RiT9gmK/hyttPxiYdt0F
fAdHySW8CgVP/PHFRomae+ntOxiCKPSSx3rfQb9cBtqI5Vyu8VgQbzv3Eou3E06x9z62l1Rf0TqH
Lw+EzqrLsa6l/9g7D0wTkt2mXEsdECyFbIxMq2XBQwmnu6zVqMz1F0Ow3Weyq723furIn+zpPdMh
toIxgMdDC3MIxWSomOXWKwjdwOLStnHCvHTQQT20dsYm8iX13ZWZqzW+cYQT2IMjh+zweK/fBLMW
179885Ve1iVcZ41RIifxQGSAEoa9WBlePxDvos+1rzZtaqF2J6ekN/655CKVz5hW0sU72G3KL+Kw
pIOWao+chDPWHQUGND09W+loaRExXwFqHq1hNuVZr+x2Ld8fM+7hFk0wGHG3HL9aHcRIUSmjrFdw
2rT/xD77TvAvb4UEGkg60eO1iP7/PFFyFebDBmMTpaWMFWQlFpBhSfZspj4qy4xXdocexUAk/tkl
xxyCShlh7byw2JzlXQvROudOj27Qb1UkU2HWz9eGVwp4thC7gWuIUK6eoJVFmgQxT3ea2qUD1o2w
Xg4o+3G3hr6BNW9+sdWaKpQUGxXH/AMHYgQjoNUMclH73w/gpjJXksaUMogpc3kWJBe0Us5aceli
GWDmbShqTXU5k6nQa78oCq24ykBblIQ1KCDODm53S2Xc8BZeol1GRogSNuS5NkZiyiJgQ+lZ0klN
z2f5AOZ8rvACCezMPB/HqwLBJ8HIc7v8yFXKonq2YR8Hh27Gvj2rGx2sgQH9TPEsXGGXNBajx/vx
UaN0S2jvS7hdGKSjOgVeHT4zP7AeJ919rIygNoG6gv/s0PhYF3J8+jxTVJHAbQqRkleo8BO1L5OA
TzQSXqrO8RK4frX63Zr67TOfzSJnszzJ4+aF6aHp6M6zNNg74Qbh/JgAMQSIJHlQ4iaZXYxalcQQ
z7xmM3+1urR7u8K+d4vRZsYukppN0L91GujJnVomPjQebYX05vQ7uC6pyXn0udQnNaQf6KkPaDGn
OWSQuo5g+Ln1Q9T+6CyJUhBjWxB/7VWdJa1sokvI45oDbtB8N5wvJIwZWu8kQa2daFmooh+duIPw
QdbkbP9S3oDnMbghDIDK//mUSD4MHqEagfSrkVSgJFVEg/6rAwultBZe07UUQBKyFjw2m2kJh8re
kzEIdZgYCGdtnpFW04Z9FtiCLwREcgxSpzOAUAkuchsJdyJ4+Qn0JmC1rN/PFNhflWl0FbvHzlhQ
lD60qD0JQVhFXx/N9EymoSLp2a0oTccccGmtiK3Lenniosy6qzX8/CAgYjNVX/L6Y+reMlCpBmuc
rhp7q7V61aFURhc54ZxDMn/Jsn7k/MKu9DeekOq4UQGnh6XcqSzHIHESRo7lnq4MmZmCNyZg6gvg
dJIu/CnviDXw/lBvjuh9j+rDFnpxq1SPzJAZB9Ae0N20NbEgM14kOiRoi6OHw135MtiWMXhFvL9j
n9ifS18j46wDX82iZSCrIsu9GtV706425he8g/7nf4VBUVm1emeNt+JJ0ROsPOvZ2pXnernjanmx
CyyHZJ9X50HQRbe7pE5JsiJs4gGNyyVIwIyPgumf83Eeqgf7iXjwmuot86fju3serggKlCMQWhqr
1JEH89Ns8Osrob8znHc/VPKRcd1bcySg/rffTUykawsRGKCTpkcRUUQzAa/MG+RpuGahhK4OxAUM
wjLbOh/xbTwKLoBBLigKH9H40XC3OTs0gbt9VB0UmMwr3oGM5NHtol6bXy0uBcpO4RWgMTYYxoax
TV23AOVaBZzleX5byGU+hMzYVP85OTL2O3YZqa3mV2cu916thyRT8m8KjWxXCbfr4bMwbW+29vk8
J1ssq09oEQYTiFYtIpi97vx077G9GnB5W5guvSgt/tY7tHp/0UAMtB18lz6h3PwIyKv6iiWGzaei
ZLakPkZZZAN+yT8Zmr+yCH3wVGdChkvNlHZch3/X2W5CWTao600SF6aQgbAd0Ay9Q74D/up+72fC
tyjX/ICwu1j8u7bq3Wbfz86fKfPJSoqF/my0kafPFGSE/OYEaj7Byx0xTCK2kdsY3U5ejWV8hFyA
tvzBYCrStmL+RgXZ/PYjWQiaVaI8ARmF4wm8/LcA6H8ho8s7EiOk3U031RN9cjH7dVo384jMlgqx
0CGsehtS0aqiLQN23rF6Qp2/rCxfhbmaknocCC8YQNd+vs8sfNcjCtYI0pM35OhYne8mSlqy6fjm
IUElwYvAYhBXtEIuOsWvLNGbuePyFP1pEbJXCLE3YnthqFDYPXXuHBbpPDOr3jn5ChHppovJaHJ4
3I5oVScQM0/2dIi5o+rJeXebNB+JEm1uzL4cXhRUM2vj6db4T3SyqjEIrAHOdjlT8O9yVeJs4TLG
klBAz4DTLCkIBuDgjxYfv5jwHPhQILXiRw2MOLX6l/beC0uyvA//O5GdgpER9JEzPii0rtN4w3Fy
UhXZj9ztb8wWoNQWF/9C6PcpjeqRZpdado+NXOPIVt6Uufytsa7WXILNw/k/20/+/weE6cvzVmt7
v7sZ4B1rDmuG+Z7EucUDEfho2Bq+AVzUenONCzp5y6/VDa3Wf1ajPi6lA4MM3mf2xQRtE/1Jg3y8
SNOmGpIqoOCdVIoM1j3yBYqRE8zOPhvKSfHyNg5Q+vnCrV/6nm50MDVziggRjtdLYV3iWdySX1FU
sQjhq0aZFRnl2F0+BpPNo3AJtzFzuZhxxR7Dz9gntsg/iPdX0/NUg1GiAD672J37DXlxbf/CQjba
ZBKXAy9QD8BJfvx34xc1nB2Pgjh8Zm80wjAXjG9O+OGjZlfkWnA/YT1L8cuP7Swoxx2aHsToJYAt
YmXMSmWYBzvOxi/n6jWmyaQuQQ5gW+5qBL8A0N93kPHMZO0agVryiE9Kvd5d0vi4eTTbNQl39C0p
cShW4dbSii61CBIzxCoxyPbVCN/V2s6aLakvECnrcMne7+MBrfcmzUtvXS0iwoA6wFpjlqRuCvMi
Sh9FTlVVF/p1Kx4Os/h1xiCrqieyf3hXLATpW7vGib2aQOJHZZHeRKs9tNoLe2MW/n7Hyj374Fpo
nMEvD6cnr90ayd4i/rTijoazRSKkxWdNVCpmJlrpAhlhDTAxIrz8jOrDV/AQobp4oX3Ia+zniMl+
UWB9mNFaMRZbKZ+E6/cc0IYpDtC7kONSh/4JWpi80I5uobpiTst2sirPrDynd3BwodP9Y0BMkBPp
7iR5Q+2N1QUn5SbtTOV5Fvmgw5Aoavj46PsgftZu7XeIvcZ7Gmg/HpPZlPlb+57bDN7KzeCXO5yW
IcfSBUIledP51Qkf9zOeH3N5rtgov3QlY3upE6OR6SyRnMnDNv1/YRUNRFxu1qvcDPVEBMDLa9SC
kf4MzFua1M5p3WJp1PzJihDTSHm1iKQKfKIMYfToaJnvrHIxlLhz+vHYaM9+HflM9fEoCkChp5ZB
vDPlXqwSs5bL/Mp4L2WXv7pm5rddpRatl9n6bOX9PQg13iTVxJ3Y4mUwKpHn4q/ZYeKIQuTrXRUN
ToV7YNX/0e+yyj/8yGC/ujHxP46L+XHK5MubZPtxAfQtuZgKdnJtOKiHDqMLdTW0pqWm42povzEO
k/PTIhiE2LWo92sQIMXRn33Dr1FDYiDsK2rDhoiQ533Rpb8z9Vql9xsblhAaA/TJMw0oGUdsPPnP
4c7dR7ctmAeCJeF/3oE02eVOQYJX5TkVT9eSj1u7LINDHzZmn9c22fD+G6KauUkIhWEpefE17QGL
pbT45ukwYZ1Ku9pur7jWu92wHnm54PFI4sdf3P2O6gKbDExYL+JO+QpbUsCYd6KYbtR05W/d4Ssa
VH4ZR1rlNgxvCm0VOxjI3E01pDczNvbOomWMj71no+1h1afg/XOncrSReBZf9uexKo7jV/eZAqvz
0XS2aPFbRYf7izRXA7B7MnH9WNgUm7kJAh2CVPHY5bo8/1+kbi44xCcleG/fZ+wi2kWhpjhP86iy
36M5kshz9jESuy8pnCDqo8E4dTtNysCG5/VaIGplOX9A+m2EgGcqAmzkcUZUdaNmbcKdTNOqI36B
YIFMLNs/NwgKFnqSOqUe9JTP5ADK6agcYCOdig2veWMdhkxSI1vQ3oPAQ+0gUxvF8DaJyP4jIPo6
tzYZgZT6ynWv2gqwEOjKxxRaNBp4i2PhZ447T17+4xCy4JAZJdKdEzO+ZKkpjSqfaaCWzCS1J0AC
7fxdzDUgMZ1hhFvCOhPPyK6e2Sd5euLc3ZodeW48LO7rzZhcap4ZfbOXz44d34U5kuoPyoljY4Ds
m3+3RVhDK5Qeq/EXRBKzHS/S0R5sEMb10NYGEuCGkHqvfb896xs+dRZYzVyrdW58/NqYkRio5+fD
lcn0V+euk3FOpFDgX8MfDSIDQTV4EtX7mF4v82sGFv6cG13e/LEKVhHLduPVYgaRKfnskxt8f7eH
dPOiId9Hnwd/unAPRMOQEJU3jha/5HO8oTy77/OlxARGLl248pYj0lg3On7probHgTqqxgILtOVs
h3YOlC45SqmR7db6rx/oiEsxos/n5bUB7OS0oCe5oNA7GNfD2x2r5MXa1AkaIwFXQnuWmzcUwP21
HfpKAHR6DjVnecRPj+WUzfkQ9P8KI26yy8wfM43GlpHKpm4jtA+0hIdiT0vC/Vw2BWN2TC659SDT
8zcYKnFa896ZUHFcPng/5LJjY/XYE+M3BAkMNtRy3e0ehe09d2IA5IWumVIwFvGLe5SE6LqLcktU
oa+0KQLnVFHOkUb3nBbAXbNGZCHm+iT6wYE2aZDvukrVARmDgE/q0YoC5qxpiBb5O2OYbfhMjLNi
350jl3sr0uWAfInV/jr75BSTHfcyWokPfTSF//nnxnUn4m4stCrBTxX28BDifO22MWtaJlrzjmhk
IRk71tDYD8onwzmaDN/OtuIwzYvdwdTAHsm9TVF3xnpBmuEHOwNHexZx+bYW5brxXFfOsBJa3GBP
KijA+VmmXl8t+L6zLtgtJrTc/RCMtvqUF+99pMugcHZA5XO9HX1jjed7q6TQkqa2HMRHnv6eX2pX
Bkj3/pgXwDtVwLO+MSMMTCpWJYLBJh81sC6DB6JbnmaefnUKpmL1YzEHuFuHqw+a3hFF9jHPdwmi
5m6jofHli8/nzN53D7TJIKYib00MpncF9257X2DMjnPD9XksnfgzEHEK95YHwmP5bBYXmSguO8Jf
Rnp882VnrfCT4poQ8ExkMJwBr9Mri1FU0+dSDeEn6OnK1rpCb0fcc/UelR3Z4Cj9gl1KbuHqLiEV
NEJP+0SLfFDU+JtVPJ16i0rt33fTT4pEM7Ex8LjM35+kLmz/pAvWvN8SeSK30ni3beQG9fkryVhT
WegxxSTafPewW+rCCpn4CyMpLZVRvSdX1IGIrg6bbLn7t9dxkVGpcgp6XkBgbeaH5LkoHm/IKvPG
kO9+19kglJzvXGYVXyrD+Qp01cqCsIiMBr9B7DpI/WCw2O8F5L/sn1fYEeTfnZzbq4choG+a1sh+
WE1z7mWuMR3/sceGLC14oBCCH8fXYljsIpDE0r2ZIqLzRxVhWgnwZAc4I07RxIB2UDSMjlnpJfyo
cV8J+irCwry+TjusygR2Gbs+vduekDwPZMF2hT5O70w6V/g0YWAC87kHlEWl1wTHOSRZohT4vVEN
oM2JarXK9WR+R4DR6ECtsTdAd1/YWVkST2c1evKByBKpVOVBSZLu/5HC0He+G1AdKIFR7YIJTpc/
ELN89voVxPtCaVtxh2PCUJFfoQ+I5gUZc8+rFY7auZpa9uFFP2VV+YO+NxkpmlL23ojs9JtIcdbG
A70sY1oZQNBjQgrX68y9MZ+2YBV3tXIIdNnExuubjt5yYBq6MreE+Q46uZEcjUBk0RO+6i28bQWp
bLl/4Sg5P5PKQ7kqCPrcbLrEUeMq+tdeH/BIDeb2HG0JbNMjhY1gJ4n8qfclVmjnf5c9eyRAur5W
031SrhzoMpPuxM2uyNIHEguO8mHMOD79WH2qVf3se3SuN2B7Qamll3LcP8m3Ug5Et8UmcCFNZjjx
YiKSx0TQGAfijJYYGcJqHrWc9GfLH6cJe2ijjB4ZGMVzVNDbJrUWmnI/8isyYsC9NJpWbna4YMBU
AKmoyBQq7X98kVfqykIoguet+kwXVKWBe0OnXYWbKIPvQdUNyP7WVK+OPRc1yNuI9Ep3GDmrH3xr
iPTk80QXLd43o5ECS1bsdUaL4Gm3CQ6H+K4j8SYJ18evzOmxfOFTQxyhEYk6fhAx1VJ46+kY0ojB
zyHH+enuIujzawMFxq1RPYY4Nax3oYGi6YUSRJTLdCfe+OKQct+cku1Gzhrb7liKgaDg3K6969ML
U4enoINSyT7+koZPSFserVo9W4+ZQm0eLhrwl16b2oxEVW5OBN9jGLEtWU5frpFnn/fQmGGiyook
pTmq7Zjwt90985JREKqiay+iaJYE+FZbcODsEubuxsVi/sBFlwlKeXJ3WK0jrDND2YPaMb42A1y4
TYe6G7vgeFAjJihxWHRHMacb6HFYQEiJcvT9SZ1ckkZAFGD8yXnU1doMtTg9e+bPSfdOvz2gNRRs
oVN/xgsm4tfOkmnCHGLHrYPwUkqcCJTL046UqVK3edrqcJnz6eYZ57otE0UUyG10qOF9QsXAHJBj
uUeoQfhr+gVTz/KLLU5PVk3ANqggcfH0++4NOKbwON4bCFgJS9xZlpBKGbp7SQpVP/Ujwzc3N5Hk
s+v5ts9Wuqevrm1Ufc9Kj8XQmc6l/lHNctjYM82OFYIKCgoSsm849HktLFFQg9wMiN76zLPtc+6F
kj3urSyTABwri8bNefyvXFLPsBPcyzgjoXzcIIisekhUpaqRc8IApdVxVKlO1Ite3AEequYz5Hcc
PLzsnA3w3ZwE7JODdElNNbu7T7uI8dtBT95OLfXsWWrwKuS1ahm3cu4dgLSqzNDG3E1AvNm78j1L
1IXWBNZgytIUYesGp06883A0xZrnMuZMyC3p1R9W8SJ9PDjvdXsQKFJbR1vYEDC/QNp8poK4r+KD
z1Rav+Muv1NqfIZaUCMcnJhHarmhRB2qKnUN+sJvbXOEGrs0F6OxU/CnqlRtP54rCUKPYbZytrDS
jWiIEndPyjH93RGedoQq6k0tvZCFFqwitmBQosYGLJ4fprlsmzhekSsLdyarxRNEqv1fGwQoDPUq
CTXq5jZqf9GCeLM28N91ZBabzaAnRvYUPHZKsAzJJ2IKGrohRyT7vGiDIqkf7uqp9D6DdNuUHC6Y
tjEIE6kyvtpCduV41IezNBqfvURm9we7NLGrV/PEaKbRHywmWP60CwNeXMlfJiZsAlGMVTN1Q9Ft
aAjYobpH8qMGtE1oouCXuidkd4ezRAc/3feI69ukMA60oBbWBjkPQpqCZGrXzaSENzVA6kyR+GYB
SL7VLYUfB5CNyajW/JJ9vp3PGZzgpRVFek32mSRYypER/lQYnFFisxQVdjvXz8oubcdMQzgzDGGN
IQaWvXcL4H5Mxp4D450h9wFLBwBFwg+4/CrIwc4kwLcWD/VfLP6ZWHKJhx+WaLAe5ayw9/VhHf57
58A9Sq2w1ueXbWohsQ19N0guiETxCWHc3/z3yecbVA9QgJWNpqGmXOj3Ua6SQavMWWZCMYls2TLM
8JN9cn+h4pSxdXglPMKOmAX2RJhsHI7WStMuUQckVhueAbfDym8fjbby6qb+u/a+RLijK0KP4SiA
l1yMYBnqGRC8/2y5NAXdkSDGSAzyLjhuPrPylIXNPmPP+iw68jAi7KRRJ4ZQsn6pPthJmHhr6RiS
UTlq2tUYO0WGotk2oxZBGczR/6bjFMPLmGPo+BTFjavcw0MKgBDS9fomsdLg4wKQtXIlFDVvm8m1
Gzw5zWkqmF/tD1WlIWR21z5QwTW0eyoZ6TUX4amw4EzfeSJiDsRYNarpfoY1rpT3qu3zUF2wtJBh
iKiiLl3rMADGX4oLeO0sPJECmow0od/PKgvGLG91gklq5nZ1ZC4bmgmhu1NBRkBDGWnZt8QsDnAk
s7qLKQWJTqK3BPcHt1P9guXoSmCocovpjUBz2XgrLJWiVAvcn9ifQLz1p1p8r/MUU09YEJfLKTER
VEb4k+NbWpYyLt/Twxz4e4NP06JXIVFdZcO6JCEia5jdpQkEoJLYD8nAUMrid0vuhmmr+h2QtppE
GSf6OLxEqus43/7fbA1x9cgdU4Ki2P0eocNW+aeTanrX0kHJ0Ai+gzJX9PiV/KxA9q+CGTuIOvyK
woihe2cZjPvL4mPjXaBaDgjHl9bEWAH2inhfX0Qz/iKEM23ipdnbwhUV+H6zRAWCtNkCwe+7p4f0
jAtF6E7P3bLC8HJs/TlQxWopa3MSbII3WPUdBr94vKrlImmHjkGzrFbyVcxm4R1lSrvz0/E9wTVQ
ErLTAb4isblgMZvRpKJ8yNej9WeHzNEYEpNgYkcWDyCJXKWwT++n/BTlAnBdqfUFSasGrJNNli+T
HCT43S9bSdkD/PnIj4D+8P2RqJlRgHdNM5CtjrbTTOGByrZcgWJt1lXoUxOeQ97VPp2xREa0Ur2y
/74iby16Hc+UdJZMy3UVlSBJNHTtWv/pANzrRpN/6oZdlXHe2jSpHyZ2PxrnsvmLFN2niDIsAL4J
+/0R4vYwBwquLpXfJhV30mYRJeF6jR64foXfOymaxk89Y91Blzj0bWxcBeT/596eAfdzylxZZfWF
EVkJW4ZcBES8eG1AEEmiKysC+b++qe1imqSDpFjPFe2kOArTcHBEVrMeDMo49iZE+3V7mnHkh6YE
GTe7NooDYPxF7t3blLGDf8sFn/0BxEN1mutD1J4OCT6lWyQMshQUnF+l8IlrXHjKGEBRBxgC/l76
Np2TkOA+NeawLc5zFcNxgP6qv1dU0FYLQlCToVZYYSVXbB81Q/lEm1RytuIQY6yUEzVq2u7BJ5qg
Gn2Fsuq1MZYcQfIurZhqdTJpSVqiq83/f/a+qRZddJg92BzT432JgvnmbuYQGJSxZDhJWhKVQ4JZ
HBYmlOspDw1AeJakrtH6MZxpYe6MMEmFErVfnfxq7YmLT+uunLFWHP+3q0UGth2sD1X5VfftoY+x
0piJ/xQ2y6XdeBt5TB8LUSjYodRPVnoV5tL/LyzRDDbQOU06T+rGri0L5gcuWVKl1YeBruKAicC8
VXCy8H+6oRZjUceKWHd3pieUrpOrVMv5F6SRk4pEKeIOfRJ5JQsDefUhep8OMpIrF4EF13CnITuR
n3AchcNFtEzQg/nvxu1Icben8TfyuqFYzjFdXl9LyWAftvKJTPsjcZQ3WLVuKpYJ5v8n9r27vnBL
Um0XjTRxB4L4e2TG8rIls6mvZavrKvTo/XLVcO40E6m6sPxROO10FGOKTYVlKWYu0YHcWY4d9Gct
GaDQm1SPoukgBW8RiECOuvPKgl8Xbq+9nXHparPMhFqp432dRTMlcfEhBWJxGyW9U6DZaM7t10RW
NEO5kdn9i96eurFjeR029RI66H67dj0HLgAcqx49hz3He2a+a/hllm/JWK0ktPZF20+nSsNXnJtN
PRyzZSt98ILATMta4+kWodYAz1Ead6g3egxvcMeDShS55+5C81j5jNSBHyzx/KDGUt06AdCohYLc
ofpY+4ufbizFKbnd7D8FI53KG4JsyWtXIE+yhKpe0Kf5wSqUdFV3J4sCKrzEizPyQiVygaXzOu5x
buR+yUzQE0GL6Wkahl8r9yfYEModNgScXDp5Q/KthC6eu50qNnhIzy62OfQqj/HlchUs/TIjarjt
Q6xfT6+SPgwDVoL/gOkAy7OJqxXLgwCudYFx4On2G95jQWlWJZSbyUQl8Ku0cviAfYWJInsUFeKB
ySbDOK8N8W3+Ty7CfXRF7v0u/9JA++uz3E7CJKrdH5K7r2DiZDkOPMl6gufeMzKVWCvlNhcpfet9
eeE/j0WFkl7FkyFpH/B/noMCEqLWfXalvugPPcndBfOerA40Ro5v6fYbrmfgFFZk/9pf9uwl05VK
2fQb2aaPfpvwLr1f/ISCE/0WLGuw6co1elqUV/FBw1PJ2iCWYKxGKxoOT0Kgf7mu62UAJwTwHBGp
8I9Gv8+QuHznGr+hUZgGIUjNdjOvlsX3Lolj7JKbR6tja6qL0IzxtEcLDEayJmUWQtItfzb+ikxs
2BQOMHCz0ra6kS4nYu/aToySEgf8ij1egq6z1p4G2JMaVDrKwxNXm9e+q2kN3V00YGWRRNag9b5x
9Dzf1YXEMKLeUzDRYn0cfj7U0mpCH0ZEOh9MFvInS8y8eImz8gdGm0Gb0xwfTlfJ3uxeqdW8B8uW
Tn7qfXuXxKyAh6G9aFy4tAUWFcQaTj6ObXy3xJt60zXR70kXLR3wD0O8DwUokZHft/Z8w+QKSFg3
NncQvJrQB/X0bIEe5KijY9CCEpxrEizxTNPYaiVnVhYwlFnWwHGDSiCjHZ2Db7I4EnQ8NxXFJwvz
UJ2OScrRdpSG2SRC/1PsixardXBcVjJSOen5SqildvdABhpsF3KdtnGizhzKk8fzlysy0rClQBlw
KZjbV1nnwxxXqzuRpxW4ka93aC8PhZqxJIqn7rKyUGxNSjmy61IGfqJk2qQf6d8azbrQZDLnpk11
3EwaStGzf1zBscgYYGpplZ6gLvlwdtkHEO1up6iEv2KOfsBIQVDqjfNv4AVAblWc+Vssq3qk2od6
74D5hMK6WxJSLkHMgh9h51iJvBYpXR4aiMQC7h6g67KHHlgScU4ASSvvQL9bv3kYmzxAKwvzFbMF
TOpQxTfVhbkucglVbmuMKHWTgyOBpM3ze9YYlmXG6T1x4EdCl8DVAwVZaGRyZePxdJTXsz7N8k18
QrQN/QBnDGssmsVdCVwn7MF3KpizGONXauPiCfDjI283RHhuYLTki50fYMykX23XlRgaY+nxxv/n
/0nCi5jyQqytK/sZVrLnFPP5+JGdjQkZ3vPUHBePuC8Fr2PW6qLLjB9q+2olNSHMFM9Xuepgone+
7eldLlffoGKO4+aGsHyZUEwc+qsyWR0ml9BFEVw1LFpHG7El55mKBvorJxyrKgrGtdVQ5CCNvJDp
Zxd2Pog0ClOwai0EniMYta+30pQeOJumANPHtY7V8sYqOVKcF0jsdlVsRANbgbVWNQ4a06ibQp6K
C+WmpXOEvjL0i7C9Ubfn3RjuTij4TVfbZklB+jP66VFldXcTo5EzA0L91wkA8VRtrZbQ1N+ALQvV
ETzrB35Sc5y3tK/6CpN0RuWscYxghfxsbTW3Jydvc9BQZL0zXLazADFNhAtsRERmjGhm3ZOlED/6
TaWjYMSW7KkVuPp47rxgj6C2b15W8cwHbFzsiZudmwhRbq1bXFkkYcMstcoPuELjgP+LVoq47l6i
9C+v2LR5YbSlQOmLXfXa+EcINhuVpRvAlMyZq6eNCKrGdqsbzaKvLICFrbRwTrMLFa1/PK7Meuhc
40C6ODRb9iRYjld21ztk46HMAp1zFPAAqxFgf++Olv8biiDTVPxIduzbjnr66mnldtNz2M2JwUoS
OcFRDxPX95/0RDaa21o1MU42P6ffZ5fUzpEk8ZugTxpBe5FGvKiwx6FKBV/ErS7KZjPjQpDz9PSM
WOmtW/e31VDL4LKx4Pr08GUpAUsQWHxREa74MYUOiwAjF5tJ6qE+6dtU9TkKRHNlVXrc+gBBkxzT
5TTd4eCrQ1XD1YzmWR2WzMzA5Psj/Nc8CwDeVrMNC9/yWMbGQ7vom2CDO7mJfFiaex+tHlEMPhKE
zWgQI4qrfwQOzErFWqY38rOwlz9V7VS4mqqZQn59WWIfkEYU5r+4mU+OTpGe2P69VE8donTStmL9
0r5wp2fqaPnDsWUOJzkfgR58goPhrRU6rP0d8yqhxHADNEqeezsh5MEHDL/T88e79o+AMTkaTwHq
GoFfMbKgoUttwjDgTD107abEz5O4334xcpCIZf51CgJLW5I4/kWN5PdtNQIlTz07A+QfbyxVSDeQ
1PEmnFlGIPNbKHQ5AXrloP9I9N8oHTghq6Nk/VSk5jUVpWWz7+2Kj8CC+87VqGvo8xztO7YQeca3
4kfFj3cKL83wQnCXYy2a185tQy+LvGqagIDD9gArXGXhdK6QC1v01afcr2c17Es7q1SmxoXIXCLi
afBBkzA+49l2vYhzCMf0xX9vejKqq5rZmbnbF9fCQ7RS4JJ5wlkv9WTl4ROrbt00Y41C32DANvAC
xCB/XrCzqq7BZ5kH3n612EXkSeL2cRO1hZDx7W6DCxsLGup/yE5yhcx2PHve15eylem9eI8lO9zh
MQdNbI0Zg3H6f7I9ShkawpIOooqcD3/OHM2+J5KWP+GNWdCa/uy0iuSTCE+F/uGR2I7iAllPqMQk
z+MhB997XUHNugEsxDhKyHDDkAY46RGuxjBIXYJtsJA6vqi2XUcdqzYZl9XWqzie1CfkpAN3Rasm
nyM9WHJkwCszGlkpKoj83CPZs0g8Mqj6ksHhMpq+oqgrg7uFAuth/IBpaB18k/l+qgjWanz25xuJ
JGfprWuv0duMKXyhAP9LMiqc8ycs73xnnybIwmvLH0gZUED3SeKPfGn6tciIgHckgwOVQXnxaxkR
lmi7I+Y2UxaBLrHZRgMjNg55pK6TB6aJFu7sykYBcquJqSZxcrG3l1KAQbEsRk7FRW4CzoSZ2/+o
Mxz0JNt1n7mge4mPLPAzhAxxZrFeA8Yv8g6X2bGSvgxfvnfu3/9CadonATH8s6G+rztm4zsLRtMd
xWFZyogIWY2t9Iw3OP4l9oOlz1LIiTZhhUUXFUtMwgQgXQOXR5xR63Qwx5oxXGRFHMsY2BbnwpVT
/caWS/pQL6DDtyBLyRw1HF9CcIwKAmbQIOBEaWrjWLSMPSfS3Umt1IbgIemypXDLKH3HIRVLKQ+T
60zgXzcO6hVzb50MtqQL93suAFE4vQCDGmWob5JPSPZ7L3m7km4YuwcMJDFth7avF0vl5pgocCba
8qFuDriTY1QMMrmYeU0CstLlrtuRR5WCqwVoYrBj+d+5lgN5XjzsVlfNAR1uXWT2IEHUpKzpkgjs
I/XoIr55DptainDXNPX7AL28ySQ4+HKNMmy5F3aJxTqhEVxaz1ODVMz9hOcg8rXc8NxnAqefaOF/
BL2p7mFW/zkXA+ygjqYl+Ivb8UmqSQI39jLbMoq+mSxIf4D4iZZAG0aHudKqHGFyAlNeHepklgY+
hM44nMCemMrJzrS1XW81oApEKd/rTBau99Hq4F/JeEIXG9yJw0OQJqPQc7fj2Chj9kDuCXtRnOvE
ajDGzHUJUuYSiQOHT9mkv7PIZ6ViQYDJ+sLiFeXOQa8P8BowxbNcQLaLHRnBC+lhtsX8nhpfX5lp
MpYBFjww/funzGQRe2Y/oWMSsFcvnKZweKKHx0eV1eS3BKkS0IQP6NH0G2w+xocqdHOHgSQezDL3
bPtmq+rhwrJq/HGeZrwMljoNhrvE/n199awGLduEVM0bpEUZXUkdx22mlmm+xj2dm6IJZeQVLNcF
bP4YN5MdrXeBJ1RTbT+KY9auAXOy6HsKhSnsO7YM0WROxrm/FlsqzHGL/WwIq5eAKiHuX6HP7STg
fvxjgO6beX2nGGIJ2cILqqIp94MvtDFDD39QaCKj+dfz2M65PMqfsZPx7aNNAfU9iR39VJuubtUp
Nf+JTx6lfNoMEHRNdojnH2hAdyKt4iAGYHozG3tTeYIHn3J4oEiev0R2mw7pczJk8rFUNJzWSQjg
kf/8+U9onZw0HLejGC/wgxqub3Kx2wf+ivDZbIVjLt0xWk7XBNu3BAbB2I92QLoN9ciCTk9+l7Qo
5jfYTfobvQZMVSjIr8EKN+aJ9SCgoQG54nVUZn7lmCHu2PSUuNZ+4TU7jJ3F+ZIoo3p5RlvMq2LG
/qU09ipPbGnMHceTBuouMtt2NsSOlADA/C4r679EB7coRfQk3+ahw+a+b18JQC+2qeNV/nZo8R4x
9RGcKNN6Ph1Jk1M1mcTXy1j4YGbGqkAGTxl08RppyNQOu4Ls9boKYuJmO2Ninf4qU9bIacjHb4BM
5ZMSLMiwR10AEdQIXsOktI0G2k+RTHK3CfubM7Ie59C95yngxYv9yYi2E3DMyDnmIzCcwv9LFB1Q
vahY1G7iIjt1KQeYPS7g+GweIwpC906DNKSa5WtDavTI1JQR7w7e53hWgvg4WaMIMCqmlNiS5bfb
oZ0leTu6Zac/GTBVHn4OhEVc7SjSQ14IVscT9sMDSNg5sesNs4b/t89sB6t8Eykjx9jlMeqL06/z
FJaKoaX0Zcpr0gu6Xb13W+SUUiJFNl3alYaB0NsvpvX8aICsmI+YmiRCbTV/s7f3ohVv5qwWoZ5f
E5YAXP6rer+XBilzlkAGtDyVmyi7mJ5hnkqV7TzQZZq08svw2W4p//LwXttcU2S3Ekbxsl4Ul6TF
hMYmvSttWJ6Ou2fGTOdwz3ip3eABZlrHQ35DBxsyIxzx+DtHH9LAuodx+zZFfCs+iRQOuPOqoELG
qNbCo8R19l5nidUL3LtNR+ihNGqP03OEjNTrG7JOBc0Gn+efIUQGJnC1GR3m8hdwg8/+jg8HwJHW
7zt0WoItwKD2kgunwVmgYBIMJiTdjIXg0oi7zUe7ixBsZc9fjNV8wzJG8LSoV2PGtzrLwErOh2hd
mElO6qSXiLibuRZIujMwq9mJMXXrWELcnCN5MmlxFGwGXMZ3Duqo/rIc3eos7U95AydDNvQ9R500
8HSJelOGmR3NagbK7tTAzAy0xK3pjbQMj85Q+foqtZ8pGtq/N8RHzvh+Rciomc1iZF6lmhAXfJvC
zoKVxoWfzk9978sE7ivYQPR3vDPIbIPmUQkLPGSF5veK+Nsn+fk9NxW/7YKhtgMcodZX01rKjA1l
1UEOlpWBxxTPKiWe19JnZNtzm7khyvxs5x7fGyJxss1wMowFwgChsLVFcQb8yodRGD9GNoz2bfyj
InkuFJUYmOvZ+v/Fgl5R9DooGa7TWYarF9m3xgNTHZ2VFDJZNVCIi10G4NvN8QfFOYqkU1PgSXLe
BIAkuaosLdssL42+eG4Sn3YP+rKA5chrc6E7YGL9sDckVJd5ykeXEoRVztSmG34mJpxG7viZgQr8
VSV9sGbpEZ1w63yG+ZgisqxZVaYPxSS9lP62344/BQOU2QZbKuuSzumu5/rR5laciZ1pmXlOK3vJ
0IJyCYgkvrphAV6HjO9cgGsuYoXTDn0sO1ALEz5+Xv2MSH2KMdN7NqlbL3MJ+WSqiVH100HnXmiG
UCDGSxzPRKjZPkOYIa8WBqWWls9GKL8McWjdhzeq0QTyK5Ym7YPtjWbVsB9z0dokqqyn1dNXM0TJ
2QCvQ+U53ow3mIqWUwlAgz1Ow3Ejcrel6MqTX/OLDnivBfRNM7n//BOkNgj9FaEJIJD+rY6ioVqk
8H54Yf0AgxoXdWdeKgsvMDfakPm9oaVFPY+5pE0ZbISTus9FOpgnh+nu3/iTcWQauQAsLsH8p0qs
ySg9yb4fgbvtRGhWanvp5Q0udZ+lGMAcdSNCro/egpB6gKhW6igEIki6dA7UhC1obKDf0JzQn0Yk
cRy0sPtXzdST9RjUMbZpb02KViHCLl+02///vPWQj6ntSZntoOFMuz3b24cOMiLkgdBZibMBxGRK
4tJ9vAbcx2lmV52LSyC18gOtw6s2FlpCu8ceV0xY1eDHDIPHrwrDMNUvuDahgRRkvkpp3WWEWm4Q
9pTs+NzWX0GSnrnpNeKJalqCwcFkATWvdwYRpD/Mq3N3ZkEBlj6jkiysSvRK7ec5R6nG8Ayhw6Ry
skxKHMZdizFIQc5HZr7e6kO9LcnEObWFLGT/VL6GTEXKQg+zvMnonUt13qzbSrAZja4DH8k4PJw/
jRJ+lDjU0rFD+WrZKFzq5EpLzxMlMwHfHB7RG/pI8vEMaIqz5MmarSgHG9kopQNcNOFcVJDvrBJP
Djy/jAivyXMB/oatHe9aCgHlpJ2hMbj2Ayt8whyKKnJVJtb7SWJy5fs/5i6HHIHzELM7gA6zXRxM
vOM3iiNHgDlggc9zkWO987YTzyrzeSgi2iGHs4WJpyOWDB5G6GWHAwh3lqSsOgdiN6F46gNdqh9h
dge8L6K1/yEUr6/diSrdbE4jr95UddJ17rhEnaNnoOFSB70uCaObJpko0aBUFYoQrjDeGETE//Jh
daSGLXPsNF3tM5QfXioo2GzLzohOjK60xTaSfFuinEQ3sSqieJCpgzoVMoJMiMN+Lyotm3ohsjyE
inIEUIo8OccaGHU5KgUR6mNZmdmsjuUwkOJOf4RJ8JKSxY/W2Ngt6qgpHkVjeKXZN3C+3Fzcaszx
Ml+GyNCyAXqoLHTVN3VT4LAzMyqFRL8u0uhvNCCca0ZJk7krVKD3lqUnUDVDmNfXn+gYLNe9lXCr
ITuAcvhjBBLmjC5jgaZyHyHKPtC2Lpju2ACqCvmmLaWA8ixIzY4T6H+Oqy6sNiO5FyEZGhsXXeMa
FwaMBZBDwpalO39PspE+dFtc25YwX6l37hHC7FxTJQHYa1qRDTaMo4t1XQX43yNMD4ZYly7um3q0
iBQ6yhJEpZ8ZYs9i+ojzIdyMePbYmXUtvBe0XtiB2+tmBfNOXV/u4g2sYb1gqRK9Btb2FeW7YmQ/
/eikg7eshy/XkCSd28GGQ5KEcwXrAVjAbW5n1Qiy3eniK0c5CbOqxwroUEIi/8KCspKvvoRWTSqO
heyP1O7rYHbe0mPw+tjIKWDUICLq/ciHeSLzvSXl5Ak19Wdbj+DRlAgSrs11NdjjWYKJ385mhhcq
yvz/h8qP8SU/OWg5RgmSYA9gMKMEaODauSACb5lBdaK2XnkVfkVTnhpcYYyRarkjEhL86SQT8UO2
l0RRDBcm5yPsnX433je1pyescpGqi2EzAgXkTFjWQf1EjESxjpaUu2rCJt0PnpWYT1srvdTp4I3y
Oyfo5bVbWAZsKjmUD56gVPaetKgARZQKAHczvPgzj9vGjcshJlSeb+eKUJjzwDizEdqjv6ajLC35
Z3LkmEiZKCmmcfqRB7WMnE0iKjglPxx64fzm5Nu0Of90qCGwAJwl57DCe5Mca7y9qCR5XTCaETs+
0XPzyBbJj5/GyLdkwL899lAOEWahDhBhSdWwtssMFUkujfY70VuLR2dWUp1xRhmsGAxYnEpB8Rrg
yRiWsNqT8PPggL3kPi1dNwUYssQxsq5HS7psXWio8ZLQ4urr+hcZRh2oU1DVJ2RVBMM22Ub/Dy0r
V+lyfKS1eYydxaVLkNX+VzDJQpvh4iIsIz3/BT+gVEObe8M28urZJPdYS+Z6K6x9MGAsSjkvNJEh
kzKHy7mlXhv4MCQKNYSfwUWc5iHfIJJtzJHqVRH/KTwsjHzDz9OuX5cGbUpCl9nuXynWZsMSlzGl
Mv7jirUC07Lwa7GROa5aUeQnI3sul9Nen0698Xpg5n/qyokWHOOOE3vxx6lRYCJu7BG76zHH3+/6
G08rI7HU1BKUUH5DvG4wVc3X0xk+CH1c+rQQuJ4QyIHnjwPU3Nl9LBsNCS0FJ/yjU0oUm5DIhjzn
gaSV+TCggw6ky4eNa0SeuVOVpOFHZgmaDvMQbblzL0iW+IkUKkj0gfkbT3quGw+37L8bxC57SYzu
j5WQGET4QMK1zFgVR8cn/5IQZAlL8Hj2aQuj6jtR3NmJqucXWsE5ATdulsM8h4/MWXQFCXhtKNVO
+GO/j/xbw6MZSKy3Sk4KcJkGetXaqQ3z3BmgV8ryjeB41QgUMHyrm+L4Us4E5H83Bo2ZxrC2FNDb
+bLtiLAXs1giK7eY1rkCkoReNNmzK+Fy29S4Jo4KjwoMS37zmgNf8XuWk/0hO8I+5lHIum4+5V3V
gVox+Ozl7l8Uvdk5cy3CaMfkI+p+RWubNmXF81z4IjqG0o4blI0i/I4VnWDxZ1LRPP7cvqQFtBDX
7ZQ3cxzkjazjiGkxCHCpA6Ed5zzx3FMxz93qq7be8Ml2YGV2jRLvRpHIIPyTQX++xSFAqCsJ9VUa
EjsPK5x9ixBWqQEdcwzvuIA7bdrgJ+SYRkUrB2pAI068EifkbiljVf4aNe75dm+em1mX2AQwg7OW
FZXuzNegww0ffuRu/8KMaC409lKLU9xsrLElieoARhpQvAemDzpohfqr5I+AwLwDF2Btij9hQdk7
hiHLjLUOfVQx9lNkpZEeHOER8Kigepe1v8Uo0BY1oP12F3W66O8hDT8UNjfCdrMc6a81x08k/Kc1
GzQNKEzG9dvvp17BrDx2kwBnI5F15V7PwWLb1s1UP/CCU0nTEwOH1a0GYqMndOmUj7tPH2E7Scnv
oCia26HLEw/pv5qp3UrvBLcOko5x5YCJ89uIh5E6wb2MDNWjr69kDzdyt8kk2xvYOJTi7kmEUjFx
/Le4RIaDLLv0Sprhxf7RG02VgI/kt8uGaC43TMjvV8N+qaxvZK07nl4tXN4qMd+vThfP1ips5ovi
dRZ4jF1aW18xusZXJwd7vjxIqz9RFuPyDflAFDu8wn0BiHri9RuJdoGEbM6bd4/SBt6gnDOpL2Dr
RKQ8EW/SnIFqhXKOyJPZQAnmRARrBmJn9J+p7mdnK3WeD7Mm6H7pwWnlY8bahI2kMriw+qoMzgWl
/BhcWzDEPXUWeOCgtREOXyRZxObihNjQpnyYEzculrAV4H1Vm5ff9VvCrV4lq1BX6BtIw96hRjN0
nBmEqbW1GYOWFBKBUg0d/Z34/iUEl4wIYKDDOpwmSpyuQgQiPkpKyTXKT8+2SPuvVRbjrj6mZHbY
Bt3WhYICEAvq/fPrqZtzUPAJwBdgMboqzQFIAlkkZQEOmRbv0cTC4rIYpsB0S74ZJTgDd0WBy+hX
1Wq5iStdvexn6vUofanc+/QioMYTk1Bcn2BWOfLNy8Bh1qXfjYiXeDOZJUpLcrj9BPFWC754os9H
tMxXweTW8fPv1binr8MLYJ61QO77OjxuPblEu/wo2+66dSiRk97wZ2EYxZIqxwFoWH0w5qwsi7Jh
bvWKBXC7RJtEKqnQeH1YMme80b5aaSG7k1r+yIYKmQfff5k9K+3RvIbK89Ahw34PXvy/tRGr7H7J
a+AiiHespzqsna1daRBtyNlj7yJ0fw6Ff8x8SKvuTtdoFcT0aMg4b5zk9swdR7shbvyrWsaDmswB
qlG+KrI8USuJQGX+jWKj4g7/A2TvD7HnZhosC8w1hwntr3Hi7iMh4WUlGbE3hx3XSnpzl6kBmHgp
nWAV50lzNb6VzPTZ5rNqWcRNr6n8HCR6ciqmLbV/Job4BzI+VJvQvvKm4aMA43L9dXkK77iW1hVi
OR7UuvLdukN/RfDpFIm+LEN3HTMQsvZU8VgFNMmBqDDXlt7Hl5/jyaeUmrOlHWxcPbxmG5y8gLD0
on6dKuGt2iseJ9N3EkVrxKS7aRxf/LbFaliHvTCzlV83Ukf2UuoVp1yuj4KKUZLycvMX0XXdgtBN
0Ai54rPgMpuGS+1y1SsMqixyeVqfYkknqpa+RYsKggxpGDUw1T/LLBl2czLduny/wipyCBksV6F1
TjQDmW5X7jbWSXQR7UiZISOp9NDeFal2rCTS9B90CMdesGikahE9SP70ZA5vPBz+dZFJ3t1d/fMW
IrsaVyfUe5ZOeI9AqDNUaDReJfPIwlw1ZKLCMJBkyuoiJ/GoOk6mn0glLcvO6CmL0ovR78P4HpA6
Fz+h3tfdzXkWvyhpB4MrfDWPSHEDagFW4YPPGk/iALrPnH0R+C9GzCg1YsIz6tucMoXzcle3y2qQ
n/KAdVZs8F0RaukLuYj+5Cgkmi04fy937XlzY5tdJwJ52fe3ec123y2w8lO4AYHLcJHnFO/R8WVs
WmJuy9RC3bzblaUJ9gIoSfmXCumEi3CTd7r2ZckoNb25CEAhKzCfY3saejktliGMLMPoZMmQPDF/
WeVS3oloyLHZ+oUkdNObYHOzlSRWhIlb0LwxthFgARfDmLMnbvmHpBHlAZ8FDKaTqaJ/wQJyFPn7
mJt8OBCJ5ZRUWKEx9cOUxwAzer1JCESuhBw11duQi3aLL3gsn4DQe10ScG08rr9t3Z5akyhSVb0m
OqIPaJM6SlBYq1coYZ65Gik7zLks6R53zPE9mhY3V8+gy7a210NE/E/1i/5D3yldr424JcI4WVJP
XVGO/k6V5n8shjE0yzcvuxqYGTNKona0eoSlVaRA33UYvBlJDEjuDNm6upaeHZ5Jx4pxr4bJHbfC
hcJmVTGTssWjmWC+6PQNiFoBPi3PQQs/PtxohUquushPPFa0375ClDZNm2r+cOVHOB+po/+fIDNU
WDQTKMbPPCKCO5qGYjOoJSUW3KKQG7NMgxq6iWXn87EIsUeliRTZ09pMjWBCzZ2ODwHn3vEO/tAd
HsgjV2Ivp22ef+IHeRDvJeQjPWrKI8nhP++2412PJuyw5sV0XEcmD//T+uxZBksZkIVoQ3Ol0Uqo
8yhg0Eb9mfNMiSc116r9YJvZeS1RwMXvcqKOqKKBN5XDrAROiOiR1K19iS6veNiCHOwBPIuXrdBZ
U0nSIh8EHKLKUjaFpMvqLt2s1IRDkwVyqofpGSwLyl0fu4ozzZ1l5gMEQetnlYWTOxq1NkGqDqQm
ZiYiy6uCuS90YOYuB/uNCIVPegK6FnSDPPlzFCqqwRdFEfIJtjYdLgbBv0NhI+y5HrnbcH1M8y6W
x8kGQOxCSptuhEFgmU2CAMLJB74nRVaFmxbWGDUsoi7ibit6uFd1w212fwpdzr8tpTTJG2P89PNz
oRvNaNck83jHTLAwvMneUU2KqCjZQCRvj7aLsChx/V6/yXLqn+bGCnW+7zlgrYIXwz4/EtcsfxgQ
Nzm4veSBNa2WO098opMavYZXHB8Ud3rrHCgg+9ONP2M5Y9KwhCbFzkk/UpgWp0EwREy546AorP3c
GQEIor8aIRGZ6bxNgpJlN7/hyyxLMXQD/CSkodhSHLVIICIldQVfHlSX5tQVQ12xuqOJK1PB+6IJ
PB991A49oANER2msgr9QTNrknTrY9HIzlLAFkweKcurSp2nV2y+RMCCHrk+B1pzTf1r93ickUXY2
c48OmtnNTs2uul8OZvI9RAsibBV7GAvLtQbQeRssd7CoCFr1R1WIu4+OfJPv6zjYnlr8K9scS2TH
tZ5PuwSNWuQ9sB61GnLnMOhvLQI1OFpEY1m879+EMF6YFPv72DNWmAvM80GH6TvdmteOWTY14sg0
3wDYQpVrd17J4QjrVxVhqA55S29MvvZSbeTi7KOKYRgi1pPZfi1AF4S6UXu3163/Tza6u+UWllUX
ByCfkksNYGiALgopjU9eUGGCtS8338r0TNpcuF/BTX8r41se2PSAvJhLf2AxuR4E0Ir1wnnk6WQ9
ob6Bqb3ZiU+feRX8a/geQ6nXFtFG5q2vmSfX6JZtylyF7e66xe8SBl/8Cz4DNAPJL2+L6FJaga9Q
lC5xFKOU4XW7JX2aw/c29uIFRY7TKs3mEnZbl9LDAcr/qeT0X0ia/x4t9yJfmVr9UVIWQM8bBXD9
m8IDtCITOVrC/W+YwY5AFDf7lyF+caJrCOZKZwpMOkw7aVYVpFus9lJ1re7mSSpNmVz/kUiGKEzZ
FS1MdzpNLBn3Pp3JccRUM40YgReefz+XDi1hIAs5W4bAwdwMQzifmT3C9L7tUlxPaOIvVjMOkkDT
sTLvgu+my4Yyb/DB/4KOo0JJDNyMYu9tj7P7Duf5qvdPK1b2McYdrg6TyGBNOc6gQI2piqVkOV/o
THkjyIPGKaxXb9nKRfi2RC3tceHr8xOuKOE/Q9pEQuw6WxW9R9g0+/q7sRwg8H7y0OAiVDSXDvTz
w4WTAnZ7dCzVNJy4pWwl+p6dASHMCodMxRXX8+bQV1G/wHUaZBtfDwYVq421w2dzSMQf+2THTHLC
w7YdrNu66hlN0PDXzejjER+FRXbSMcWX4Ouwsost/F3NGZmOliHuazdzzR+Mgfc++zrL3eLUYSk3
CELfXAt+GDecOfRkAaz4pTUGvz+I3URLFYW8bwLb6erKU/1XUnTknonK0VuH/lLPCcgUL3Aa3N+s
n2DKbJy+7I1dN1M7jvqMIHUr9CG2rf9bRZOZVedZiKluuulB+xy1UmCfcb/SrIOcgNTumKKImSqE
oOeSGrMK8JyCQj58Hz/O/58MT0h3TosRnQvnmmAMVeV4GX+rQSh2VFR69nxA6VHFv/n9+prUv2fz
emlQWnhF5qVOaBrvDPaRpz7e5dEOV9bmbOyoip4Fd53+0Yn3g6CpK5ovuAP2JSxfqx7UXih6Gnq+
j5v7YoHFAco/v034GLDD3DsHuBGXyFhph86uBTB3X7jTFMTAxg9Rcz1lYrAq9EHXW/A5VLYo3vSY
gdSfrJx7+HeV3dxpsQpYsja3wKG8h8qTW6Rr/7BTD3x8/2n1RLsy6Ds7dVH8qbT0PvBAmAgU0Ofh
KVS4Q93pnU035lUIptHtqeFXMKXKNORNz14eumwTAu+efIUEIOHxLusEjicWW5qtl+fYaDgxSnPj
o/HGpUVPR3IGV5Ms08/qE1Y81PtX0tEJtq7WFhQ4+0PKE4bGwYsHsv/LX2u9PKpFfTk5NATpF4q1
F/D7vTtB9dfXZHZvf6YjcYcx71UzelsJLPMQq/3G3qzQfh8wuOObuiOuPTj6bbzDxvk9y2XdjBO2
FCTbxLqn5BxxToQ3xipQ1GnYtlq965pbCnME9nuvcc4X763WkeSEqOB70Vay65/cvAU5yv5VJKvo
VTuS1unEoJx7i/aE2qnqCRZMJYX4Uasyyvo9N2IWkb1Sys3gQOBg9i9TKn0PPWSa1PeKOsSaLeWy
goLaaewPLYSroul41mHlNiwEnsprnCxy7ACyofGoHHUDh523lXAo3q/xa1tkSqeeKPyZpG/rsdpk
RQfT6FY2yA2xeeEa4wfR8C7BajK05AvxeB4mw3t2lDLGN7xZPCOy/9GJvttGabvErD1UMjo+0fA8
spm+AymL3t9sKa/eZL6+vf1ysIdangavR8/lTzvX6ynTOrdyAD+xiAa8awO7eRX3jlxH1bQMQT9H
N13y+gHpMhY4KJSXjJ3OFIcgwbxcywh+JegpmMvXWUEzUJwiyonz5o8QCLKjTI+QR7bnu2DnTI3M
htCD/MxBtrLu5o/dbuD9/uFVh07H2VhDZxOnXOOvx40hINbX9KP0g7NgM+vlKw6FFEMj+Af7GbdP
w+YUd6n1Esv6DAY82dPUnlbUfYjgjztrU/73ZFd3UiW7b0OJjwkJZL2YyRsMFRZxeAApQNBq9pLP
ZexjN6n8YOgK7ZuPmpYXOjO9Sux7sQz14G1kQwXlO3vcchwKn8Wj9ioS+Q/oB1oY4oEudkIlV4gz
UfGoi03Ag3gdJGNw03Bn23UrLERLF58FoiCAYT6eC6+qovmm/Bd+cNZdvjGggDhnzV8xEsJhGby0
H+fqK4I3iwcOvN3RpqZZaspekA3Jh8BpgheS/wIIkRAoOKLWq26FBfcHhAlMy5FxDO/CYQfdXMJx
jb5RyNyPW+pcGeb1WXbesC7G/czbqiGkvl62YzwVdG0z1tZwfzv0qQ0NLxY6PMx7Pp9HFvp0l3HN
yKNsxvzDbWd5jBBlZwh4btZSirFzf6TCeRehufzmRZsFJqDBIJD1NPEskwN2OE9gV1owbHqHM1x0
0loK8Fna4zaqWhJgTmlVODQi3JYrmNIc5+IW4KzWNpzIKezQ4EsZEfmi55klRUmhHqqP0GX1dBII
Aaj7rv1jQ5NEjSHAgY2i6trMs9xHwXULp7HUBJx6BlndRaTr6QgOWiiD5lqMJM/gB0ZohDoHrmHu
syuIeyP3GpyNGAmJAAmE3gAd9YHCPH3WEPrgwEcKJiHeCB8QMqPtrpMUDhbzIHzJpDMTZVp/1llE
THTZ5SyqvYc6A6UkTxCLQ4qd9EWJ0tlVOpQYEjQAJG6kQgvRUU1vFdbyVIpWtbOYOGJai751nAlV
R50IULcu+3hFJDKMPGsYiQMrEI9fN0pUQUaNGxSCubYubmpif8vUA+nnBnatlOROFGnYgZLX2htc
8LhiMo7icsQoXJmmU8WqOSKZoU6DMPTfDBTI5uLZZGuYj7vNXLwkxubRH8vpT+c5urCqjvZosz1/
5GldWRaXpanJ7jfooqb9LQLluRHMA+gkqR9nLm3teCX4ts4LIlh9YPxReNpU4qRrXjxI48RbrOZ3
qenFL7tlSqQXEVVb4KxkcK8zDWSIdLYxX9KOwsd4zK0IUFvUZoaixMJQOhQ37cgfcWmby5ggezGG
fGuTYZ0ZPjQYBed+pB7RLusU2MzhMzFKuRMb1JXKiEi9tXHYx1KimSZCSLOXDOjyBh20VvyJ+R9Z
pWHJFt3y/ya5g3iE0SRzRl0HohX1ZikBkVh10IBoYH564Or9yycxcslW8xx13A6o02fF2QOjaCMQ
zC4fWlterOrL0oB7Io9s75Twt3SurWZxwSYBQsnYqE68RDVNz/x9QKcj9Q0s65txXeLVl4grIBfZ
zCp/aPz7psnP0rV0ADmVpJgk8TYY/VnAOuOa7xvdCsLBFCJOcPcKpUxvycbYMn9kRDYIA/ms4exM
MoPsHgZ/FltAkgCmbJiW2viW/nYnLwrkBpB4w9YtEuIi9nH0bn/k+nLfbdbfQ373shQ96a+eCPls
dc8KK7BJNaB2VTdJ3sglHfW4KZbJo4LarrpDAN6/zlcatWJKdTpvV/YrtQlwJnBz47p6cAg0pWeV
WFA0Tz/Y/TpnRRmJhBJz0jpF5w5UAcFVX7gT+0vm2d1krxPL5rCYGMqzkFPoZXwtQUyfPVSSh7RA
2Pe3Yd4ZkG0ASc/5EbHCm8lkW//3gBSYarTtviQEPd9JdhLfLof2yFi6Egmis3jhUGPtJkggB0kM
n8kTiRe5ZKrQ1X4X5XTLMr3RUm24kcXkTbQYVDeaq7f5CKgisDOuBrTmGoNtADxQmHt8ctkZv/e5
YX8zEJ3tGlu0oTwdp9TKmj4fu3IBVml5aBv6J8CXw+lvYny0RFUc8IxQfs9myBZOZmW8R7zDzk94
rugs+s6CONlw74BsgCgEd1YWLPHXMgSYB6gdVZ781PPc/D7jKdwjVAKb1i8prr7DUaQ6K3md2SXG
kY8Tyw47BW/zeAOZzJyEHlzkMliUvvoy+iumXqglD1I9RMj3hSK62+2XTpNaGK22Q5uiuD58A/v4
WehVJK6sM7tki+N0HAZ10/nlpvcrWWXrAWOAt3kCOQZJKCqCv8jB9gaVGWMbyh+D0N1IPZJxqdDq
u8n7VzaZe5hsNNczHk6LmVNjs8GCH/cYvWZX8y0ZF18TcxrLqqfeoLVQjK7OjLoZfQi3Ih4PgfBF
YYHIkogfRBpH+6H+tzEPxySL/jXSaRv71LS6PXXgGhAFyR+zXQ3NmQ1xG6CM0MMQgF4cUqKEuzNB
8RuqsQkSJbOsX4JHUx0mw8ZrCjnJUtCvfQbVC7RiE7S5C3ykM8uRU9hBBlphWAOj7yd6G9OKP7oQ
hO3gTNRnlKSLh5+xyrOTLhedYecpbROjucfuewlSfsCQz72+JXiITGwdAYaBg6BEVuwDd/alyX7I
ZT2rxga3BsFcalqYkVPmkeKJqPlonFmtIyRYPWRJCuUKGDww4jcCZVr3a+ad8YG/P7BeDdMWkBk0
EcHJ2cSPqo1e+W4cgTD7s7QXoAULrBGonghAxXlqevkJnnxZyLCsaaOKQ8ru+lm52NxQVYrd5j66
ndiO5DDfesp1S7Mgl8rXp6GvzPCTIRPDcIxQMVB2IyurZG5wLxCKLppkEoOYA7bJ1DzmSBu8KcyW
QiZplMYi9K0U1J1wZ0T0r6xV5qHn0aSmzhjd2KfWE0L/m5SaReeHHIsGmDnR//rBWOdL8TqZHiCQ
jZ8kehYPxS7iHl7P6gbLsPpdFzXgK5oeGue85Qx1PfXVckCFmlPkf775mij69aNPbo1eEgcRE93x
a6XZZo7px32WOdahs29FlLx7hpZ8MYX1wVjUPErNqWFV0wBZ8QTqrer0XdVgPIK9WyKN7wjlcFTZ
RL44vygXIina/Hvbtum9M16wbjdcobeLQAc9mwQ2ZtzbEG/BbhPPh6F+UxZB2WLg7pl1Sxx8rYhL
3lEztTfR3809CdthYCNZi89guFFSAwNjLaNxaDmJQHrbLoSAOGv9oUEs9Y/aNg0Cm4ANGCUvqt7l
u2yqeeEUpTh37mB7YIDgzSpSlRKz9QC2xnUpCO+vPHF3zefLh8TXFpFpZtsYjb453NivtYgDBnuF
g/x5S783bNS+1nA7r+ArePb0LvBXIJfD4w0xu3NCQsTLs1aUb8KA9j7NgXUElhhjnHUdcUm3EmxU
s9sn9gK3Nt/UEW/Y4rka+MQaZhh6pvXNRXpV4tgZDwwNxMjt/3tIdvQcgTij74rhzOqUM3Jz3Z5c
kUFpIUpef35W5f+mmAJHzA8xFIoQTasV2lShFm59fisWIwLPKffauUqDI1FKgzhCASTc3rszza6y
J/Kxx5Nmbj3Y4UnLzz08u5VMlMpfs9xfQsFXGmIHRYOQIjsn8xpypBvO/LAzHeXtoXbPS34zNY0Y
TUjDrls7as6nuSROIVeqY9S86GAI7s2mWbzL1xomv7yQB4hZbPHunivA4LvxatbALmfm6cP2hGPa
MMW5KkR1R42S3gDRBjpVyGa6NV7pGDkJUpIhCyGxP4P2zlgVMzaP7tJwZ8U7DO1c3b+9dg30KTkK
tKeQPdtUerdierCifd+Z3yt3hBiGRPeWPtncaU7FadIIUgCm6fcDOM3zZ6FPb1x1V+dnZDXtZvfI
ea5Dq0bzTmbg126p1jP4ZP56Ldg3gEtEg0ueAIo1V5qhmQo+yzv9AoARQLisrbpjZ61Yn1LXoAhO
E4AqSVs3x++UK+ucvEU5nRQ3e+Z+wfmxvLcze/uE0EbmC/mvLzNpk7ZVtibNfGspMt8DmYrIaep/
mzXkeknDrbbK8nkvSi96ht3WX8D3kHriwwz12sJYjmy4jPqtMHr9dK4UeCi0pTY9Za22r22qKh6M
WhFF8D2kstrKqr9zdkvAT7M0Swpoz2gjZ0C06KLlKihi64WGhYj8k/zwNxEJKapOUYWDVBwGIpha
VtJDfac9dMawVlM5kUN110k2ZBAHc6E1MkiGc7D0jDGhx6HacwSnarGq5KLrMTVgd1xZAH+RgUjl
uuQKjGmkliMuIJNL/VsmrLV13QDnUQ2EIQWxYIcSSAaTrqsikgJGy0DmmMWE0ycLQY/s7CtuGbvZ
d4q8DEudbOj/4n6IaSOY/ZI8CCo29WN+Rsdsjg+zo+Sl3sQII6D3CmFtNUryxYOWS3BRBpEvPYTf
URKsXw8MlLRqtLE0xjuZcMzxYYp1p28LZtZGOZ6DmpKD7icXIOr4wNPrWYoLRYIsQIqBCQC3wRjl
ApvbSwe4EQ+8YBtoa9/SDtZ+J0UevVf8sQuywwxXvptcjBmKVYZqmSj4fwr0hOWYfdl++9T/nsE3
h2gOvDPFal0w2Kt3BL5d82Svg2FtHe0fR/7o2SHoqMDhoVHNT8g6Lx96EAXsj+i0ighFpF9jjwLC
Re9/0uHXwSnn2RFsJ/5Kp5nT//Ml3kjnwGrpmDkZE5a9A42RXEp6uW8UERjq6KrgClx38DXs1XkV
WkoXrdF3YDIe4glPI1Ca9pPz03Ym8HFbLjwsH8dX3848nMcgLUEtMVRm5KNUBkGZSUVGRHGPuTLI
1io6ip6eg/v2Bl7fSV7j+1nc32dnioJeNgGMLLDj2iNrUpz1SwzVBoVMrynfMqjo0tLN6b+N4v3W
xiMBf8+qh+zYvhgBn40RtO9TVpqKndZI4JaUMXod3nH0048lG9sM0E44pEVxbX5MEB5/+jBY2vXs
hnICHn0bdxRfg6smVUll7Y4WXruX68rU9Yk0AnQpyjm1lWKO/u+g0CyqCgbqka8qMoiDQV+WQHQV
dNVeMZeHJiMHfiRX+tgE2ADVUDaWvw0ucVpHLVi/LpX1qAEbhcKRrmMWo9sjfVhtxqCrAnyVe6YT
2ig/Nxa1EYuQTvfxa1c5gHJyOIN2E0iu4FvwrM/vttSdItWXznS78lZAccgbLqeBFczt7GesGVbH
6i82DxCugMqJd8fCNCnIUera5SK/r370ZnUf9Kb0sko/55/bpy1m321rUoreY2J7ZeiMleSqRCRy
ypXDLU0SDLqwBBe+bmHgTutDlOP/Zfa3zVuO4pooz4G60/hQlULtBjoNg8zEtter4hLYCJT0jJ2t
Jdgkrv5u866XCGaC7DPWiAwAu9DRzsp8thdFZnE5T99GXaonuT46vF8x1LJ/5CbdnBbJWyIExhJE
qS+Sjv1FfEisEFhwAPHbPOn5eMb+PiUP835lheBsRSGOiFgDSO7W31f5yJdpFNB8DWQ9xOJJ4S6p
P9s8DDkO1mD8JrxfRsdkss41rcHwrElkYIKi6eEQ0bMTmFJCc/IQrRNHSUzQj6Bkwq+7SiB0pxlE
HqmzTo2I5a+1heJjQZ5GK+OwjFsLh3tCI895dZPBSnlTMqf3k33na+EUXjHXcrkzGH9hd4vjGeez
ORfppprCG466SyBJcHIvpfgaVtTxKSd8WE94x/cUWRjan/YuOOrmgX6aUk6Y9Qvg2n10PtiBqBZ8
YcVUf5GJLpdK3mtXgwXzCzSjqdaPqvZjqm3zQ5aoct5bPGRYXJvSQPJwhW6qACwj6UZn1Caa44kl
iw2edbbwnntpjXToK1u2jNCbGjQaUr3aUtI8i9+Vtha19aEkdF0wBm/UMWG0DekMgdbG02ngvMVj
MkwHiICvM8opQcF4wXBoANQpPOpthGvdDKemCiRRlkvygLcfDc/HNglinhGKysyoGpsk1OARBp8Q
zpzh1n2wsxlKxGDcdIQmHaz0tHVetyH/bFGk0DcadTG6lehdolIutZFSw8h5kdfwgNOYk5yqH3pG
/HIIh/N9RHEljyhxHfb75KNP90VumDXk0tH5RuXTEazwvuECIS6XvLmf2QNom2fwopN6VoccojZZ
JRtiYU2dR78rDU5koCSzzJSzUqgiCGEsoJp8wGSPobc3XO2EiNFsUDuYCk3rScq4mWXxsOCqGvOG
1LrMzfmLMiTPcmbcnLyNATkadb56/ZMnC+RzqQipRPzxVbHbdiaw9uQSTer6X2vZn9C/JmWKSV+R
T9bIGj8EVxnd74lcgEpIQsO4MNjkSdRD+ckAlc9mmXW80XSynB/bjKBv0Uhv62LzYUDMQ0G+ykZy
QINqumcCkwZEKp4M5hNUS33Q6RoVEibSH2d2o93HfPLxyJIzZxJd2ku4VU0zPv/BuJqBVz7ZjD08
HAxMZKPQbAM/jd3K3G04b3JMfVP0Qj9BazJQbkYY5SKlVRsD9v8wMRaj8EZVRMP/B0UnYQQkdBj7
HSKUZGrw+R+4gaB/Umv7SepRSzDSR3NyBqN0dmOlOhVk2k5TnBbqdfK3DuO3pVJfgYy4SuCmCI9S
eMvpm9xF6H56DuathhJKeut6GcdSgfI6WMCM9/ni5GYXWDU/vq8zuyMTcDx23WoV81WziLT/4kpp
uT19IO/Jl5vaMUt8npk74gSFO6sSZ5RZQ17YUo7lm8rgqN0My6hqLfFDHVWSZOIM2rKS9nBg+2xO
bl70moC2DE2x4Y44IbyQLBosyPod1UDj1+hy0ilTHaT55Q9FJIviuYCTrUwwqPbYFn/8/P9nF6L9
CX7DimWlNbraJhhXvD8mcHSCPVe8BT8SsMm/Y7sXJs2qlLjeaUesiqLFvsIL3GUi2CA87SG8Af0V
gTjA+G7FClfjC61IuCr6FiKAXTQEdpi0jN2mHjRxTwXjpiuRxqI452KBeGFXmyxSoAJEVIJjplJ2
BNR15hp217Qo2eD8KFfc04bQrhm8S1QCvph/cjGYJXvtN6CD5aIhKiEiJF8+hqDvsMpJ9J7wqF0K
uAxQAw+Bf7AfaeXPHbSLjqvaNcY629/7Q7PFVW2Qi768IvyCvK7BVHKHc6RH59CKM4XaroyAkGKu
LBGGk1UYeqRx0YlLuFM4w/LvSZoTvQS+qOWJSKyS0I1UOgRyC4Pl33oynbGbC/1s7vdAtPZ8xTUI
OTOmg9dmnn1k0NkrdCOl2SXju1NHJBMlfDpmT2lEqEac5u5r/Ql8tRzE4wbYnsscVCovRWZRTTve
dFOgSkT00NCmMhwm31rXl2Ok0g+OV7fgmbOQgrDmr9nCREtNZYDUDjPxUA+kGzf3P349mnnZ/9N+
irviV0y0gTJnWSj9LhPYNn0vmAClxAI3sqaEUC9G4py3oP3FL46RfGq3DduKXkhOu2U8hDw4v1HU
GY/eQ93Z0ZuGz5rcLEmUZ+8KX59mq1cvi5hcCnZNlOtMM0HH3krogZdasgKk/nIXPpCUYETQSYhX
YkFCX+WIyjaoOXEgdYHqzevBQQOyzUUpjX+8GE4XKWOeqaplq3hxfwmRt8wmGuGMH4U+fPRqIr7K
vFWPyvVTekTLjH/TxO8IfknRAtY/qMjDnWT448Jf0JQMwH3x7TctBjuZUJXZ6+oFyTunxMMB5+3u
eq7fetMWXbYUfa4XuXqI+3kJbhQKTqIs1bNEwIp3HE2u/7mvbnrF46RqTUqQygBrBDhKlRCYA0qV
4ypkClNQOoBaxuGxfkBvsX/St0S+UtkXCFjwsXnFx1R3LX66vkNszBqkL/+ekI8PE2sxkOvzvePp
8IMEoCtHna5baXwsKUnJ1hokDrwa4DdZbXVv62xkWpbszCQsCwugDqm/YXN3MRGF20sjw5CJ3Iso
rsVxvuwXGevxkN3cQOz4cv83R0d+RLaEcg/vyRobmgvhFFe8YufGRbN5Zi6nqOSvSXaV9vJm9zxZ
hfNkaIvDIdDUbuwOh2Kh/lVDy6PK5CbOlDXg+JLO+Z5gNAUtjk/B4bNJJQAC/ZjMMBk72mX6EowL
qGcGA6W7vRymAUyYQmWVMojMMmcMeTMd+I+teXVor5Q33lbcTChsniHupqu8tRXtmUaD3o0LJDjO
kjFd3QvShx50kg2wIB0kSbj9XBHsg49iHuFgZJv4+9B63q2QvvOaqPqQ8ochKOGn4CabV6FfPNB4
JdSoaU505j2Q2G2Hx1GIEFElk1bQRpk2TOUKQswUwCHMBRQ1d5JarwKV1ccqogzIfMuiH8xJdM46
xVywzG99P47BEI1+Kgi/uLMd0TWb34eIQ7pSrOBj4gaxZ2wYgghma8y8I3NDCJ77UK2xU3RZcFs3
ASJ1eH4xUBnXgYQQc9CoH4BPgMHJyqfAvgT4umddTqRbCll+t7VFsD60r1fFO981k8OmBAXHzFo6
AuCxe3sIMRG/Syh7iYcLuTDtHARo43nRCkXLCXv+mjwCbHBtKPdg4RBzz27fp2REeUPMcwvtOFVg
a9swKB0XLsdil238s69MlWtb/nN4K3/NrwoIdCqWj34qO+LExi18Lo2usQjdQBELC/eFPEnRciM+
yOI84DhfSFf9nRBTdrLPqN3A2YO7PLt1srfTPB13DSJYa9LpgKpfUDaoic+o2tBk09K4NFGqxVtx
zlcQTytALogr9R5U3rwT8wynIrvjNbtxOFlmdBTFLcJXIl10ouqfaBeLawhtTXhU/4flXM433roj
7zpwu1a/YeqPeCRkOl3zKA+e3y99u5Dzb85OETaWlmQu6qmXRRFHk2jlopgFvxgfqzvWLi0mmTmy
Ws4iFNjdJ/J9zuDctf4n7jR0cbbXyEe0smE/hf8QB7epo4pEpXM+FZ6Hfp9KjBQ/GFYPc1TA+DoO
AcXxBNazdzSL+9DEdTzOA7ojDC6AWpBFsmzxVby1zHjyME4AI/LoDsxG35pI9Zt7NX6/ZS7KgZoa
2lnohSAHGRIFn7NYnxl+CDf0UlmgYAocZPe/NTnhSVXgO3AqVVmdp2qwVrnNNzo/pY6vizN9Diin
BcdZ+mjhtw3Ms+l0tFUAGYXmoLmUPGP5uVFimWL/Yerp0iumP5R3fQXHfSN8JKB2tMpJgy/R58Su
bEHrEMrxxSf8Cddk4rmQ2qA8dqUxVyE280EzcleiAoqDY9LjxvSnWHN3aPblJ9fNJ473h0wH4MRB
Xth5BC6JFKlqF8dm7WwRuQTRYowfqolnoBVZKjAr06Xed2s20wN3GhKVASP1ANMoWTbiIqae4ReW
N+uV9dFzl0KA5EauucdHl04NWZ0Pn1qsFEvet83aOMJokNDeD4Ktsl/T5SWCJIre0htxFzjxmKwG
8iGUdAGsn9G3OszAcGR7e08Ai0UXL8LXGf0pq5J8g8dNEfs/YXxcQbCEVkALBpowiUiVGUnoHCRB
o8ncrLomvDPeBq1vy/qPFsDAmWE5ex6eYfKW7+X8lJPHS/2u7ukPmAOaezTa6lbPy5PjNkbTJPlN
76ywNPbXw0SWzyhqbi2fDzsjMo2n/OtYgHcjbEZUm81i4SVuDi5puB5EtpTveLF8ko2UoSSTb5MR
dxtPTXSNV36X6uFeHAhdUXaK91RMX2pqF8ojgq6tmJpzpcAYJuT6M6CaKUYKxnale/iDRR5cicPP
CDlEzMj0BJcUdKr8eTa84SHYsJApS1Uurbh62Nf1+gdtptvjcv57uo9WiydNkTHDKcezw1zZWEiE
gYw9LRxs9gQS9giCZi7Cd+AM6nF0LF3hebdszUJRMPymBnnNglekkMntV/TwypMHcfuqytldsmP3
8nF7/iAaFMxvk5OTzicARLWznXmiIid634WoFJ0ZhoRARc2IUgNmIBmTbvY2asrsPvVeaaprYyRF
70DiMhQ5qoAEeHwmUUygZRHlEGNUkizyUSBk6mKbcQlBgqevxT9cuNA+61e7bHENNawsgUjtshDt
0yU5srEYL2Qul3g71fk1rJfjvBvrVpwdR1sbhPy1WMqHMwIu0SlrcPlYLp3sp4XiTRzS9F7lc3I1
9Eg6cM51rP+97mftl2WyuMAg7/VFSfx7b4KWwvWzQ0T1Cd9kwskLDDxWB2IhnfwLobqqPt8WdGhl
VLg36hX1roN8iLytWJVVwB7MSt7fY4HSfPJGa21NRgpAhNIFRWIDJqed1Vb9TXTknDw+Q/vSmCSH
NhGZNG40bfJCwp3Hd9re0h3nWUjfr+D1lPwwJbs1hUcXauMooK/BAQpCjBKph1MgZHpK8CQ+aP+6
o3E7+CVLElAPVT3rAujkrn2qnkU6EjsQ+Xw84eO5r1+mjCat6vAe0HI/0iRl07c610eqdv4N7dxo
FjJEkGb/ENrldnHHzUyP9Jxe1N7WFXREiCxbRJ5xlGVJAeoXfsZ8sSZiyvD70JQHtwkwX3yLxLh9
rNw2LznGUKzhl+W9fPlCMFTLpQ0aHK/yHq2zzZfMXkultjyiO7taQXzdhJLmtVKvtH9BaN2YujY5
hAn9iuzp3dOZUxiByoLLnPB5xBOR7COErvQuh7Y4vtRpY/6k1dlhXFh7Iy3hDKc0g8fu5M+p80BB
QqK7wW2VdDoNlpEy+RjfWCzIPSEy1GUVJTtJZQgj635XB/oAnvK7JuJA2kxdW8GOw0YDNoK+MoSX
YFkQ7mhMlmKVHeG7CFO7glIG0oD6dH/m42VHC/oGieaQ2lw2EIrlj6WBZiWHjxecgao8gRapCxsn
ox20U8Qf+nqemj3I6BdB5Fnz6wzDFfHN3sjFfHYd/MOqeFypd7JHBri9ZbRqKMcdZeIc4OSxFyp7
HnVj5TLfIbeQpjkcTVivoVN9vXYEFnBZm9sLtKl0qFEX7k1XeL+rWcG7SlY/ZKHede+2VLY9TZSV
UBE/rPgeWEYuy9T4/YZJ6sKgXn9ItNbiuU9lwRXL20+IJpjmz5YbLgevFOBewGv5NEyn+gMLWqGA
c/0ED0B+mIRDW+0kc9eQtQGtnVeYogxQ2nKjbREYDdNEwwgkQB06Ike5S+tuqkuhl6lA8jkJtHwB
1pFaMt/hpkdkhDRbenqhzUs13CS9ZuOdulT8ydfMjbzu9vhW+aCeZqmVQ1JRt/6KsjeVz6hoKsIm
XjttL8FtxxwGvQSWhAGo+5ZmJXhatr0KwNRyYOxqcTbVbCWauP2uMVi5SWG+g/hTeHASsJtsQ6oO
uTSEDxlPtZBLaOQ8RdauSWdm2s5Pj2TNi5Nu200DjK+igyV+ZBwDM9c+Fiz6SeblpF/cuD8Kvwhd
qt3sA/9WF16Z7ZmUR+pvDLFvafYuOxe1NFS1iHo3oMa3rHWEYiXFqCGAg/d8Umz6/VBs6LJMYF3f
uXhSItwI9FvCgscKKFqRA0pdQ9qSZSAUnVTAEeE6lHUmYvscFuOjQLi5q4SNhq7Gyq/FhQh4Q06j
NfH4OLidytWh7CRv8nL2SDmT3okiPipnL+oHQcZVCvhx6SV3D1vEIq96f08uJpR1KO8nMnkHPeXg
7d00Wb063N1cOrWQmK+iPX1r0GhFwrhpk7BXvMrHAoREcC8NbRYG3FHeX3m94fb8UcXxMm7xildy
b+aDIyctIcltKzdC1fyF7CnDSicm7TSvPg3nfK0C928ziQ9u8BY7Pe27t2j9lvbz86VDD3oQGdoe
CDuuwU1JVh6LX80KpSHngOEBElD5Yb4fzhA28x/w/9V66DB2JaO+CeROUXLTxRVjqotsGY7K2uCf
Pxa33AK0WqhF33nwSVIQruCaP1ei9Wc7VqZF/GGKviOVt6Vwn7FJ05c2ZglOmpjCRRjfxxv/Evb8
/SeZw9l982XrStDCMvjMYWnqpfxpgC6wc3Wzf16nx500cEm70LjsGOg+dZW49Z4x08CrRrsDvQVN
3hX6xhCGbAJ4M2qRkttU+okp8OOt/MBS3Wrn8bSpoYL3m1Z6HKjarTcBBPKSU7d7K57PiKz44e6C
i4eYevXf/JKdATUv5ODxnnyzTlonph6yh+YvKeUcskpI8aLjOnehhzuRZ+LqP2v5I+9zIMTLBf34
fpHY1uaiDGQm32l1gNvK322iITfVm5VUF7A2xP3W0zdmWAc3yJL3IHhIwA4duu6sSGQ5pWr1TEma
G0wzGvrCoCVSf+PVumLoU9KrG/2qs0s6szT3R4mgUvBgd+5WZoFVECA39Q5WiJeoTxqPzMJQNU+0
poiiMtw3UYxjNAHZ7y1796iryD5KEv5vi27wf+nqeKK9JciKsz97K8rW8Q+vZXicj/YXAlCh1VQz
aZ1HMWsOrZO3x8uJMFtqsls57eYEx0Ryz/s9lEJOowpYegbfa1rhnmqpOiCIWmUWCu+9JaW6KFpl
XTTPoElDGY27GEB4LacAhVMo0xGmeSvvLMkt08TiVDSoX4kkVAcwrbItZrFnKMDNu8cFHm3r0VMc
QKA7P7frnkP/N0zboa9bSZRcA47JMADOPkAeYQ3sxxx71lRU55XyN+psX8htQ/tGgmBMoYlCFWMS
KtibM1sP+PSydzViyB8O2CruirsCgYCSlpOF3V7C7DAX4BEzvl/rec2qeFOGNrGf02c+4UElVPcO
mB38MhVHH8Qv5/bF3gMKgws5i08QtnKbZsInH8j1+RBD3Ed38IWq2kks7KSdmCREa8sMeB67/jQP
H5+WjIZK71T8YnznSg+12hN+otuLnVCqJRPoFozT0Tgjn7iM4UwbK/fuq2pllcpG/OFawerVBt7F
HiOpKDO7T8NFt/KuidjCF+/QxdI7kGDXpvG+t/wl6T5dnwUNUzPQPrgfdY9emCGdbDObWHTneMgl
swE6UeuMtsri3N1S1tJUz9zUZkfY0czFyc1clpVUi8qSPJJx2gTKuXbOIxM2aZxMHopHI1ZU4Et8
9NPzbAv3ooEvS6zlUK1O35KKephwPWffYJcS2n4jiVDAQGzTu6u101bDTcvEoX4n4TYWqhGS638A
a1uSJd8uXykHgnPZ17RhgPLUvJafIedqei4P5xWT8+fkcSyAXBtnsi3Ey7Us14syJEgakVPdYD85
ijh0xt6TINJWCm1TEzP5p8H5JhoA5f5/NzFHC4g/oRM1vDr4XRxkn664MPp3U1lmHqrw17nc+bee
FYJvZ3/DxcTsp7TTY98pxAuH6FE9hyNTr8+n8xn6WQqXFAjpYFmMZQV/Wn45KuBY2fsRUIJvOWy4
mN/StJWOwUdwdLCOh8dlnsxkwjWiblu7C4TcFMIJXvLqaJcUVA8lLYJlnMapiaOZPI+QNF+PhBaK
K7LHw2R2isL9EBsU6H1c3tpZ8VSfgtR0wOWR8xphUD4MfYegEKrRQ0fFMNZY+1r8jJgEXLTSJfUW
GqEJbpordRx1bi461zvxHnPNM5nvHvGE3N7/R7lbFwonUiGr5htez7hWqSOwD5S8wlv6Ij4VY1Oz
xK632DXYKxhOakVu9yxUJBVdtPRzylHWWtg6yBDZg2U0xRXx8xx5gn3wqkf0glB77ecKz0QtpDyq
y5gGbffDSwKVmaKi4RM7T2yQ16CsuJMGmV7yPz8adKkTF1+Eg3GAIjhgDNrlFmS2HTZR5YiWajKC
UYth6d1Iu7xA7HOVRC+xjYZ8Q7eiddpPnrtECThhFdjQvNDcb9754Akr+XRiIDwqXKSo185lCOng
IeMBl2MmnqgPQRDtbQoWVQb5vwvhroScSnm+iUS/PeRT7lJjpRdtxjwDu9tRjfXzi91BKYMChT9H
cW8TIqlMG3dGGCITLg7tCzWqP5ktMV3kMwIRrgia6WLOD/tJ7oT3exxEq/2JrxaoSyxul4wW61IC
J9ajIQCnhVVR6kvPEKewGVYNOWuLREXWmhOJj3Ca1G0zhZgCLSyBSps5RHXasIDuj5J/Z2+ZFusb
7BaoxkXSx72dDosCpyWW1BDd8Ak9xyio2yf6/sOk8GINoRHiEXOGyxKdC9F23UW+s2y98ofNKngY
Q/ZcwIUQXZ/wA0+XI7xKodVJlp+h9niHLdZsCzAVQAkQtmnfBAuYtUFKiYYhGABTf/dyk9AFJci9
+eOOc7CsI7GMAzZalmyfTUqVxiVK+xYk+mqRxwaWnHsfOFwBF5hRuXsTa8U7p5t570Yklx/Abxhy
cbgz81yyh7MnbtkwLpz7M/43nMFPwmqOKOo+mHDZcrC/uEltcWB3fjPBcUfKPuKjlsS07pzSLOWZ
/gHiytXasXeJkFmRIf2ug9DWl6Y9oLETpJKOqgB0DBL5x02ESmZvFb1vPHdtKupo0X8PZdSR1Evi
hnW6XxfWPHM57o7ohHx5sleA76i4NbnMnHCndJZI24rfongTVCwZCsB5GGiATOYNH1wxHVUuM88c
7y+DLlmBXW4vK4VHEhUG+kS338FPN52E+rl4mSgCh28UmsgmumnFnYfFFr1C4uYE2qLTFgFS4vvw
DsZlvlr3W9zXT+8zZGuqmeZhtOa5NyO+1VeQsPpady8c/g7Me0TU2QkK6S+TaBh6oUfxd4XHKomp
QyCV9uryqlGISHoWYGTxiKiS20nPoRpiFYmN2hhcVnkTTOKP4/E5U1upiHXnZ54MrJZtRvJy+/U+
UhEXZcY883JxnbxOA9B/1YjxcMqDjXH29W0x8/RmNKyu+Z0j9d+OoOB04IwIFYDSDvz63L3tQAwn
/OZu/BelZQW8sPRT0z7e3wc0BwT2m5CLQQPs/nBNFltGXegcZeEZ0KEbBZh+p5UxkckAo07wl7gF
AnQwRHrONy8dLPeG8eTThZQaNIRMsb+sZIzeTiO1QhhGyGJHSIartvSMsjDX9KnQsUWrmqn3j7Ma
D2lJOINHdGY6Tx7QP0qCrAeWtmCfxzdCfLIso6HHX8TESRZKJhU45XlV8+oqLXnqEx2ttyRn28JY
zH/J02fz9ng5/k7B8JjvcTf7j46J37mtOzSHKr4D5K2qvnvExSvuHgp3AZXjR+cq7ffuu0UP2OWv
RFxwSrgA4LnV/1kny/BPxq0mC9xRbL8BkAQZS3EpnQHdKNh0Tg9/pLiqEwFcPINtBvJev9KS8to0
QVk89wqKvxYw8470EFHc/SD37A2uYs3chwCunZ2HRPwePMQ/lQK8ZQ4YHMh1CW6pfGXSiXpBAFq1
VYl+NuUqRtVRiA4q9wZkAm4tm95+za2sdRS1yq/AY5X/3TMgxI/sLz28KDyb9BjTWnKnqiwxwslX
kVUQIbjGHsoRC6Gvlam4KJe8tWJBMZGhUS0fnVuT6ke9IsMm1GKpO7qZ53Og5Wr3yCX1qr+K38rC
HSMus5pdCl0CCXt21LisKkwABs6mnfhZE9OXoHx9c894tbj9vFV+TmfvA50FvRf5+Xd3FVOVpHnz
zw80O45xjBdCaebLez16G+Hot7XzsiP3Ay73II8cz8pYER/DS3/U8w7+DkLrQG5wzs2aWRaixAbU
2WP6Vg3JiZrZQj0A9gCya5I/P1hREb4D2N1BEVI8eRrQbABCFsHReJ+xnuVmkNFbvJaJqg4DOpAQ
cTL5We1tw++sytnB9DUks0KhQ6xSt0ciz8yVC7d4HJwVxCKtWhD0f1WGEGvI0EWD1n728qgsl2TB
WtD+vptrPBFHOZs5a0QPoaKhOEiu0mXQJfITvkv3091gr2J0Oyb3GSOoWRCfBWFT55DFISr9EWne
vkP8f9/E2SFXelQYxaE6prCne5jGvf370daRZV6HgOFdxJNVaObsVlCatlHouC15m8xND0/iTA0W
Sz6+7AbMr4y85r8WTep6+3OJt1EMV+HPvzD10VbJccFimP1z13u1gpht9ghVx8MeAndyLBJdg5Oy
pN3faDrFyidQoI8Pi4LAVTCo1NXPTrRdIPBl6NrNl4zOEQ57sjIRlEzH/tb3R9GSwXpHlEPBuK25
1oY34EP6zkHDHLEjMkqV1sMJOr/49WS6rmX3IREo/y8raN6YTKPYN1F6EUeFCWAsBKR+ADsR0Tv8
j0s+tqlPPripM5ryBQP4uu2cRXj/TQPpeBUCgNz66vkgq9cZ1E65UyWNkFmF0VYna/MKhT+NU1sN
lvVfLp2k0YdPVp+2xkiiPMzpaD8U+G5pLNEUiBIlj8c30g+s+oPHJ4XGRTRYx/+op/RxTRNAFGX6
IVizdgREDVOHKFc2bz2svy+mzPyrJJoF4MDgFnBz59quU+hM99CMMj/f+eV/Iv74cmxfMqFE1dYO
M7Z57Pll9c08iUwdK/VwypaQbAQLx6BLntDnALf+U0B1yZbb7s4w8lmvdIPmpb5WZFISRySLz2DT
DcpKR7cIlRJsJBCVcpYQyP4MHWKgUDz2lgdWMThNUGP1Mda2brnDJy9BX6uZ7DMm4kiz//LD2NKx
BuP6paKNApp77e1oe9uvN94rZgf8k730eBkXoxC8w+PiCuhFTCsard1PgVNY1Wc03hndFa5oSLYj
q/oAKhX8G3pidFT2YJCcDyVi3/5vzZIvHKw0A4w6a8kvIrb+Z/iwg/QJLA1b088bvnOhOVBoM1sI
MRRSzpP6dbZrJldBoaFq9rfSHL2EX+kHBN6glgX7qsaeLejKubzBFdCrgaHVJtMDoZQKd6i8GwU3
4JdqeKEFkeG54FU10b8JBEnI4/4+B+rIYgYkVCkMffomEs2EkFJKU9V1e4vCgDhz+RgDDiirITCB
tRzmo46D1/OYb/GFTkyUxfQnFIV72N9eKIiKGEVVa9nOzMjPniPSyI/LLFQZbQKxLZN3NFoib1GV
JV6o2XFArYZ+1Ipei0usKRZ64GJWJ8Hutv2wu+N4QP+sd5y2K4LtHk5t2o1sOBuylCaZrVW7QeZ2
EFsl1dcFvQ/tp8LVIsjFSGOXFVcBJ8P6fyQ8M+SD2hSgPz7Qeaq7K/h3CfmhaYka5dZ6nbEJMDXi
zOsxG0Umbs1KxnD1TcpPld+L2vTKmdFZr2M27Y8gZz2IlJZPtUVm9HH8M1jSqut5Bp66cvUv5ssF
Suh550Umnb9t1Y9viB3zrHy2wBTzkeJW5d5EaJXdQXGXFBT+0YYZ4Tjm+u6IQwMHJ75lySg0+g3V
ls17aNbSMANXSwxV/ABmxAEZYcI4Cxe/6FmCgnsfMAoI6SLEYP561PIaq0n//LeONG7naIYtZ21c
uhPxgp7aNGl8wW9Tcx7HD1Ry3JnCnnHtPG/bjnX2IzgWjCSlVGnn28HHN9lCpuu18F+OAjCubamr
eYNoFKnc4c8qf1IHYXci4rtyE9/WE3VmckyyA5j7y9skYu2UYDKja5L3LcQGsSwEy2jisNvgigCw
UDqoacsFjzacmaUnu9FcRJHLSKXFKfjKXME1sysH0YNvA1U8y8t/kTuE9dobAaiS13HPhTuj+Z+K
V91buogqC4CCPTIPtNZ9OaJMmZcsoR1RqY0kAqC6F7mrFr+ERKe2uPCw6ziLdZPAfBKV/P/ZuIv5
Bpd8/VYML8+30LfIK2QxIrljnaPo+FHs1GSGOHhL5X+81mdvINCGhncj4UErLYqgJC3OFYpozEsY
9QgUncqquglGnLwXM6EynTSUaeWqZC7AmJdm41gwVGN1T3zrRPu5lbNDeE8/7DVoc96Th1I/bUh7
RwcdVNeemrM7zPs58+Ikr7X6EFrlc1oTIM34NpjPPt3OKE7gyj5z/zwu76bvz/9Te9Gvver4VoN9
96wlw9wgJHAY9sz0lUZIBrB46Fd2sJj6cR0E8cHigKVVbSrHZMGYYN1JANBflFPnMa05vnPjCVhW
lgaeOocSqUAfhrBNg1jv1V0ARRilGeNaPrcnfr1zs1AYOgD/JRaNm1uSRpPqzE9can4r6JHBRm3H
weeM28nAWzp7pnTpb9wpI6uXB/HR0UJp2Upq3kyO4d+rQiGkctm+5XuS+fci+9ceq8urqr0JwTOa
wvq/KV640MfOAsr2sQDHZ+RzxL4iNf6aJVwHCJeumf8j2UcNsPkf3hw6if4NXmliEziieuSxNfDv
Jn6bCY3AbMYbWH7gIWBAdrBP8ygdTWYuSvIQZt7JjlYMXJ5in08BhN/kW61Z4KShT4bsUuSjMCvC
lYN0E+UXiz+MESjfbSVXCVTtLiC/Wy/0FmNji2E4F4R56k4eym4BcVyV+QfO+PffzYxDhprXHgJP
6xRxgQDhjXVV62s7D6Onf819L8ewC/YgIH8+Y20CKDI+y4XRHTv3hfS+XU3yWfxTGu1XuTYci/27
Id/+vGY4T2bTu0BiobDZU9cVLpDzvET6qtiTBuVFk4877bJVvenW+wv13OocDZOqoGjt+PD8QJkl
edemJQ7GVOF2oiYv6LnKP8pUfZT78Rs9I0d9VIjX7XmhUvElWusz7rsSw13g1yIDxZJc4Qfzm92i
r1fM7lL48rYHXDlIwN1eCrhbu5M6kCy4B5rpj9Nn3cQ19iYRgW43UNyr4QPLIKHZsTY9XKjnrO/I
dT69a/RK3R0JKJNPGfv7lfNDxVLhjiTugqqEzIvIoGET1qYY8y/szz5Tq5cxD09FJKUA6rCZ0k3Y
Yb2cT2LbQ/ImYkAoOZzVdelq0luF9zqfgDg56rx0n9bdu3no9l01lpOd3I9RdefbUaSNSWpqacSf
xk/iVck1bLIvX61rnx2HGob/4m9hmZCTcAkcyokZCVkFCci3ZZlBTGSzLZoxpoDjsUlPYEHYCBas
hW+23rWF8YOT4ZmXySADDRmFm8fLAGnOZA7Ifwm5JS0hlFBgy+cyoMbiRDSEcRoY34ID9yfd4Jlu
6q3za5K0kgES/FggjLAYD6liiOisDvOvc7TF0btfx7+2wQ/lnFMQix1XwRb2nz+Kj1lsiAygbQ6Q
v8+dMnQmBcPlgeZVsFh/O8oCdDZ+Xxom2+Bo7Yu0DOUH9ng7WgZ1qXOyMhqHYn1v7nmMZxaraaIq
tvme+NWltm+3FO8bWW4hMwQZOnwSUedoaA/KxIh+z1AvOQRGdM9lFzQLvwwAhqDqQ1eagvRI8Hnl
bf4zcbpVIpc+lXDIG9DPE+5GaLoHfAXmYhmLjU+UgJGqfSt8axljX9jDjE593jHKre/OS6bSz1hk
Z0sm3V+cc1q2RWuuUSe/UdT1GG0AJSkqCM4/GVkUEXJhaD6GCimrUiK/0KWytGYAVJCQAWEQMkqR
f/RJS78EKa+tIagrdk6IGdX1DuGTgk7LW8OrPL4FxismpIg5wSXzxH9Amd4N4Leyaf164DQlaJdC
MT0hjnoxRDq3kfk0TLIE0niTm+QiBuAuJCK0WbJar2lDu8lYUz852uBLNwcB5HAkJz8cbVAzIMF7
hzuJcLgZ6JCNyvRWIX0GcYQLY2GEQhsO+uss+ckNHmISDHdrSpw0lyK1Ki9CpZAkHvVnYaAWdUl+
7IKmItgKL3CxcBG0sE0T7I9h5dysi0bQmJ1E2EXzTsLZxZyqWpy/y40t5AIDEE5Hhn5dSd9lMYlV
IYY/Vq7HboUCF3eSy8HPM9DuaaNjWAWzfBUQAnk3yinHPkK9PqHa773TC1/38ISDbTJglSEZYvha
DMQ9YNT/zTn7jExikzn0lbsv9V3kpGcUMSZclZU1+6N5hrnIoMmFjWCsjhe0QeLvd2US77miDRmq
mCERYbkUanTOh1q14/gDtkg//saSiXWS2InoNJRW6rBw724JWtROROoWR+lVIolM+u/S+Sg/S8hC
Pxw7PbSjOKXnhqitsc4DAaf4z1PUE7AMRKoXeylNyKr6ftgmtNjGJGZ8qu6/VC0RaocGpMM7PNKR
QG6EPVFbZqOcBqx7gz6vNhmXWK4auSKjs64+mIHzOa+m1KOivOjBbnQV/oSiLHCB5VsfAkYqwBio
Y47A1UoA/mnJATahecvGyzNA++9s/e6a8PzYHTm5d3/4gw9bf4WMK/A13uhbxyWRBUsDpDVkADDB
c6QWz0gTrpKlKX0pYJPVBaPi7YbVrRLuI0XHTmx3m7maJ2XIpeE78JY0kZM78VdmDcY9zWkaDhBX
wSmA2hfeMxMozmZGAJAalVHm6Oc4seF52R70IJjnPN9k9i87sMHgoaxrcm7T6Zl00mK+X9fFys1A
2SmBNOXB6zssZWTpfOER0jKZOBRjNKrmLfe2dBYkiQuDz5u4l5YuQe6CvH3eLWPnCJ3BoYjuR0Fe
vDG7U+OQI2qfxCMLzyJgWQl6g2dbydm+V1xswOfMdXnumwb2ZwThdqrmrptm747ZMUf/KKzKbxcw
F7qmSD2IvzGtyWk568vJDgK0w7kXdH4qhqO8yxuyJVnBijWafmB+4XKcuI4XyMVlvDLAJX3RSKmc
HBRarYWpZfvqyriENgnq/DCYazV1AJ3U8ru5hi9nRdwaEcfduXTPDiQLpQyCgfYv1ThG0lZvprQd
k79VEm9FU9Khs+2pyNX80WpjC8LZ0Wn6qgmLdv06p9BOQiQ7HGV3pEyXOPF/0CJI0YpKffjISS/A
et4wQpBSHQ0A5+TRSWzb+EW33npk0cDEWYapL8dHy/VsDEUjqg+Y08xAQqwErm2KGFTQLp8poHYl
gA+swMv24x0MQa5YDYAZw9eJWnxIJRysAPlq7NSZDbt3sXEm6ZpDacdKGr11faH/HnrS7OiKeEwo
2bERIn9DQIldmfn7JH8DXuNEpJDpfiEbhNoR+XgVbk9llgChAdYfZr89l9YtsMXFHm7gIJ87R5w9
dHv9e+oAvVWPkoBdRyxyF5kqLwsv8nBXKoxZkgdx9cEyieu4Gu/feKbCrgINMPuRJBzrir+E5Pre
jKkIGGFOZ/IdKPxavtOHuM0duOFhEA183Mcq6LXKDewCqmw8bSSrwoH5Jxla5coL/p2NQnFsR//v
rqVrVl7YHTnwaAd3q6uVDPtpQidVM4vV3iOTba/YYQFcWY+BeC27xRUo46uE2pLS7zRome7svBcY
cyupk4CvjIZDZz9GNm9xCXppt9sNmXOGi+bmNKOyV96PP2T3npTdKgKnD0fTsWJ8Epc80vitcX4r
si8uZKL0W0LpTg8FiZzW0Jtw1E5SjHBCyaftbBblB+3s8Xcl2PSVq4UheDPap2cOoYcirCYJEfN1
7L47KbjscR7X7L38rVqklp2iRBHbmtNSOupcnTAOvST98WZfQwlgqfjcHjnGnVR/NXLFEL5ecktB
m4dttVynyYJGAqp2zYau7IjCBuqbXlr9/GR32ljNX1wSmmzSCeCzqxTFU1byoJaY8qH2y99+3+2E
jMQJ1/7Vc705QhTHbsrF6LMl5ydOD9uyGNPKM0V9dW/lDg/dXNTD7wIvvuFUXZUkN9MwNgfwqXJ2
0f71KNWrHmLms5PL3LfnRZgJaq4GPOvWD/hQ5dpUA6ei831mwD2zm2GWz1BtpdRtKW1mbRtg/Tx1
vjUOVT5Lq0XSFxNih6y5+y399J8c0Gjggso+iDaOsQsRoxC70jU6bSmE8OAUsb3tA2ZFQuY76mwJ
Eq0LTJ/8HpxIWss0ANHLsw0WiXgiZqxZwjgSi5mzW/sfukf3t78HVvdXUR91mCZ2tYR3hTdaxBfc
l1u6TyKqDDdvOD7OIPsQxDQnxb3rqARraZmNzRsTAtFqEGAi4f1f9aF6/6l7x/v/PuCBWurL1HbK
YI+XnIpjoDIx3sWtNolDtJwBsG0kcRGLL6e/kvWDy3Ds3rXbt/RAG1nICFoGDjPZe77izV9iAfKu
dOGq/c7NASVNMCqsVqWhP6I6Xi79EC2qeVR6xR5H0Luk5skhRusZdn4V1uI+PGMomlKMIPuieudo
AZHeBjtyuAgJC2f3fZOf4dwjj5+6Jgjmek+Pv3e55qSZi0pM28kZUG342M1/Cf0EStgSE/uXcb3f
vKeKdEpsjJwDhzTuqQbIUra87bD/X6KgHpvl7WEyg2FuVnRyDrkoxP3SlLLhGpqq6vgyXM0XLr0p
rBKdp7D4eD5IUfaZHoj9zUPQRYn7QCBxmJs2u3Szl/fFQ3hzgM3s3w1yjaFdr2s6O56Su4Mjm4AD
Pm2Hh+U3GtrEiQvtXc3O1wOBDBSzLdL9Qv2R4OTcGuACi0ixihj5EmOaIzFONr0CXWLltqnVn47D
0wvlPRV5MMyQHxF88Gdaz4swVag5TlW6HjY1/3FTgWtqDu3SP8pOn5eMzAo6tCZ4uLfafSFXu2Ut
W30jNixK4gab49VSASGoxBpMVlq9DI2GY/XuowtRV70/IYgskLvWQPDYS+HzVEc54vOLS2rdQV6s
Nd8S7VAVdXTeyVTGSQi90QFVrhcHZCIzSxuSSb75Cbpec+eYWye8B6SmApC3bT23FUC2V4wtKCnM
UNDLx293DsfJk+Cv4E2FtpQHIg9KwCg5ENKBt4qeY+AfT9IpWxKUtNkSrHouPJxpo0Iw0LBNf6ai
JUJ9dKiDmhIjt803P75eUr1Lmhh4hgnxVam3YIxiCFX7k59NOoQqoUt71PP9EX07/ww1ot9JUGfl
agw+6SlnsjIm5x7mjdXM6j7+F7fMCeA5HG9u9Ff4f2w+4q4EB5qOIsSEaTdmjft2FEirBnTqE5Z2
4LwmQcEhWUlYwH5ClHLNWx63BRgDKQSQ9zrCxTZf3BmHCAxppmGomrJH0dpMPpGk/iaIPW2SaHyn
ChX7rWKLyS5HO7G8jcrxwkPyD2s8mbGpgsGAG/RxVQDp7HrpUnjrfuv17USYqg4RDSozJF1KK90b
4zFCFxUAe69pTrqupydkDB5U2fgBK8wJi7YflAe5/QyXj75f+7t01E4HzIVuld8nZjBTG9djbv37
nfC29wEbwG/p2Swh2avI+ONrVnslrCmwTQrteXJmRamSYpvZSNAqYeCOAlgnpBmFpyJJrcORRvk9
cOZjgRQ+bjh05wecg3aEmmJvaRI3J+9SOzMM4j/bNvFxZQLqB+pe4+39fPL0sn2QHQJ26mll/B+d
ZXckW/j1zQ4KLnwhObQGj8LStYBJ83YFo7HUkk+ZEh1R6yiAWqnf7o81yimgvlFtvKxmgxpQ4grZ
Hfmz2hvfvcBTzFtNcOzPiHSJtu4VdW/aF436lRPpFw406q/6PAvg8wWef+RYrw7EWqb/xYNTgLOr
CtybPJn6j9fkn9VuBKprcNAZdL4KgxlLRwacEbNVRgNsYA3Uf4EhjCIUEoMfSeaZeS7F7HLXPFuU
c2B/vRyQ5EjU1rR0p1KN49g9P7LkxY5ssOr8VBjtgzrqh2Ft4KxDcsziSd04v5M7RxyjgjESU+5e
TR+Ex9oLa9EhMkoFmfxHat1iU0Tb9uXZreNWYGvMPYMb+Ru2AKPi+f7REMqJ6hUEC28s12xKToLl
zakqLilJEO+3wQI90OuGFLTcZeOS741W8YAcEpg174ewFHy25LmAuGy8up5DX/LtQjVNfK8Wladi
TFRdS0UmlBu0p0YDgp3ia6g5Wyber6HQMX3zViapPP1KRii1Oh+jGS4Md60OfoPpFPdHQKaxOCo4
XpJ//H9PdOjb6nFft695CLLb8gnt5vJXoNFFFO8M+SYMk8ff9ZzVy8vdAAXOSbJ3TJXhUC3Y9wbn
yLAwRMHTdxjnGoD2usYQR+i2Hi7oXsHWkJYstf+Xr7PSodrkodokFfggm27lEpMlz+pfTmOxC3mf
aVz6w2pqwzQTW3Qwlulre11IRi+IM3eWTgQbeGUhG1fBeJacRAXUPppa6U9f2loFl8hKaVE7WYib
iv7myWNTVmWXMNfeERWUL9oEJw1J1btuRYpBL6p+FzoTnaeMMql4dWrYPwHC+nY7C/LzgbJcZr25
aA4w6JmH7gR8EhTK6dOGwm082igMmRaEaKG8TsZe/DI9tGwABEIZLBz2VDO/q7wOLmlGxDJe/QcT
rOam7W5pVKt6InsX+kILPX4/VKO/94jxSepX7JdVXroNteYmH6/OWilfaE6gjGhQEuf4NxkpSL7h
SgGuYnAf+sx5sa1Jilt38R7C7dbvPiRC0pIcE7vuvLmkzrC1+eldX6vB18RoK2/1/oq64PGpw0Fz
FIUIHGCuHBvyTdyF+qa4mI/+0cXKYM7ddD1ZZny/azSMOYlZd+zxHmVuEUj92YXYq4DUEcq/oOzE
Q15XzcW6iN1nKLu43ZB0Q5QkhqO9+BH136OKB+rZyy4dtDigyAKqEqqUXzq17amHTZqj9QKM+idq
xjRRz4FyCR4aa6HNOQBajedrFp3Tw9yXNzpxzD5Y8Qal1Y9XKVkZnqZEi+wNWDkRxSVHoy4qN9eW
PjMB+RHwqq8ibwil8W0la8zh5Sn5UxUsJo0x0aIjnFpwEL+yA/eB7kF+RenEkYNIxqRny9dJFnPV
ehp0glzY+rrNq09fUvuWczNTdH3HDlIQHiHhfz/IWtcVeaw4UVvKok+NqQ3ohAISrejL0dwtdiaW
ajJn9qP2z8O2r/003p2MG1tjlEPAHYFs+7FUcnwTX0Red1/+ZCBLfJ53I/fvNu8oua7eoTWoj3RN
38eIE6fq8TqE1LZNE08qHBWVm67Ufvhch+1M76sJsSnbzIRAGdCFqRreU5RXYCQWz2OAu1NIvBIB
bA9xrX7mykvOzw2DGdknMMnJlYL1VnTaf9vsRe0dtsbX4Qn8CfEFeNAnx1nRVSmM6KL4zSYiDOlI
1w6R0KfG6EotMyZiQTKGc78tlngrU3jWA+Ix9qAfXahslmRZvrJJUddd/oVVMoHslZkVfM36mZAW
ov4egGQ3NkxpdOxyY0i5a89CDY3PCvV7M/hPX+zxDjzKIRn4n/wLkKrS4g/gl855IimrHkhy3mXp
YHYaiLwGpQKp3/oMCpdoxWItG6XY2yIWOoq2PL7EttkoY5kyJ1vKm8t3JYW4PtJADLZy1cfbVHLN
QEJX8tXfttIcfI+D/xSFQf/7vHBZeD8DpSouWWfByPjyBRRZWa2cC5pfOH4Pl3Uj3+zqMY2VX2Lk
5ikYRu1o2Zx56GLOG49ouP/E9d1h98s7lHyA7YDhli0mHUmNIY0ofSZ5EljKz5SSmSYtpPT6MqRc
rdyGMyJ6KE4teoXKSIC5FSh2HHaDFFL8V/l70i2kmQr7VQBVD3uP8GRhTSEFTDfFUMCj9N5vwSQd
AcwtpUj5UqYrx/GTuz4zON+cHcQid198hJBsmncUKwyLLFtsHKZo00rTveT6oV5jh+IIJx7R2JxN
1/UgGYrDR926pbcx6td33t1/B5oMkwGvfWtl+KTi2SceB2ruJlDRzivl8XOmz/EjszfkuEwAkEsr
7nI7a1wa7Wc9F/VLh7DH+6gQm44StV71U6Oe798HESiPQrDTXyfGGIH3KNi9gr30xmBr//qQbwGm
MX4biW3HqaDUveIJYi60fuSkoCMMcxmeAmj3HQv/JEIUX+V/82bzbTgn3vu36h+4D81hxN42Y4bf
/mfWyoDsKT6vDKv6YunsXIhT38zLsO03rGJzZSXbxksdwJR35IB+RJASzUOMBueZx3YCFHU+N1gu
/yKG7I/nOza04xvMZY00IgMRh6lNqR5yrrN/HanTCS69E9lGeKqFzbzGxPTTMZiksXVlZpYNL7LU
4WGVC/FjaElkbqsW4nGq4ZmJlv+kKY6NPlxgRY4sMqCBj7aDcML+ins3oMH7LnKFAcsBV0UMnjjt
oSigmgf/WiqRvLWXriozijXi3p8xt6vBSSZQRYi2f28GlZQ+SOJlFwO91zM5R1wsqYxpwCHHOfW2
HlJDm4ze6bwoRVPOpg9DpI/IU+kG2MlNDZsC9yB4/XgA0xoKdCddshpxUVq6PXZYgwmajPEeQbW3
a8Km3IegiV1qsXl0MBWvUVg0dIQ1i9H9PIa6SrVhVz5tq7laMxkMcD6ZSV3AKtcLnH1Eyt2YcDrK
3dRkWXRj4W1vwXO/Gj3bfPtecGts9nq9+3ljRzzNGpRu4mA/sRAPpAXFT4ug8I4DAPqgzuV5Q2Uf
Sj/5uEHSQXXjDR6pmhomIGZ2XCKsp3pKLnvclDP29D3ctuZrHRnWT5L9Tjyg61PCsIBchoEaq1YA
LVXfgZCOAUmhiOoiZo+cdQgrJYbkelt/870NlgDYJh5P9q2f2thnkvT93Xtvzh/l5UWCTK+oST1s
OcoNqFbqKg5l6gRY+sa55OZwlfs6mjFr9QQqMYIRgw5jFWKBy48QMor/StwBbrEe2qmJ0OkaZZEj
rjkEWfhubxXrnUGzKm8De19FD0Pd8hiYbWOx/ZXQR2FxKPcUeAWwYcRGKfH875+gyB6eY0VVjiG1
aSVwTyn69lB0aB+PCG0MSmTbwlhvf2Lqbhpw6YVnz8sURosLeuvnAG9UJUhA8bEgBbk3qbbjRd9l
5cn0MVtvCQxwG5upmvi2sXIqHV+lb4O41V24eOkvB6sI+cMx+FprxGkryaAHmgXYw4/aAQBEBhNq
gZQHyg0jsQ3nI4qV0bqhUevQgKsgvHNxCtNMcEGVPx3cHPme3Nss/p425A5I5s9VgXBrqDULGmBJ
qlK/cChZqClUnDkRFWxU03fIYhnuXjveFrYuuC07n2lRDG3YLQBjp3c4EWTybbt37hRWERbYnbi7
FwA8s+iQslAX7V6fkyFNdsPjXJNQ1lVWa2Uo4eGL/Kd26xRTNedZjiUQt5vhrG+gCyVQqFqofGWr
63pkxPGjsDIdEF+tkm1b5N6FOYr2yJb40fRjftNjDyHXQnVnZErJooUXoY26Zo1BPTxt1OY8nxpf
7l2eYXoaoPscR99bYG09Nh5QOrocFSqloKMUiQDhyKqsCkVzx9i5m45YVZUHz0WGQkadisU7Ec0i
avN9/yyWFL4gNZ0LVfhbf1oeB0vRBUTuUe6hZfqdWh2fsZTtcLZIQxmKOkLsqQLKVoWUPxjH74AM
kqmnlpgNpCv8005JPiMuN3B0UNMoV0jpT6G8+iH+0C/hZnGOxDE1j7ZUNNSv1ypc8l2QkMDZ0Zbv
hn7vtdLhu5mJkFRMepoM3+b/0uEUrhPamLaDcbRiKayE8fWsUEb7GrquAR/2Pd2T8IdM/EcBmWgF
BiQdGjdEY/njTYjPNqPt4fQKWoiXSWoReY5tGyy+9iMRehczHXZGhz9sEq0MYaexEGoKVWayvZ5b
lchadoAt6Qds6U1PNoFB5nFT9RmKL0RluODI3CB5h8CRUjtxmsNUX0Y3MzV+wL58phPidllrykqN
GqEhPUmttwwBbcy8mF5le02DhGmN80OOIrvdPbXGaAFc4Tj3cFXEHHbKfE624WjpmXqMHGHRsAPR
/zMpEL6SJiTq4Zi3SmRm6xr0S0CV3nOoGx48SiViSuvzeQynO/jeSZoNdV/uwLb/ELMVLNWIcz5L
//bvfrgMbIv0tDAZGdlCpveR41X2pZkfA8t0F0sAmrx8BY976wfEF1O21p7/2T8AA/OgVx6l6zDF
nPrsgqsm2ppTKc581ujgMDmDSdsM6cT5xupaglx48U10hCk0v3tFM4Xd1UnlPYYvE7yKBpMyVx8/
abELOZ8akCarIglfWnefAjk4l4tSykPB/sId+aWw8uX1hHl+tS8tx3qHG5QWYgPA9wIUjGzC4oB4
xxV1efmmqusFd5R4LEDXf4qPOPXSFQikaJzO8PL85aFyM6I1jV46nfID7wf7+j2fq17np+YpXbMq
jD95Gcx9Nd05TfzkZWawGF1ILFpZME4khq2TnVGZE4wQPP9jQrnkRf3iJ4GEZblGi16D/Xhupk+7
hJ93j8A4i/ignSuMRnPdOl1QphTnItSDhEqN0duer30kXvSUI1B4q0nEHC3JgxLSpEGOZX2jrtTe
u6JPvpS/mY4BAm3eksP0iQ+xyUw4PRUQ8/+3ZsBSaSxkZJzoXjJmBCJQdjp5sACE4QexNRukJQWf
KFLjfm/p4lk3Tc5vdziToxiJaL5usVV7pCfGXsL67vKbpHhSJUHL13lxqiXPqez+UsPWU7zPrayA
1MD5sV0vokauKP0xw2Tn/Dxik2VjEcFSlFnaBqG2nt523q4rjxpyhwUfNbxaKII/iWyS7K3l3nwf
BKzXzNZ5/v/9IyQ+DQkwlzTM9I1dXBtsSWkEDdUpCpETLT6XAwP0kZD2GdSYM6CHSVs4tmidMmP5
n9qUDro1qWZmq8IkjGxbeUq1bSv9b2I5phj0c9ZSlkzXGTXdNjq8yoNNNvzLRiNboJjRKT9FQrXD
V/55fdQsdSHoclEKsYFK9bF4beLU5FIaFsS6wwtw92txq48zgtyANkbwc5v0Of5EiQvyKdPoLrsJ
X9Td3LL9gfTjAiPotF9Ng9G/ec/ehuV/uYzucRuuDe4rdgyP1BMdV0/tjCdvlkfjuLsNdo2h1Fpv
LcF0bg8Z4BjOJ1nD8OF3DvGQRvYI1d0uk14/oFah8SJXkcyIy+KbUtbWi8Lbedc46q7y/jgHkHFx
ufAcrTNVMckC+aRVDdhMhL4uBwdA3NlqDMMn7XEPyWjwG3n6OQ8gP2zKVPHBysSQjo7Gj4ipudOL
cb8KrJbdzzcgjaAL3do8jjXdzJ1hmTnxgQ+VyKnDmUL+NrpBJECZKYNxWLEdmR0rUdRmaR23DBvw
iyCtzKHgk1281zdlxdsly211ACih5a1DaR9sEfeVi0Gx/yFjYWS0HPnQLULkCx68uLg34G9G6GOb
M9iFw9F2LYkh8Dg6ykUy22wLIv3LDPS5Irmnly/d65N8lIcYb4GvSITCVYO6ON+xsJuSN10ZKotH
daAOFrjEj84azCvzeanW66d8BuG5SY6KjCyQpbUWpEHMpedjjBZz86TfYDo963at6+A3nfaHYppO
HfNYSEP0/MJ8RazARdUAwYNp/Z5K2KaUGSK0bO0cguaGC5bn/0KnaTHSBTVrFLTaDjDYBKceFj+0
JOyg+bugG480S4UvT5dKz1HD8W17A1B0xVIq0O5uLmtFBwdxdNG7auVz5r94gXHISQHI3OeqUpWB
xrBLyDwppuis+vhZ4wc5vu+IMuqHNpwe3DhiW5W8Ob4D4dCxnAdWFW7E1weFaYso59R0Q6USIk3A
LHszZiL3SABBUY+RwjG6xWvuz74FYmiv4pYj07qpLZSEm6fgbcwAfhB8RMQT258MCkt+5+aB/NLZ
AOgUJmnifcp180v9TaYwwmeNPDkGwGxo8w360AG2qXLVEd/PMLLuVzDCR/qyK0+0KP0LHk0/74de
jR9LiS99U0c8aiXwATFxZju8Zy5pvAMqs+gI7zcsTHf/+WLbOiAegS1BwrlLiLyjbjZg+aCLQfEi
2POlZwpdYmilyXBCYWk+S3Z4DZ/GoUBOvNzOPsOZPEqIZUKGZbnUFj7zeOWqHhjGhnDMp5upe5ja
/YKcTss49gDhVBiD3yxPWu6a4oJJn3tnn7Yner3QREhi8yuOmw+XAY8VB1T06LvNFqiJ7r62QSWU
YdZ4nGI7QogCys+wVC8LMDbimkDJXRgEsUjSVZ/gb6Dnirq+A7cSNLpY/I4DoOm75ui77E6IU2V3
Slr5Y5guada4GVqbmtPJtNAeh1ResuQ1cZWvr2aCSQwZtRNyBlixs+6qgnRN7TQs9JFWUZBTgqVR
wiiJDHygQE/96cLFvyTUCu/AzrxTntdqRuLwA0Rjn3NNK0oQvZBo+Hhtqnbea9oVkJML8Rxo7dVD
wSpYdskO9CoLzlvng5BDfsRH45iPGHF2eNcenCsJkShEPGhrHMqZoGuU7F248avOeVsxbFa3NBHR
EinO+q7qiw8os02jnHVZxrUqT3mbl1OdkLjX4JWwesKa8pnAaS684TnouFCvVocyH4lv53qUN2zq
XzcFv4FVCbtJ4nCJFA0r99eVo4dgh+s7tuEyLVjYWccChyIKYYbDwWs6xaz8VpreSzQeKKvwEUSQ
E7DJFHu5KxOr1S51k2AdAad8+CvCB9qk3kmbcDigCXwl8n+xcTbi5ezeEq6cMX4/xNvYmYxf5M+t
H5pYZ392yy3XlSU0293mOTg/jj6JwTpjSb++xLKE9Dg6uMPvM1OzmjCR3FKEW+bKd031MllEyNA6
E/CwsGjZkozhwpK++RB9AaLnyJBvTbFOmdgWzKmJNeAFJng9AbT7+gLFKmzI2+VPPL6zgLkYAwEL
A8lAwjRIPzxj+SKT19BD+bc4dm2RsZ+/jtW6To47Vs2aCqlOYdzg77eAmiYBOw7ouTTIzn5CIqWE
wVITu96qgb8urSCyPyVqLZfK4yLkZ/FXDQu8Ee6VV0pVu1cwZZ2hEr+ZjrzI5tPcctjxaXr1cD24
gzwRQXV1LdbG/gJmnilgvUS+ajCsLZqH7XL9e3FSvlYRZgm5FdUYOVa4S/S/1UHwhH+FXyPW5BbR
Yqgzp0VGzh2Wnoosy2bH+IwoMmhskLctjarmbs7RvuxNij1GpK9gTAx2/RhaXzcLiOwFUCbiYgo9
YC2UshTfGYZm6YeXYwMzux6H7btOKer0AnbEuRqzqq9veLBa9fQfw3TC6JoRO/FiBLyDGJUEB1cr
FrK6bwZb26H5/WY1khvHB3PiJ07ukw2OrKM0haYAlW1YtTe5j7OsyHDulDc1eIS5fYtlypgnP0Xy
K7EBWLefYEukjCpB08gU5a6MXovELv0hFeghLsWnnHbpkiGe465NsGFYtXGjZLzosjUck4gaPrC9
N1I0hnMQw8rmHFPAJaut1nTbkBsTS3SfUOTG/I03vy2w+LX+CWcbq07GlLgPyfZJi3X7grSdtn14
WtdthKdVKcc4wqU+qn6jdHM4Vq9NXmp5dQThyUyZTyTy/Slhsfq0/XjbTxWQnxgx/VxbbYkWn4Iv
M5iYO1NfmVMkLi2aSsc+f5Km0wywjZg3Sd1oov2FXUXL08dFN6C0yRWpYS5JMgn8IEHg/ghU+TtO
+BoXxAPjtLk5phdIsfH9ROJLeImfb7ZaDb1nHTY2t5eN7c1ByrNpcFouUQuTvLo9qV/n1zZBjZlN
YfaUxuhsT5sbbfdkDNVqtd5v+n9l3T39xveRyQP7/Purwo4CLs09uPmUOL8moR0wgSrWl40IWfiv
0KHnf9zPsp94AxNSUFZfR4gW/jn7IEkk2JTXooj8daaLqzfGoggYmRhOG+bSdistSqnBpxL38QG/
vdkN/guIDkPEgx94NlieGjG+TRlaC8Qo3InnTxjlavEnBdYjd0jG+VKqSSkIJneHshBfwd+1DFXc
GzyxJLAVjqydFp+rYkHRtK448rncgLo1LUWOyHp4aC+RpILN6HSauXR9gGYbpDjEF/cuqDdwnQtZ
ZcZ0hncCrr79Fvgz5fjgkH7Z3rmO+8dZP0yaNLUC2pbyWMHiv/hHvmnDZo3+5w6LfksbQ40eLiTS
Vh2+krddfuzCnt0VSvCUj8nlPE0G6iHopQW+FoCIUV1TjBnxc7HcDKqcpzxScTv+iOx/m0QttW9Q
kJKs/wYK9HpCmXYap9aQTFbX0fVD+rrdF9c8WaRKzNIV6osUekS6E2V2YFIHp5x5th5suMrM6X+0
4DeFFQKtFNSvK5ZQ9RBJXkl6wbCzj/eOm0nKdC6SpTBuoVGrDQAzL1QgG5zxG8zHfQH6HqhtZOcA
uSrdbjPXZm0dZoc1ACT8UqmNCPipbRq4sJ/XXhL/gMKuV9DOZawkQ7OKpnetg088sXqnytyeM75F
eUTWdKsxCXcJfHNtZQP6FyxlJRehJPIwZHi10tP8HYBza0xQ3esX2SoGl2szq7lmBoTvva3Wj7XS
s6j1/6GrMXprZb6/71ENAgL8elS+ECR4WBmMHhLcX3cqPXKf+BiWt+i6NZJ2HwNbwDeeNd5qSvB7
zSWyxEivRWDzHlkN/y97lZNQzRf9vW8qOMk/AOKrAmj2PFqxuvBwIlyPgvo2LtHNgxrRX0RjjpcV
ilxt4eq0mahotaMiD44VkWT18ptReSSfcwdmh00Z8qxNNYWgZxTqVPGiRpn3ts2PzpFTZcFIt8zU
V3uq8gYZwZ7HSB5zjtHIXT8JbJN46zWK5yCwzM0XouxmWVmuuOM5+v+oHybi9Bqwvifrqkg7iEwu
hMAEF4vMTSP0dVSaMDYFulpGInysMfsnDHuLbSnlYz1KhU+uQvXFEWGCfUZP20J+Wup6TLvmO6yp
dVqo5JFRjxN9PuZfl5d15C7vHzRCYLVa4diYAHfWgS+JqaaZmSzZBKzbkRY3E7Me105A+X8qtOjz
0cSv4+lRb6KoDW7uNLWDAOICmNKiD6/ihUWQvr3duAZ0dFBMcOxhEzCDoDhKfEaM4BLOaOFr0ZLq
5aZ94SJYms3OdPcBzNC9wJjxhXd9WsQg9CFlhbvqmed8rgIywBk/4A75vFho/jrnErj3C+2WSFVl
Bdwf/kwA480LTr/RQhzNnk0xwpWElzjxi99PjD6KA6psBrR/ioQ8aJDCa2u4+v+bMJ04F/CPPJ1A
4LhCucIUm+InXGl1sDyzvDkgyyGaOnMBd3OXRPATkSIf5ekPzA3UnLNrcGs3VEBNnYh2GiHf+NFd
JQNr6BD/Gcu46FCTX2JGgyjIAfB/WnSAqFFLRj+NtZKERAUIIMIwPLcaalQ6EdY+XqzSdm5Pd4s0
WikU+Hk4adqjKxRWLDyx+hwDDJchJTfx4wVMVCqUw0AFECXrU9Ctg5s+1Q43x3VX8n4t8+tA1rB6
BmZLLesFX6RCQDEleC2RiX7SSnQ+yulVClcqjZYLd9tiPsu3wrablxQcq9hXAkI69Pp4LJB8GMb9
24jvdsctlClOuFwAMyZXyle+ZvHGK/Ti/JD67r6t8hej/B65SkRfW2mCeCC1AhZJaUUlqoGnW7b7
H9UZ0Mc3d/wothTKnh8stIG+SnOM7MeAe7vCoD49PfBHOZYluDm/4Ct8yey/qWWj2G74LLbnOkT0
C8e562tbRcusqfUYrnuswCLSvKWEQRQEpuawmyguOC1X8YiuajRVOO0F5uFPQ+UnRiDZ/Cz/VRJF
A/khb1DFjzPujEF2Yg4+F5NrkHiIGO/s2mOJSY5MtvDlHGGKfh80jJNK/wdn8fax9pW6LULf0CJl
humotZisAJ6QanoI18Ou9nDGnhe2L9QzAVzip50k5ZJL1PhlcCgpbfMMkT6R6jqLnl+zlcmVPdsj
i4+D7kt4p976ZhbaaMrRtFO19e83VTZ2y424WCaXo58WSxyKncejDxz/jwkTmy7xjSrmuT941+ZH
LLb2SLDDkrhwytpo8A+C+BrR5ax/nIfFaYqRPuYd1rrZIgDwq6oeXsRcxxNVnENTgqA0rqy6dAT0
aEGbJg8jbkjoCg+//T98Ptx4aMSjAgkGBDYmA2S6zg3AmkF8EYrku5MjYNd+/eY8+RmBN5sh9hXo
q6rwA0PyZaY5nfE2SBFGE+dACLB3dkVQu+e3NdAe9Z/F3ohsA8iXmMGn/ZfWYMMAuFgf1vxcn2ea
3ZPQvGgrDyoD81L/c7ZNW59rScruOfPgZ3eOYNXYFDlu9gLRLNDJF4iAumAYECUnneiZgZub/ZVX
UCdieDg8wLqtlA5ZcUObeqb8tD0mKWggYImUXo54Ta31ivyqmAKdKZT5vcnayUcyl+p/KDAdDOlC
P4NJSdvEZXsxHAcbKsHlTCijciN9GtcMyUgTK9xmRuGx97e9KJom165AmxKNMJhJdh1XO14NPjX0
Ic/jlSVg5f1UEWpy4qloPJBHd4hqRSWmnjGPLcinIXCiQ/DeQpZuLnVU7B0Ahzo4ymrQqclaoFIO
uYI91v3GoSsTefrxS1TozA/K028HsuZ8gSljpW9hnQRWDsI9/vTWtmM3dyY+LKjCcVZFSabWXLNs
pm067uN3BtTdnkNFZtQ0s/+oo7Lo6tMcAzjP9QxpEfvEtbkR2Ty2Id+NYScXHq3gVWwSGt4mEmqS
mtw+ro7mjWHmQeQhYo4e1KRuWD1U0H226t/rSSK1F8b8YERJySXcNQsnZbT0FucW/knSCuWHRz5q
Yr2R43qIHsZDLiY+k6yVjoNvgr1YtFzXdGMh75dK+JOvwYlkYjkvaKEIlzvkA3kjGLeLbiIkk6oA
H9gEa1x+F/HDpB+Vh+icDDE15s1adNlQJq4KvZHVEtOauLBPdP+927QV5XO84VEIwvNxLq2bREPN
mJ9tLF/65UwSZrzftZs7RxNX741itcQOFZFrdZa0EmdFVXAoSVgorvaROglbo+Z2wDSENGEZbPNV
rNikKItzWasxGoEZZQwfkHerlBqvfGxidai1u4mvbU2f/O+xRhpyVFSbZU9HcNUF+rMKjpITb8EK
xYCN0SEYahsQ52YLjYjBjwntLwo+QewT8NXOjdMvegFNQ4QuQXiAoqUSWWxNrsUpMnYXYkRt1TYU
rvP5qXVQezsu+JZegsHFgIw0ztgbQFWgo5Zy+rWEQh7LsRz5cDncWHPonokOnWNlt3YMj4pjtfxG
glMaM6hGb6yj2/jHe+Zw7VGTbd2KvnOPFrR+UOIvi0vbKC8dXyQP+r7+03btwVP3FSBMg843WfI9
SnejbmNrbedXkgaPRS7ksweTpykzbZjTj1x5wZglbrJtMfUleZqarUxsfjxYpgeAPRGyjR0Q5yPE
fL7UXywxgF5+SNepcOBhJQPjXjB0hq8lzycUaFprWWt91K7Tha5w8ZXImHn7n61vwm5pxUty9yfi
uon3459PgAjwi2LYTL2BJ5Yvs+yvhcwpdeMDfFtDI9s2QOf7yra+FchxfhfHK+MZLPHVt7x6usNq
GUhlMeV2no11XervCo88R/EAdCFrJDk+bhi60iLjISVfFDgaFb3aOJLkP+HyXu5IkTft8j7eOdZv
6mlcCYu1GOd7DB8oC7yW2pZOJVjt+OrB1/sb8mc0zGXxrnIQC98Y6jfFlMP3e+6sI5aTZAWjViAP
jxjDXCvwFZoSl5e8wWMAVN8KAX8WIWSTaynfJooiYwbQJJWNxlq1o/PVRgU9DZK7hB5hzpX/8SkT
dWUV0BgOKnKAi5UHGBvxtw9WGqW50HCXTvHGlj0zjNbqaUDi7GPhg74tSZ7LBL6itUaLyJ1OUwHx
zFVHJPtzCMpU5SP0iFawFqlkGEazidioIxKah2jCI2illuCxEYdZ8fl7yBAzBn0R53nkhK/nQ1/X
nNb0j2BkZ3uhPt1gCKHUT9+sEbZyYeUSYjF/gMGgt85qOvol12zFCgmnplngaBajTIHlzCgmiseI
dY/fMFwyqbVxDQtcxw9+Y9ZtpYoG4CfDJu/dOfDaztFPBWonSdZ2HqahSdILmuYk52aAZ5SKHu0L
4NkJJ4OzS5jFbmhKIv+MfCyZnaNf4NHtJqSjo+Njpep22vlSwW7Ke2GDeIr0rpptGjg13ERV1CtP
zhx+m8optaYl5GA9UG2W8t0z6nKhrPdMW/u6x9shZF91sHUN4W042a9a7kyPDf8OVavaIf4tZypk
BgTiZ5yBNQpJC52RRZeoNk5jC7UtgiP+SZD2FPmDRo0/24BDpnPm9RXpwdaxOGXqIO3rz8VPULEa
jo/ZnjI/V4m1e/v/jNRRUAO7L8reVPuN8Y7jfdzQXVdqaHwRkSTHXHKSjBTby01t/c3zJkpywKYD
8QAFws+3GKsAipwYa0LfQWcWVXQCI2gAKa1qyq33XqDaItoEwE0XxnKxGbJsgt8BtZlIlI0Jvl60
vzAV8q7Y/a8EJtxjEIzpN+VUKTBy+bpUthW1+j+tU+WSf41Jz6piJT/ZLOI78wxom+DT26EPHp/f
w8NIfM3l83peDYhSo2ojr9cCH9CxbN032RW1Zqhky38tuybsL1pfoGvM5g8V343Zl+S9qG8xSQ7G
AzE1jfdCv9kDV0Qx7Oa/fbR5hdZQZZmBtnQY18auzM9odSKaiDtzGpub8B6IKwhdc1Hgj5EFzyIw
QX5MCibyu5iOWFKzybqMUrPTRI09pnksYiZAbWuf2EK7pnoAwdkEZ/R94V7+Fcb6xu9jPeXlT++J
TpZFX4b6kjpmCcXBAKx0L/hGXpwGcak9rpWhbmoZrjYYiWzlcgqJBqHDeU31zlyMF8FtJkZlxbe7
8Bpy028WlSuwOQDdJRXjk+GPp1bPjGCK/1bLYyHkvAsFazXwQUY5UYpP6CwucUfjEKGxACmKtshA
RfPLZ4iBV0Rvgqc5kNBvep+BgzDSI4uMX3tP8Z1xNPt7NsWQQomRialdkBte2B2xdoiJLxitkcwN
T/OqyVA9NhViVFr+6KX272Yt9keTcf1tl9KBbv8rraCAU8aCCxaHcGEFhoTsnLST70AE4t0qNI8f
VGelzNag/frgBSAvHeL8GkDwm72sPgazEOrYB9YkQWZ7k6mqa/VTQjB1CchJ/ScquOCLDsOB0jWS
aC+AOcTvsw1qr8lZUHSwfrLKBjDXmSjlFbq5lLAjtnaJipeh0WG2uZ11cJJc9I/O5+dmibSQFTOk
DD6SRMYa8K3svjx1OhklrSdx4QO5d+Xw3Yb6GvQrUnMspJZ0PMeay0DV5hIrTKzV5fwiMPGpOHM5
P/eKhL4FTv5lSjXKYsoa3EWKy9Ikk0t3iAJ6RekApXl0UDwcjmZmngLDVz/0NpC+Y0Xx2Ixts9j2
k+Z2Z7cWj9TghyTq51gR4P8bVKgkXMy+GNdNVyyugd78tge9kT3F1oADzgPy91WJkQ/nU7Qxp66C
Gie11D7Idzwb5bvdu7FmIwrtSLheuzw/Bm9DPcCgjDCex0stSU1LewSr1taq9MvolLmqpbu9dcGx
RjyAhTTuTg0boHi5MAiJcFCqYBPd+0cXHrS/ULo5I8fJ6vZ2M915FLURmD+Zx59SSgrAhXj7lsMg
fK+hL7USP4KwQmrDPuXQSGMqE0KCxL05ZZbTorkhHCWcWk9bfcVoisu4e/9a8WZtIlxQRJrRCLHf
A+UmSWe3i0zZiIGUFwIjyFKHaX9aL6BRiYbvlhRdayY0+TAUyQSlXqM697DTSLd1bkuxuV9eyR6L
OIcQ11tH0/ufWzHs90vxjsFV0K+PW6ngS5vSOfMmKkeQTIuIH7aJLlms0YHekpTMI5LYVQ6iFfTb
j1Q3UH4GJJGg+r1uY0+GAM0xMAHa3kvqGQKDNg4qJ0YIwcdYFMdQSvSwBaJaq0VsDQ07vxwZPrJo
VQZbGOn5cQMCTrtnZzyzLHlbH4tQHOrGRmTugID+p0VdeNnUP6MnLRUaRWafQCPtZ7rWZRZDnE8s
953kEB+4I8zE17dRl/S5ETGtr1GxJLuHNqurzI7GWKf2Z/CTA8h74g/otSlcOxfuwpaY66vny4Ty
Bi6hmEOoZH9L3cqUJLNvSjCsxwC8+Hxpg5R068a2aijtbttcBr7wBYmkHocqCNBAl+yyRc8zvbR+
RtL/YHk7XYJdhATlvb248eepwX/12CY68GeTv8TIGY7hlkV6s7YUdadhUzFIYqJF8Nz1V7jlZ1eo
OpJD7VjvHgch/s0gmitPo2kjsi4Jt2JyKjLk7gRk/l+C+kdMY8Bm78Euym8VR7ALppwEzjo692r/
x0K3Hl+SwSYGIQ2vQuu7Nts+hTd749GcuE9soJp4I45TJWmK9v+btGyUW2ImNIP4kzcpwwk/lJgj
bBfdeS8VOaTN6mZm2ZgJ2/nweGdEx54GURFV+Ix3PeWAbixIeFWRD9Xn4jVXICog5WyoFuR+/+9f
pyqiuZnEKsnIlVUixtKEky4sm0BAPU+1jWmjAj+l4JyX9wL6tFB3LdSvkmNEdUmBe9ZWq7sJ8q1Q
1ffxYn0ntMgUFNBUDpIynLBaQfrhCJHHdQHVTwDQqUts0OOSitptInRUCvj1B90QOR96F1Wb9VLq
/+lVztdSB8CK7VJDrIgpApayIN7BK0budqiLwrGWZn1xqleuK6+D3TdT1Q4XWTsRDWu7dqR+lwvZ
CIiELCICCXKBFuN2Csxoa7CJSuTg0Ch25WzTO3FuieTeeWvXujEHrYKohbXzGCzOT+sgi0u163d1
R/lqgp7jzijZ8004GIrdqogF29MakhffSCPGupjkU8t/YguC8sXqNWrm1Dsoud+gV9dWgt82WunW
7jPYYUUFmJOuErVTEijikO2Njpz47XaD3AGtqIV4Qg2lIn5HX/D6uFnALN+Z4+HdGp0I116x58U6
9XOdR+fpURuGFrbk663kc3XKWAPs4u0nA+GBZpzDMi6FHoUjJkjNa+zoaxn6MjfijeO/ORMvuReZ
piHKABuJGUR7r0I1M1Z6hJXpfbyq586XRIQ5kTUTnfSeJy7bjkkSlrf0tsg1OdUwWUfumVEkJMIN
425PO1DhjLichWuxobWnpy/hQ+kVa+fGlIn/iO/ulnizEpKEv9UHY49r3uK7YAZDDpA+KhZ0isGI
bHD/z1JAysrfC61jpRuKrmFFUQldzxEbCh/Hx22kGxudw2avk8aVT32ar/+gtW8puc7wRAZCwSwp
IHfUJwr5V/rQtrKeBTkjvLxqApm98mBOyR5zyoNaOfmlnvY3oOHRIYmBX+LH8CsSOM48Yj5Y4GHU
9DTCD51dsInIr21/TYgadzlZPMZmSHLbynUQiiMmB7jCQa6HjnlNT1opdGfF2tHk9Ax2VZValdf1
4PrM/nOlul097ozGACCZFckjTlX9XMyNHjm7PfxE73gYXoc8AyscNjMl6LPTjt60Zt+ku/b4+I1i
siYJKjWDHBL9dJhRIZkP8vq4oMsQaO4US1UHW1rQwZDW2om1pWtC59w4berNdITMC5IUKaNVG+lp
A3IhQv4xWW+pSo0tjT0dNBrZRmnBCsGBkzjQOsDw9PjEWPYVJsMvvvnBp6B2D6MFZ6xnSnwYnWoN
1tSRdteKccM4E4Z3xgKPvZ02ExHhDcFUeiGFWX30CZB52q6iICOXAORRjeYiiXkEmtN78/Gvsh1y
c1CgCSGUZOayA285ijgpshcis/D6JQj/A7J7z7yl/0/Ak5yivuAiFzNOdnZJzIKBpXF+vkX49sKU
vIq1sCXny3156wIy/83Mfreuo60aQRFlIubjBwI5KC78x2EGpS5A4IQLgR2XSMywgnSbRevJd6X4
RuQrUy8IpI8GkKJmqPxdW0K5TjuGBarBXSmfg5SBQxZhQSADtcx6CaWN2+KW3LaBGyWP1oOrq39V
51Ok85RzwpDaBe21Uhmp/J3gXIycNhVs2ltO8H8GflTqsPV02v1B2R6h7TYGc+yW9pdo301LvXBr
vl2h/B7vMORmmv8rWoE6brz4gF42QsBC64ex0lO1unWOnQWEeA+PeBeABSa9LFiiko+zWXCormp6
FOzSGqiMXCzakVvBDLlAhjYz+ett651keobB7KyWAiiai8qi5wdn1hRwIL+lZy1SGOnXQaQu71Ie
oiXdvUr2xsnGvjWf2EOg8WbjpnH2dUAGDumGr07ar2TjLSua43Fdnv22RJtm9a6LRfPRH1uFv/3C
myt0F7S8N9pStDflhcVW2oFAJLqT6vpiT0nSmNPujsj1sN25lhaDpJfmCfAUqcrqWs1Y3SYf49dD
fp3b/4TdvzqyncmrtOquV0gpWbPKujZUd3DxskSLdPNuw6vigMHytdWAhvl1+gpJ9txrbi6/LlXd
piYdRHDPYHMgH3NK9fZSjL1GJ551pWl9TkfPxmJWbucs9D0xo6H8cRndzwlVorqbDbTACdFkXI08
aypq6p/17l4/tfg7BFjn26UweiHm2Sv5XvS3xCNOOtIITm7l+zKPvSXv6tOYErqQCWf6+MLtHE3F
i6DOKQCnqPLCOpxYfHPe307LCHvMCDQeTq/yLqIRlD+fsH20nIlB+m/bS2EQVigTSNiij0xEQ2BS
M4v7C9QY1/v5HK0qzhJsFn3o+Qz2M+UJr2Of66GUDWjT7cRgEzcBe7eYn94gxAoYM+Ona0jtDEHz
cKh7OrBICFxyNZ7DKWQ/zOD3TRg9rlAN4SAQbL5krSGfeTfijUSVBt+iRSjn+ciVKvhEloKhlFnR
5HDPpUVDX/o7hhKBry5EMyDUi/y6UWADb8b9OA+9f9G01ZXIIHG0ZUYewaDlh264vT5OsKeB1f74
krwvcGf6R5uk47kjUz90aT08AP9cfXw9mgqr0CBX56a5VvS4aJUp2Cgn035sfR+utC2eiQPqWoLx
FyMxHa0PVZjD73kEgY2Svda6uZTWlNZTX2DKVdT69KHW2wJT+B1h8cf/knSfct1v+N1ni7SMtTkB
eufQvUJ4Awzn5GdFW6KZZrHA5SdwGPmaO456/ct3dsoXwIRULOKqQ/EgosuACX1i2rGA4Fik+prw
J63yvRDzuAjB4eJjEwBDyb8AUQUJmxV4AEgjmj+LD8JDYEzkHg1tF5AXM8SQplo3r6vavJJzC1et
V4/3xQdd2oyR+a4O4mIsJ3VC/6v8Jw9fVe/MlmgCi5TjRxtW8XKFzdtNhpOlhgfzAQoCcUv4v46/
OaM55dRBqF1xVzaZR1WMBbQE78t/GXb7RnJjYgwl4x86t/bIDgyDoZDzkEKH0fLtXfaIrv9rIzHQ
hM+V3CepVN48Gb9fQGuVakS6XGxuedzJx/9UNdBIEszP11dSIB6j226ARPl3hTb/l7Y7LI7sZs/a
GMxcdlvyL9FwbuVpfXgl5VzZ5I0WmicQ2qBQPUPH8rwuaqbuUwv0qOAm6YARSPZdlZ1bWh0iBJq6
QtqLwuD+148Nppekqgb1Flrjwqm02rP8wSuMuY+F38sGaQse/x74b1/uZhXQDSRiRzRyDd9hzJoR
pINic7DMRp1COqqqbd5XUjjGRnP6knWPsBwgQNen0HN3fOWF1AMyOIdR4o1eb+xIE7uJlxk2l4TE
O6KNXS91ZjSdoMJj6JO2OC7vHOOTaxfoteR3a0H4GGMyBVrjbuFe63hF+zCN957kmASLUump4J3t
7pWwlpi4IhXlfJH/IbSD/9OdGVIRvPierQ9lHgikbtFIhJbquI1FfJiI76PDuSzVNN0pUy68fF+C
r7YXl7oEhcN+EUdBVVWW9+tzGT3imHiKsXrKO65pk/YRPS7pR5BgYOGTYxqM4fn+T0EmDzU6bIm4
g2t1yPYP3QKspbGd5hm9QrBXoTulVNfZFG/IibPwjNV8SzWtaLRs08EOEVu9FKvU7i1P3jDQqk99
VcES1xZq5EwvsuYber6YzBs6Ll5JVhCszTymE8UPQ8ds4943YgngC7xRVdHlCg01HRUA0kEC/RoB
1pecVR4Cfa+ZV4f4pji7Kq7hMDAQOpkWlcaN4oPhtAMYTpVCGM+OUVfrjNJ1X8JlVOUL/joEgF8z
UWNaaZV+xDe+2tpfVwoGUJuC/NYQGUxT0KkzFlFFOyTjvYlJc7g5tzUUr0l7mS5YuLN7v0GzdY7u
y1JQYh5KoBcMh+4oqQP816Bc2+TWwJQmeVmAU/ngntNHuzzz/k6JdbVTKf5nDGYyDMiynkQrBgOn
Q2UE09ZEGqXyWkIBQJQvPBHewPT8E239PUekGosk3Invl6xveCngGTediE7E2tSPclwjV7j1Lhos
9K4sGYtkzcDh89iz8l06uFH+2LpcOmKlrjX5jZkHbw+gezrhpbn/YAHkPnchoA+qehyW1nSzg9+8
2wdqff9Ip5b1qKkWpDyidiIdIecZbDyeU8f0nJ7/26vKkyv5rQZZUxCqRGipV9TGjtCVq/iI0lcn
O4PTFOHrKfT4cecpD3UOR2TEZILdNoXfKuaNModEQi4q71sBaNgZtSTbrAANj/Xpsrs+cDie7xTP
S1gtpmkAkmcS6XJ1gKlB8835HBkXv8Mvynl+rqkDHcPIa/dcl1HykevT6afFh04ORXeSwYDYpE/H
z78hf3BRQKgcqiWS3M0sUuqtC3B/UUcav7kLCYw3CbE4tZvhAXqnz8My4uzcXsi1UmWf6T9jE6X7
P94/gTD04BEX75NGquPTxX/++akhZjDDImdUxeC1XkCtxBI+euk1XV2r47weXyJTM2u5afMjR0iU
aJWSLd5icmOh+jp7td8l3I1LCPY+MIeawWjcdVi4msrhUiCbebGsH+4LGTpsxGQSDlJoxTq8jr2k
3BLJGPa3dHZN3oBqaHpvdLxPGXlXzz5kx6rnIl3wbsYukeOUEidfdL4FrLf0UGLGL/1or+RPKD0f
y+tTADzt0KCfCIf804toftyRk01xEHnt1GBlUzXQUX4BewCGPpRIz/0lYkOwCdZ+pp7yRcHZMtHt
hTc0y8h1ILo4TwelepOG9z/e2LY7r6hcCrB8gadYDdOyrJdGceaxmQaaVHA/j2fx6JtFtnyEMmZX
ZBiInum3raNTd7VvUPd7yhQ6jbWZL0A0GVaD1F5cLVPzZCv5nWVgR72Mn/iDUeJ0Uq7DELcmBcoC
HPDGOHHw0sCLG2x6W90BIDu04yCNaVS4X0dkAmhhXBr/lCYAu/5wbMrkah7zqOSHv1p5bAolauhd
PIBxlEl1pVTqzjP+m4Bn/qzxSRzXN7X3BsB3GzuCHbDedn9XaVi2m1U9yOuQB/o0wW90ZxssE/bO
lGoBGf0Fv41FOEJmRbL4tExGm6hLPq69heWECMSqQq9bOWQ9kvc9GG3CJTSBcMrsXkzYWhZ554ie
+9q9ffhzm/iO6Z0imGlWdZj/ZOYXAbsD8T55Z0vghSpGgWcy72t9StSGN4+vJcqdRv/gsCLHruVR
jVi5i1JLWPBAlIlTjRfCnJbJ48GbRm5NsTurur/BfLNBrQgw3IXsPHIOP5zAUR+pGkCw42IcvPrX
Nz8OCsqrTVCf8jMc6WL4y0FXVGokDox59xD/dPTGGLfmOCCGNcJlQj9f7to3W8G/C4GttUQFPt/n
MPvk0RCOzLOb8OJlA7S6i0rnNKSXn8sAJx7rZU+fr16FzJ51I32F+sqVskepykwipBXIK3rGe26/
B6mfRcn5pJDzvSM20FbOVhWNXQekegW65rKdQkh3YeidIE7uZ77AbiJT1gxVIGW/iHkzwxnC0hpu
mzCeqRSF2b6x2JUbwqqwJpBSrsQ+jy6TKLnomN1fdlKh/0ItjtCwe10cLH62SHz1tG+diD4rOJKm
yMcEh4VIG2vZG8H1xTGoSP7ukgw93nHDoprmIHUmAtz9oiAxjiCnZK9r50XiLLvZD9NVo+T/JSMP
XMPiuPH+KLn83ebac/gVJgTDYU8Swb7F6s5Hlrs2vzXVZTij8LOiiAgyzEgzT/Lx5aF+XWBFz4Sh
TJ6ZqXxqcDCIahnnE92VAqaPCSA9D3ZWy4Ha0eMEmVSzH/4Co6cpmxjl8LFQ3AwXNRhbxZgJxyNb
VsY5K6y6QTGyzW0iicjL5xrBF8SgN0hdpNlDIvpxMGW8IOxvCexsgsCD6HvnUENR9njdUWTNLJkO
6SlX0ei8nlwgtHv8YfvP96RSoLpTjEvkkW9azb4bq12dIjVeCfP4ThCREN//S3bJka7OtnLL0Gk6
RcK4SPL0g7xEa/VUMBF/WewFmCF37JmiLQanwvTc/9TQxs8w35XZj0sWcdh38zBGtLzlM/g1EkEL
nNiAGbiCnHPf7oGcA2gMLBw9QUcUNdLbbwBY5huirONXhacSqoxRLr2xu6uPIPaH9CVXCRw1YVjK
VyWIRQsmg02pPqY+MHO+1kuBFdwQyfwaL/oEHTcK38HqIKJXiVxRU/9K/GJ7bPVEKSvCfw1G5QoY
tCtXxGnaIxJqDJMQA39XjaViY3h62TRXv8/nyFys2G+28KqbXNh8hJaEimer07Iy9s4DgyrM/hzT
UW9M6foGtdOnaIsCLALcbgQXEz36OBQh7Pp8/dPB0MEzV/9ar3YzlQBTfh+D4ZXydZPIWiKtcprK
6pyaTmF4G9gzsp4qGWuBTmg73Zt+ZrIjEKGi81gIatLlzFOdeEhS4Oi8Pw5SeoZ8zr7ULO8ZDfqa
fBc1/zXsF1X3haLXHmaG2CMQabZ7r2y1Aku8VxidHtxgXpongpbFczvxFWadkZMit1smVAmBZWSA
UKvAAOb6C/DPPUMBnySIqM3TeioTBfWR6mGO9qN7Ktu9jgM9N0oAJmHytfd8qgc73J4LZTKKrAw1
Q5HsopAWmfmjxrCLa/V/jrQRX2XfxpLqjOyzyWHRRxNzvsG/u8b5TkTkgVUBpw0G/4hxscokcAr/
pqAd5JjcY8QxinOQ74UajZKh1Y8lum7j0v2gcGr+c7Yo8UjYITruftDoqy9DhVq4BmEz1Ne8yFDi
VvoQOcb5JYbfLoWboBeH8Onw/mP0YFhJfYopK1TV5a+xiuRp/Plt/HJeXs0i6U1DV6+oWThqrVjl
TUU7OdvgizSfz5QYLYlXrJcwFWWxGoQ7JMbEhPg973jU+mcguhcGpFTohYTFBUyjarZiFIEI6SNB
+0DDmybjX/9OC2kbF7zH+l+OktBSAH8tK3SD/HGJTQnq1KcNb6cLjtClC46f7Munnn/hmN1mQ6wn
R3/5P3Paqj/b8X3a3pC298+5UPqFiv4NbvOTCMvlOW3VnfebbjsmpWVejNMvazNudnxhql8dXYDz
QvAy1MqA1ClMF3jFr6/4lglZ7RmMqJyEJbPlLQivzyBO9sdDhWbTaL3Kz2LSjtbpA8cKg7GbOBM/
OXXLgFfRzg9H+PRrA0SX67OpA3Ej1bNUE5VsfaitvmzfZgb9YXNdqZdPYzZaggWPmWoZmuQzVD8h
snQC2QupBMD6gwzT1LnM9tq/Bm8a/LhRo/PVdeaiTGYeZzNQ2MDZm2bParz3CZ7hBopwz9I5Gu6a
gcEDb/7w04WEB1bmhQRx6GgE/RF4u1qgymLflx391gWZ7jy2p+QSspki5lUKH3vVV0g6eF4el+If
zs3v/EcQVS6jXzGn5Kpwp+ua5j9ALX2gIRA3RuwME+bIBhlvjRfADPcGTbcRyydYBrGbXQ055QdP
rJuQdVQvUUcWMOyqWVYjn0RAZqHXN2YdkMPJrZASOzOk3jPVSBxlXa065Ml3xIcTzzAZX9elaGVE
1lKAt53xruIceiIqrdxgW6nb+KI+2Z1Hg92felcr1bAssrWeKGhsiMa7jyxTjjf4soocsms172hf
49zr1jZU6IptDCQFcJPFD5y1FMHWAf//q+6msqo6rgG9BJsGWy4BiwBik0tqv42MCgGnDen5u5Q0
D64FVYW8+jNsKlIwPwKA1veiyl69GAPacKQFP8g4yukbocmg0Zf+01qdWet644Ja6eUpDdOnzquX
Ix7H+u+jKObqeurollst/fa8mTfwpw0jy8NIQpinZsFcfbwnywKWJ6Mqox39T++dhXoMCN+CFd9R
DEwHcD2rowvVaND5b7O6kI1E1w5SefLoLRr4FMxvZ25X8PsHQ+fACb/nQVBUY9SN+yfRt3dmgG0D
7C0IgIchPWAeRvvjlBtibmBYXWR7nXT1/FKt1pXfwlgC7zTEHe6SDqW0pMRK/Cx2sJijW46wkDYA
ygzdc8C46fx0PJedy92HjJVJpx75rGjrNtmhbNd3N0tv4oaz0+PM6Z6Dc44ZHIisfkgCqW0MaWgz
HLFgtugE8SiAJb8mRXGv8rUMXaRTzzjpLcChJ8CMXpahav8ZObTnlqTw4mLWIyFYOYmwhhSLpL5e
oXUE+RitmaeptW2aIKnX/4alk4XmozFr7k2da7Fxtyy/HMvCF34i9t/omwMKiBhBMSJtKEz9Bm4D
bEhSfxyGxQJCWjPpnE7nVA2uzyXHDvV2RXmbrbCSuEPBYvGjwOhkJ/md+iBMnJm18NwRbZSuyPgu
5oNtUN2rGqCrjrilWtB54i2nm2TDVAeA5qyGioU7dCrkDTOKwEt6eK2iVn/eZJyMfpXc7Nw4IEi3
mc+IXn2GQwNd2uYc5Q49hlE5fJjZ6mA7dZ2ZsfDM1JimP8kY1YSgWttSIWZ97FF8u1zxIryxTyWj
Wt11zNPKgGjPB9VxHB3oGoJxZl2RARmePWaD7Xmipw4325oqKTX7w5e+nrasJ4aswpGXDqaDL1ih
QdGpIgXUqwPaW4+symAylax34dECwAlnibsxTEA3GDRLGAQ1FFAakwalsfBEoiKEoaEFnYN32VGM
mTAU17pBNdSeKjf0XB/feXiQUsE51X7HGRQ6Uv8VoOr68TkLMArzr8A5K3migDeimqJOEKBMNKZ6
ss/KbD0qBiWXhS/V6lxNgXDQKKnbIIAtRQa8MljIoGAbeIAB2FcIi4Wozgbu1eKSWwc1Yqm0mqbw
ARHLyQwS6EfipImtnQIdJxGYjIxflBD38gwLO9lR3N/VlrZwai9F0mMYFr1PGgZYcRwuczMd/kFs
4mC93zmaBApAjQbBMMBY8ZvfFxPClwF6+E4VlR4mmGobCaqjlt38U7ZhqrxPNvr0EJGNZp1LFYMi
htTyRtBwtaeTSXb3i2aQ0DKmDH+WDFTS9hUzl5RXgIAMmaA/wGvaEakBsMpieyEZ2N8SKup92IJl
RQvyRruh54Ulo3E0YI5aglCESLlPTb0zSokgcOEIWu2nZhtc4ZB3ZwV5EH3iyin6tkNVVdM9i+HF
Zuyt2c+ZPHEkQ5RFAzjttwk5d2YOTr+CmO3j5yGsdBqv74CkdVwT0uYSNVUaOGNOD7I2/0pWBZEo
/nnYp9HXriLQHK0VlNVzQEC+aZBn2a378mK75tMdFoBejm6aI6ZgC0lLM71z9wIz924BtxswBdLa
xZuBnJSy9meW4Gy+TxDlZRW5jOHK4XAu5cMQZMkXpBYKCjXedTDj88QkYMzKugYz5xldvVm1IOD+
xu1HFvwMFNT/EMgHr4Z0a85hMkczh+yafUuJeTV0mLFTpVnO6T64hBF7vutctVGyU3GnBR+dldtX
FB82pseJSwGStsqzROIy8ao6BRxIXNtWKXlPa5VDgOl+8A9c8eXqccS08HrJ7P1wlgHnDlc7WI7N
7BOJUXgX4oF7vHcTWKlUnWVYWRF83D2YkFjS1970KhuHweMSUDma+dtVY1dRTjgvn5ExFYwwwVHd
YBJAUgfZPblNP1Gur4zrROf9uy2CZHss5syF5VYPqhNeC8NmDYozH8Zvx5INvSGkTSp8LeowDzKX
Tl0LQX1iEzsqQYRhsxg2uClhTHj6bKbdF/ji1SiXlWLxHW63iMRMMIQf9Lo2nkd8OFFqi+Xl1LmN
cCkUq1jqpOfTXZOI3wLbqk20JgiFTrr0vSQ8BG7H0SbDHV0o/kZ6z6sq05+nLs7E1hb3ZQBwdFWY
P8Ek+mrYqireRRaTw/f8DuRS4v+mO43fXEErjCZ+ap0XGJG2fYRn3OlJUcNnCDIPq5SpAcitf7mD
esrM++aHbmKXA0AaQdD1MpEN1SEqotw5eHWwmwU6vm0uTaZ5COy/9Y/hhqJF/AqKflqg7IkVNGkO
z+fR6sxjoWWgxvAdXu26X7IEkq8R5ZauGw3+pS8KTqjePJNeENCIVKpwuJSRkF36Z/dBA7PCwAZ2
5OfeYL8cartIYS/Ny69jfm09JaVz5VA0Rt7VznmJNFm2xb+fuv5vy4XlGs/YEoMnAZkFxnyWZwwX
jqe7IYJe1ar9XTDIGhLB0sNu0ozCswhNDafY1TV0TWbuTqJJcMOZ81qumV26uuBV2bUEmA8YL5wg
W7Zth8LFdQuyfaFNo53VkYEY6NNPecfjg/yh8MemXHMu0wR5ztVS0c/pAYvH56fldZvBHQxTgXq0
doecs+Yyj1PI5YG1a0T54tjVmDVAmvvF4CYMZnAnq95NAXKZB/PZwSysIBZcFFx805uNYPZfJi+3
73ceVLOBT3I6/d16NhQWH0+zf5jgS479yLg8OdyDy1/dDGKLL5tNnuEMtTnWK+pJn+nmP9jXu6fQ
SuxR6T97aUAMHhNiQfFng8SexASrCsV7/iqh/w1HxTaL6UVWjf8Te/QH9eXi1H2/OhcVmbrVzlu3
2QEr6HHN5HJnZQ2iVDVebssKrrh6ugivQniexQz6XQAMGvAbQnH6xkvrsTFcUureHtA/DsLdys+e
Gqs0xwF399PetSU8RAnRz75lcrT/sy3fQPUh9jqI/PyJEXXprxeaQnRQw96XplnZWYR3usQvj+Ft
EIlFKVQRQzKZH8JH6EYMf2WQbcGvqAXfq3A/iyNehTMYKnlUfEvPol1RKv55jZpsHfkuB09u5i+0
7B/PGGCt8WcKUb9uuZ48ip1kRjqVzueesApr2j+OrBSehzP6doo8e2YMG9T3tldvYKQ4Besh5uIb
6TSLZae47QoWEENOG8SHshccxq/yXuRIqhc8TH5iIwWIQje1DjTKY938iPa7oKFjTdFy0P1H+gZZ
CoxnRWsf2t2ZbUZiwt9rmr/e8KLs9VuGdsMMXdSZLUe+i+kfB5e+GmfhKiu/wWsqVjWqYfAGPfOj
LIUZFoV5RbHQrXb4mtihQFDkitfPyxF6lUDpQ6gdEwfm5CPPX/4ixO7Fjx3Xio1lZnEnLDjN/Yqg
cZjeMqedY/vLBukWTEAZLPBdlzl6j8YESTDBFOul+C4ff2qHhxVyAUuuAr+shsEE7oNeXVXtg2Po
JrvK7qt7qhm3YeJqrDqM8UQ/dCZrPMJnzcm8hzRwIStH3LLyuEOJfvQ7lne6DiB0EI6hR4MJ1lDd
jHQa+7eJryz8ukErRJ3uJ/HzKn+MT2P81oBdqEU/ft3/X8kD304rDemzCFenHGEGnVZchBgQ7g9P
bo5Q3INngYc8+HHYuM+v97hOXpQP1W4ghvvzWukz9on3+e/1zOWnZHjbPRdp37Orshc43FUhN66/
gTkZKZjKalZKEOzhhwq0qpbqmTU/i5hV5/Mmx63SqYk6xgZq3zEXxb33OF062zS9mkA9rvDWyKA1
NT+vsv9fmuVVdg9ivYDRcv7ozx8bsonBd7+a39/ekYht23YIwL+bPIkgNfecIHZrUsl0L3vQRBS6
LQKxplJ3GVU0ysNOz/AJzdzgBoLvPqUjAKw8hxnlJTgT9Z7KL0yTY7I11GDRLONQxKq5rGb7k+YX
WCLsD/y0zRaIxXbjSETo7P0sXAPBbyoMKYAqqd6l8kpXeu3T3Md97hKb0SeB5VkyYytvES0TZA2r
u8VhQ8ylZKTKMY6UPn9stLeHoY+h1ugckDg+2qjIlqITzyJqhofNKO/hIeRf2gh+YQjdZzTFSv/F
CLewmBzXr8TlIJkhX1bKfLVwqtMltbPeYh0k8aCea+RhaWNN8+8w0S322WCh3rsC9XlQKSYqw/Fz
vKRjIvnDxysL1P68UsnXRJJhuxV4LzFHZEnMvUebZzWBjfbkggKe8kRa4XN/X9w2W69yh68Z97q6
fa4ScZdzArh0J1BA3sbk8HWUvcNGC84Uv5x5OU/E/jsq673pYDwEeqpuHyCf1qtqYQkq0/2lPq/q
zosKstZPSgLjY58xsIzedKGRS08+1rWWe3p9lAVtNto7L9O0j06s1ZzJB6QDICgopsBr71tITl6m
ccVuGINk0V5qHjbe5Q15uiBHK5/Nt7TNks9jhZx/ixjjTmfckW7XVtAg/LGBvcRrX9Q7bCNSfe6W
azNwrTkw/EWUUO0Pj1/nPU/QJiNd8od+TbT8Q1ScdnCelLX2IPD95Dw0TWeiC+n2hTjICiigTZgq
EAQWoD976FXNbV2OOCeiGiki86KAyTMIrjna9nHyNx/0Q03UtaCKRQZEvPLT5gunj6bMSvB351Ky
7d/6QSaAkuP6onLcXtEIX9vZmgW7HRpmZMdo6/8eP43TTtzNBIGbOnLIg3w1/NBvy3jQj1dQ0of6
36enJTrq/QBT/K0qBwVY5agRzjIP7Hd8d9c8+sIBEoneLJzFYIA3oTp3/Ozm389JNf1ugRgpp6Fi
6b13QIx/vKcGFtpjjfI9iNrux5cw2N6NkakMvx05Gvt9Ps+ZbJYPWNxRk3mevcxr77d0/5BheO56
H/oerYFg0+XxkT1CcKZW685ciBU2QRLUGSrtTlF8qrddAqOyVGvNRKTxRdN2g5MYax4+lM6I27TI
CkuIVn8iT+l7uVyIwE79UqAuuVYxy6mIaDzdTDiky79BzDNwnwJTAi5IFgzmxwV/BSwXj05oEjBg
LzEOjjIgbfAyTv6DTNPuSzBdx+mLZd9cpxiOEZ5FfAFWswSo1elYrwHgXaaLED12GMxR6yLBk46u
odUuWeFjpSK0oHqj4cDJfAs3kiaeIUPCuEus1ZOhOP7GUtOlgZpf4MLY0F3NMTymvGObci6V47VP
w6uauOjs3fBqgA3JVZiTFCHrilBjjmqsQpsZxHNpB5u96XTeq06a8/2d6fzx04Y86MDezUTA+JDR
ef2MKz3D0StTM0oJoLogNdCzfZV+qQChrMiMrFunTB3lgNEKDBLcTgd4v8dUdXTjj6Cx02lL7qvR
15X4wL0kkntZWRXoHH4CEbYvBoXzG++qgU55QbGgHPaZYvvV6T+IYWXYLmiHtr952E8j/L3aRg1W
Dh9nBADE99xQ/YvTXM+IzzRwgOt72B5cMPBJd/n19OUZSyTAewSgrwuw3u/IbKvwupUgAABEO8TZ
0eogr4Bm9xFhPbpuB0Skq0udbzB6gfI7Z055IiKbw43ow7wBGytjXsu5l6IabMHGUXOt90aDtWH9
VK7K2xSmOwhVObJpaiMqUpBZwf0deDfixZzNPUE6w1Jq1YrpCIZ3/L5VweI1EYtbN+Kofo/ERrI9
2Gk6tkrvwnZ6IMPE2+NDekS07Fn98mRIWuIbQuNgvWYTDHtSXW0MOub17kEv8g8zUmBOhSad7kCA
5sQeDFOpL8m8PKBM2u9ZsFhg+drC90BH7IpJ4pQ+lF9LU1p/sRmYRfRj5k1+uPTcoNm4VzknM+n4
cmXteD09KXRsMvUNPFnxIWGkPEe5PERDqQZE9GjHc62XBqTs++aoWvA9otniQmfheB8jjUPmCA+C
5EmK/QsI3Sbhs4zgzY1DQ5WIr5V8k0Z3Bbe22u5i91vdKaL4kpjtfZSCpT7GrxoBAedrUwEfgxU2
LwE0WngrFMqBQv1+Zbx0tl5JnYQjURWVxlbEN6k+LJ1iDHY8kBKq2syfTfORv9nwcRQOCpEFSsq9
vHLkUN2sJml8zcomZbZhP2fdjgJVTG8kKoRg1otOf/K7cEQLSZZhhjGX3uyl33C8rI8rIBWi+7yx
jQb3C2DnHhvcq/gUtrDtHPDtKHrcRyLmlApMYaPFz5+cS6DlcMnHjafEHi0e+SwRQzCVvslXmDcr
p9QQpQACOjODa5eE7/wxN02J0lnHVqIFUHnUSA45v62ANp0Mz3V+jqAmKTeQKLIuCpviUc5RP4lv
IdT5UTOQrxpL/mcD9NlAWd/1RLVYtTc3bL9N64UKciS1dplzfu+4HIClmkm0jgLo4Zrw+DCy9e8Z
lNbHWrWcYE/BzsKjWg+DGQdfGW+cKJPE+33/V8DNOVFPIAUCX0hP2+0NWePxM0XYSHNqQLeJmvTd
pv7IifsmQ0eYt9SZYYMF83P0TrIXcSpqBd5LMNF9YCHfaJOTOFAMxcooaQovnr77zvXbTaMYYCvw
KTakghuuvBQQYkFIwrbgiEHW5jI5Y7UXC4rxS82LNOkB677mWWu43AFLxDJfXTPd3fh12RwVH6Yp
ORKQ0OZnsjiiUh325+eynSEMVv9RGjHZzBst6Dtcla37CizTyaP7iXL4/gDNPVEJRBJ5jXzMVK4g
5BYeOCimZgBzFGo2eg9N6Mxya/BISdeDeSVxLcd8vbdzCYyk3soF6OIovLVh9Lme3NKrWt/srJ2c
DKcThruNcZRiu6eWrIjYNv2nTyv7+3JIwV65sxseosCfcwF48XE6MY0wLkhM5mN/qftoEYQShaUi
+nvIkOEZ4jmKlCvkE94NEYfidJZiRTHJ1UY2Hoz4SrzhXg/Z6mZwMK+fzI6MSSIjtIcDnD0Utbfp
iipCzFXDcPYnTXnhL/nplRCCEXAkuW0YXRPTCIdIv60koRBMdWyyF6Rs4BqiUT0YCa+e0dLxVQhk
GzEg5aw40mMZOKUeiUsk/V5RRkFYnV4PXd3DV1jY0GKczNCg5hiT+5qfOJ5OapAnqivlhyEWWy9k
86x728eL5W/X8njouxikjHr0+X65TBpE25w5CH/t/a7jMMfrbHcv2ng1Lp1YzzYE3QPyIM/HVPMu
A4DZMrINAETAR7tmz0HODDL0peHeoUvAX3WVT7X2ePnRQkMWamdCVB9aNgBZUrzxjdqHUYrwpbtG
bLXix2JFom3Ia8Oag3anSTcsmSTfL3nHkWEH1CzhEZ5I2Ytb/cTIlK3TrbXvH2yR5XFxtG/NNPOW
XJueXP4PaMYolk29Gz6LUhOEHyslCG7gZnYxJJAbaWgZnymLI+TkKwWF4qm0jPRVJdE3h+v97bBK
gflwg7egLaT+DYwKPuZv3bCGEDOKI7P/nopQMf/QUo511zf6n9dXudH8xxkAkqIDUY+7qFSWES+r
Tulm2r1sB74VmfADeUDsb1+gc0bEb6Hz7dlZVspTgcgr0EkCvuTSmWN1IDx1HlyzZqd14ypg392Z
Z2TB+0KnoDqk3OOkg8tTc4Vb3ABS90/6L9yy1zMatB0naaGHGHZTf50S8JxpgwL7uiAyvtZzT0xy
gRnqCM418AHIBL0oDv2bglbHeFcvWifY5sc5opoSPOMTK11ClVE3MECnSTAYgIypBLg/I17J2raf
sd86Xon3JIs5V8XxOiu0vWNBui4elhFnlQFNIH8VSz1vFPBt5r9M9fBx+kCvUfdPVF6k+ik9G7fl
iGWqXi79Vdzavgvs+Zt4qPbToeSLbSfyk2aZmo8WhWAjYzl2APsDvpk8Ur23xIDm3FgLvtn5KTLk
UUwIKxaDAxlm5HxOaXVGKJ03RKwoQhzZIT1oKk6B+DOO4sBsgfW+IQA7/nq6W+xL28uIp6UQGqfu
ndbXg8ZeoLHMcGe6TB16ZZtvETgnqO+Ij69FzXHyDsRq5lKitRk28ylV8e53XbmHBYIi3VI0W2Av
mDc/f0CiZeq2WnNYCQvyZig6iZKo7Vb3kEpr5bVz/vzL74uRmHiZnMxI1+mF8LMHad3WB7YC/RYv
UjJxYoZXtGEizv7ZUGyd2M/InAsRwmr296DYN2NN/PxL5mKNf6UibLWTtfNq09B6LX6coQS6yIvx
XM6u0AyaWbqmjnZo4XAfXVg2lVS9nVVTwO/g20wOJSN65+DygVaGl9HZkVNFs4Kkk/MD+LQ/2flG
1XSKi5J/1uBEyL7B3bCD59zVKBSxVo6pG4O/FBTLr5EjrC/JA8oOm7RRQIL/4L7v7iI62xgqVIzF
WNLTywztEZZzrJl86gteGljsuUhLKnGTBPQvmo7ZyfU5KA80igESTc6tgTOwV/+Pu9Dl2v+7Gcjz
avpXAwE1/rM8q+D8mMu8DoisOPz6woiRlIpizZQOuvr/TVq+KlTxKpJLtHmJHQ3hkUF7XzhrMucf
q1p4xwEj7FxLjd3BHrAhjdu9HO1przW25vQI/H66tcCS7Jw2KNjQ/SgbTlrVijY59tVf503jVoNg
QGmoj+ZbICXnFmgm9ArtQq+5egxkRIwODJZC9JqXDhK2WMd4Ts+3K9miXmjZE2pNO3D8W/Ay1eaX
YjPOEGr+Mzz3Tym94X8VuX1yZrgYi31nYfJ2Xi8MyLNos5MX7IQm7jzAOKIVKVoy8SRbRDSVFTTe
tEwoIHGOkmzHv3srSyhi1Y9sUSgq+1HQkiTSC4H3DTCgktjuUxEObMQe5HDQJFePNVtEcubmwdw9
097fzvx1AdwFoRJjpmS0Eo+5qh12hpF4ozGlCXf/nI0yvxzX9QXqPXVP6eDOXxJZXEGm6uaS2oGf
ce3e9iCRcJwlldQj2DacWBfGpaaPLXax8bY8LozLqesIjSgQ5VhbmB37NKSp+jdQ6Hg918pCgd55
kjrz7nfRvBnm7dCWp7UbWhR2YOoi74Sn1yLSQL6gaCHRNwmAejHvxerrkmqE2OjfGsHHKB7mDUWb
McE4QDmZI50LXGt1ZsAl5KfyiJD/31IZade6vYMET8pJYNR6nLDHULg8rw7JvF0odDkr5XJ2LcOw
+jGKR3kn248aDRq68G/b2KGitHkqY2chq1pqWeIaCCLAfTWF5W1JYcvSAkmLPdpBEI+JicrR8ZUj
OF09LRk2OZ5h3iChSeRHBp0MId66Zy6/pe4HpGGKr1Ms/xoDjVqy6RRcCC85yOs1ZvnOgXkuu6TE
Gfu881+rHLRGyBQ8ztasqXTzY54XMjQ92VbKFGoxypM+nF0v4IpYe6IqcH+/1I1ju1sRvk6MmA+z
PuJFAf/nBOF1bs2/GvC9xv/XsaFySUsD4O1ekF6jM3fum23HwSJpteOISSQn8Qm/wvS8OXndvKrG
FIbraWAKN3exDrTaK/KQEKQotg0FerwICQNuVJP3VZVvXW7rHb1XQkNddd8ivZyPlXuwV0laDZj4
nExNmocOAP7vfTjU6eNYjSVj7r7Yby3XLFHBsqxApyO/ca5T5SEa5CDigQIZzZJO8m/SgeRXHrqL
P8deUMnUj0lYuSVj+/wUiwsuqSY4Ex1g95XIA7+DKoGr82gmUREee7cCLR0KSriymP3WWLEyQ98Y
sFHpsnwmGDSzeTNHDaAwkNtMoclWzysSo3rrGGnbh8bHHrvfKF2U2pADtmlBSpYinWww+M9kANrd
9KTfZHtJ01iiKaV6j2Jm1DliWDOA8fMmPWEvCQh06hIM6otJd3yBhykqPTGdA57slEYL6dLd9yD4
HMB5ozCLBSYWlnvfCbhiHFmDofeDppycTD4yFZsDx4rdBpZL5gaJaUAyT0FfMXbPc6NAL8Gd/Yf6
Ssb9QFcsqe04kAqBUaQS6X25kepLhTKimEI6E/yMpi9vPQMC3wgwhX4t5fzEOuZuIc1kji/oM3Tk
/uL8OUL0DI8aOnmk+AkAmv41vIbAFdEvvlLaq6VQv3vAXCWnJhAsUmS+ehM/Ni9p23BTuAUVt52Z
xyZl/i/PJOpUv30g0pHuHqZxjHk6HWLry79RbI6IcDpAlDKLJhtqJRIhXFqBrL+GBV0RgcEEN3F3
VgHF6W+agks0I1POUA+6aaF5fsrXQsvsopHFcIgjaMQUQVJnF+lxRORyIbGb6iAYX60CkLg/VrR/
fpavB3xD4ClmQBGMT9yHMVWAMfBczafBWY7ogERHLzxQWeto0UGJ4ZnfRmc9TfyrSd3x2PHvqgbg
JGrpD0pgIDcs6P6R7/+GVfhQCKvxOWIVb/SmZMxgRgR4uNpkrYOfeDXriOsK0egG76vKmKGV6jZT
F3lApuhzAs5bbRj53r3g0/wQ7e1yiNeAFdJ/KXZhukYGWnfYJbl3TSxH2ZJ64JhqZ2U0anN+ojBk
faEg3EnLAfYaVLAovyd4J9rIG3apEbPRBXwsKRunn0ef6HctUp/TlJDvh8HkF9MMOHfXurQz8utk
cpnxFUuCI8k154QuqKh7c4OkpvK606aE67udAa6WSXvOyhvOaytSyesDqbispUvsH4T3QTQX7Vv8
+tU1D9nlNmF87+OBH/Y6wYaJdHp6cSFv8uo3n0VTTaVWVaOcDq8jyZhuFcBNGpXE8q8SqabFxpMX
XhAngQ2wrf9h+BumC9PG7kU52JkjOGvsnUgWHF0ixiyD5aOZz7NXQ+RAxlGAN56vulLcu1X3v50j
tdgMXimx4XbQc+PwD2OHwUvsV+IihQTzYRmMwO5OGd//adRvs3q9sDSr9UNfum9aPXzJh70iZ+0K
tiqW303DgkdcvZLgNPaRKnYKp/F8AgvunY8tCyIgVeS9FHNpSlHp5D+gaPfjgXPi6m7wE93aG1cy
/pNs+M3N+R1+/ajaBH6JCl2z1ymD21LnkxmlHSmXTTnkAJMbsxfbA1RHlLU2XezTBniP0LlikseD
c0dTVbzv1myKKvc4zaRIHHLLonb2l28XPa/9j2dT8RWSvwvFEdvRLuqg3fnqJgK9wlhPPK8sjIk0
xD+tbmGFczLnx+ugqijdjbDqqtYFWOMWHDVnOHkO2Ae6KGRbJETrc3f+aagEyVF9gQXmSJKBvmZP
tdFM975meC1eIih6MeLdVDzAxeGRtqs7VlpL1IYAXGxDiF2KufP2uXtVzZ4l0iPXbaVoheZrjeT5
JzDHEcGKxr6z+0LFDiFdctBacLPl4SSOAS5pG04lCsTiZswynKrQUNVSK3Q4R4VmCkJzU1qPHjEV
ps/Y6ukdEL7bbe/NUCwoeHcJk52QCgo7eGI4vMuMI6XyDgr3MTmb1larp+GePHo/3E87SxxzaMtO
0MO4uuaedzrqx6vaSnTRBd/RBYQPoY8skuWwM06gYhUQ0YYvDeZpso7+4ItfvnmppDwueD1FvE8h
CVsTZi/QAS/kbZeK74XCFa4SgU+xTE/IYEd2SaWhNX6b6MAWFLg/t0Sd7u0PEoip5t9hYHo3tqnq
+7oIBCCGlDBbrpfOOUNKypurca0YzXYBLdGA6kfDgUPQ2S+JkyEsCZYhPru+lAtVB/QEbDFQj4UL
xCX4yAKad3b/iFLOUzv5+C9lXt6ysmZgHCopddsRbF3ItZ+y+24gGSFMOaGjgH5mY4MmMVaC0mBp
6MgDKSKqo4z1gY+7NqwTBLykVCXiu9XRHgFbPnzg/IysARgl8VEFmSC0SnWiSHuB5Il5v2EPyKLv
o1vlVM1FUuML0HCJMNmXfQY7/sfs55YO4afdGuK9OzDohd+HjkKgeiJ5a7nVNcoxKsJFELR9aBhs
WSyBCOO7pDiWCMLzlBrbGJpr4x1UV7DKGCfZzpbDtjPZsSpNF+1Q7B56oV2Bo7ov+NBVZCfZLZpz
2fC9xBmePpWd9pA0ivGhl0EE2e6F7cjVvtcdxMIFItlVIjP2U3Lh6tLlH4twhdI6E+4g3frdy6rV
kZNVbZs/YJXh2EvQM2M26EIwFnX4dRtFUrYLAs+DcqU7QO/YD4SXOpCGAYjUTvt9mGbjCRWYcwEP
mHDhnDEHAs/iTADQ4nhB2Wuhb8MW8IHDawtxk3HKnMH+aSOkQHOS0KICLtVP7tCSUB3aCrObramZ
/1LgbNvaBjlJChwP8igFROS2UGYgQt6soIfvuGlUbo0GbLL5scWWTA2Du6K8hfoeUqEmoR7xFIj/
/5lW6L2nD6/D+5zqBJzJRG6SCYg7tGWHbAv1OyZUtvjM/7taCsRtcTDsi4xVaOrOX7nbizmpCWwL
cjBfSE+jFVItcPmfsN3O9pll4ORr+pZcgdJX07I9QVt+1zLhr6UpV3Iga3UOAgA8ItG/D5aL4nLK
Ki3Em6E3Frt3ai5fB4HH0deaUnb1VnwaSIPnQ6Op/q4RtY5mOJXJJBaUXHkNTbaGRVmUEqFJ2Ild
Hj73aEx8yxTO9fkBoETIQZtSuHS0jRIIEhpovXq4CbA9qpKiq8lRr4hyh82qpik7WAdVZyD30HFu
WgUoKI9bCbFwijyj1cy8065/OkIKpcU/P2t4lLZc5Ps89dcvnbp32Il65dqVUL0Vc276YZ9mB7C0
7qzTdg4HB1IuBiczm7VG3FizY6/XyQ9ZLIdbtEVMo2rYGsKnn9LMl5eLTxcXMa2iU5u2M5JTxA5r
1WnoGCF7MsikAn49w6ckbYF7v2a8VOE0vqh6wOFX/fzcQkh/20ZRky9loN7UWXNxEh4aYB8gIFr1
PFOZXAyopXJI8GwgaUkIXXEG/19OlD2/ZVeHSqB/osGrvigD7O5YeUH4sqoQBmj+Oj9uYVWp0SjM
dZfymOgquvsvDOlfHwZkDd1o6YQluqaXYzcm6CNfdFPLJpYPcV+M6yn2sepW/76FkXJhbPNvoCDK
luYss87wc4Hdhr/tr8ecc48g8OiOFffS8IJptRAzu0NQHQA3yzoAQ4IXj6qfV5pMqnHy52jnLdHc
90085So/48U+v/NM5gdiewpXP/XAzm6ZFnIC1tIWw8GeZrexIXyDvqaxNddoKliikOkfQMoC1Um0
Xqb2lUDY0MDxDrBYpCU8Bx7/fE1Lb9Zg6shXi6SF+I6Znv5TVBTBzP7ycFtDb8C9BCiRMk6gxZH/
PKck0xjtfS/sckQJrGc6tMcTDMV9PJd2ftxiN3EfasQAOvpDGeD+ctbbhhWqkE9J1U4BHuLyf1LK
JUXBXuSlfWFMdWfDD5r13w6SPsRcTMTiqfRkgdNNFV4RW4a20oz69R+28H24jWBfjNyZbI7Ow9PH
iUuXe87NlDo4d6/xc0Z+wIG8oAj52zfKV24Q5tKf3WlC7+ZVYh2itwyviSo1VFnLh6vkfBt9aRIx
Xoj2tgMu7cZxkXC9vIsw2BYvJ2R7cyW4gDP0sw9V5PTA6U6No9/6s0bb0dAn9pmbUeFEvZWmouuF
7lsyy/hs0dzcPPEQzbNQplHXIpIT30gKo2uY/CwPexj905CplfcjtNlw8nv8Ff0HJfqfeNUd1G0e
EPGcr8wHXa1Eht7yWLVQY/dSZZVfbq61yNChrIqLS6ciGPC2gI8uiXsDJWFk41I7YLByU2y8GEBd
DZ0YTd2C9mPokSS0eJTmpXnFxbN1OT3VWSYA+2xbQXOq9lI9tR3oKQSdZUkvCObScK/glUMtQxVP
RHW5/v6bOiQH1nFN7/svI9Ch6uo5EdzDUfkGenLH7lASmKyAVKwK+aODZY6sGL2v1/+/tKRLMQ5z
d0wn9zzyZhYTRPdHdbkLyixVmvhXJMQuhAsJcbe3yBRuC22Qpn1yWO3fYDOC0USeqOKgNxioaDOt
j5rIFp/BBHM+9tnSpiOoMhGaKvjShfH5pmLDR6iLdf6WeOG7/U1JkG/OMkkKytZT2EHcfo3peY+5
OR+e4qlEPnF0Ht2uCB1YB9RcC8FSDvBvqgSZZw23SwnIYFBJh1m8M6Tc6EXMZ7bMuy6/nJgCuzNQ
CNYehwhV/m0Qg4a8ytElx3E7/nLyDOiixmlM7tcgFLqYrfmSRqptGySEHYuFf1s4r3HJfsbiT/Gc
j8xOmAjy6Idt3rRNWvUsvJebAVdFWh3PGtsjVkbjFESUatl/e4GXFMwpT+KPkcWZYZzC3BiAVRbi
ftTU+HD7wDkZ+ISdF8o/Ab/1Eh5pNPfEdGtopLYsN/E2/blOWsXsKYOVRNN8Q5AKuhX/ssLd9/ed
cU7B9t4O92K0fGUAK47ArRjwCYnNmvBEoaTv9qzikpD34paGy0yNLhcqbH9Ttz14mRYSeUDo/KMp
dt1SF2JB1AeWCF1JA6bbJomoV9ovReDl/0sBi/uwghutNIDhTv1EDXHPKpPDogCmtRugThCDiSJl
ze0bG7AIQDfDax6x1OKyB9e7CuXIXxvkhVeIpdJBunVlBrcoAJDgTxTIi+CQ6vOxv3y6osbugWa3
/71BbztQr4/ah9EHaVd6RgS/bzfXSfvWpA1Hx3tI1e4d/k5SQPquTJumB7Y0ekVu9nd+5s3cZH1s
O/lIYK5jzvwRL+7TEGYI9HwqwMwlWy6yie9+KJfA+t6yUL2Kxgkv9dO0d9y2yRQv+HPoyEvJkjV4
3EKH9mR0pthlMLA1e4NhTTcN0KA0kSMYB/8JvpyPbg9V8aWguNxNI9szzoqSQVSrAzsiA22oG1Ax
OrnClJrPbKiRsMtaba1/6hEzz6E/0DcW9t78tCvOxd7RmYEhS8jAjE6alT/1amYm7dCEV3BK0wNv
ho2wKmfAW7U2kGAbNeEiE/np3bv2vJiXdAxWb/j4rfHgZDHU/1RAHafskGwdtx1gvEMS46SBuZhn
0up/d9ZZw9I7vT9aPNvYQrJU8NQOxHfWyIqk/S751Pgi0A2mpyau+SGe2Rd++Tx6Egl3DBlW3um0
Ff3QBwE2KuK+ly6p89p3tKvSAyXAYs0dFFeISbdSef+UYg3L5h7iwoxcYf56/yLO/JRFPzoIXQMB
V3vPv8H3/Z98tqnw+ajkhCcNNRunIw4QhlfiHWm3Eic8XAqhfe1U+Nq2OCAValEWZIPChckPSz4y
3BympzFeFPh6lMpxlUg0Ca+Heed00qW+EfFgSp8QkDDUr930hurTg7SAj4/7prVID7XLqpJVNyTC
fEcrtWt87sIDdaaSqRBBLZSvD88jmK7kqBpjJ3t1BnG11u0FIPAStg6y2EL7vaubtV7ZBzadwWEi
/AeT+FC0IUjZSsFAinNl0DaEEncDv7X/t4Nb+oVmEkbGNhsX4sSxLkeNoOGkFcsaz9umJT1sZCul
5vgiMh6ZoHwYjgMtEuuVe2RZnIYgVs3D2/sj/FmaMujZKe7GMmDVEDiRLtxzEma8HpzqdmPc8F5e
QhyqRR3+YjAD9Tvxg6+OPrZmUDxIawaQJzt6d4DSymMe86xWpR2EyDQ++eN5lXsWZzEVUR31WHqU
UFUy4u/aMLIY8RZd3/4JySI47eDAhQ3+4008j/5e4sRF5ksYBO7XbXRWy/IA3s8LvxmL0fKK2hwp
dHT6vNz/m+Mae72nAyOtxY2anNR48jZfE1JIVXSkZpnO4fco+IlynQ8lWnLGFq7Fs0bHbE14Y0qE
/kRwH+C3r2BJayADmAP3/4frugfzIvJIbTj8HcD9VZSkLJo5FGYhQuDkgtRIaOQrZQkkbdQP0RYM
I/1KEGht+o/A6eAvVp/4aM8ZJkcaWMrtPSojOQnUjzUfUlAxBp3GkRjKgNFkgatX+Lqskyt8uKwS
EF8gUJigZndqDIpnhBxdZvkwVpfGVr2n6/iMQngCb8PpwrgoetHLVgY5SmXgejmLH1WILooGaQWS
4HqnrxTLv7V0Gj0Me2o98JyB6OXO/vjmWPU+FSAmu8jyR2orDJsJ4CzUBUme8RwN4mvhJ0jUgVs1
Misge3x/9D51MjDQte+KkmVLiuHXrCEutwxzXb1ZxHa3+aZPcGAzDQ4YKPKk5YvNuPnArJ/4/Nmu
ba4EniD8XA83+cWH1JAIsxThIDFRe1ze1DPt4inyqgUUrrkBt5HwOS4oNA1tmlt76nqsXBPG5x20
ztGRR+uNfCVXbeq0MLvFJbGqkP2yetYdL5O95vEaa3aQrs2lYnSyUGvdmnRsVTe1GS13/LZkrUNB
j7XcVKMIIpxflbEVFilxYTn4VYoD7VQhCJatmPJRucG6PVjrqjQCwLC/R5USviMvgIR2TjS9H+gX
wzCCmkWR3DKr+1WNULwyonHwDlGKdHSa1/OvGFdW+bQK2l+Jaz05lparQcMzDKjDtZ5Ssb42dGDf
JDiryfPwUzUo8mwfSzkE4WLLRpPCOuL7iV1kEUFb8lsTZbzPHQjmhkF7HhdMqV7hGaOXxhvAAyH6
h769Lp1rlrJh19EcziPDApbdrKVQpJUxEyb0FzRLLVcGF9V6ft9/NV1VAmKXQtuc514kvKqJSRIv
QnhrIhMdo/Q3ud4XCCuQUrtwP++SxQdXw4njkZDYQOr0vUOjwiFX8aoCO+BB6bRKFIy4rvi9CfBC
HyKiZnzExtrJrzzJ8V8fDfgkHM4ixl84EpIHw7de7ZGZ6VQvcpTgKUEdYfGRl0DjaHBB9hvq0cYu
l97zVb2Fz8JwqxIj35EUT5+oAzKoFSDWPvsu1C8fY1ygI7i7c0Cxtk/Kn+VId6avh0Nq/6us7hmd
H6oXtURqcl1VJFMBbNXne+3BbGEaDJ/kzygajizc/3x68zIyPY1BdtrCvZPvhwdIQ2oSuB8Z0IWg
KlydZePnCW6KLhMLZB+iJH9sZLOAJFvgy0nvUljVqYEkSRapPuBGR0dBH9asoXC0a9fNZr6Ex0ek
bKhc9CSoRW5pkRHba3c4dQTlRvu+bUy+7ypwlKMkcaXOzSc6zTPSRmwglbiPtpONGqcxnc3YzDgr
2WhHY5evuQK/WtZcgw4y/wVqtI2gAFKgle+Wk9MFeOWc6KggoxOk0SrCQsdcXVY/gpK3a5Bnkr4q
uS/deIggJqPhvwAm4fSr1NYmgpkbyopI+veyHJ87oS/sS50OzBdTZJbRLiDbTDT1SDHikMon1NU7
HDtHTH1FHOhdjTxuZddZBFyjFP+YUclbTZHYwwlPCSQKHPW9cyHohXfZBhP0mZzkSjM4ky8YK9hE
1TV8EvRCr1+FFvhCLYdHrFMx/NKSWqnwl03YKHvvxGQseifpFkKbLtmgKoxaAiUSt4ZAXI8DlVpQ
y51s5jc+JKigO1O1lB2YS0dj65Wqi23pa+p9Wboy6o3kAsvBw00ibPZHPPe+KWxG22tuAULDeHxs
BB5ohD31tSduqcIW3DClV8uZSBGqk6wncwpo1QYtppuUA+sMJF745/KB98OdfPxv41lu6b14Bd+q
dRL72Ys9TFACe6fH7hzZUZbxpjSdEUe8FhhIZWumORspl8d/LsjSm43haH/dE+tFWDi7uHjagCFf
I0hQ0cahcoaK7yB0hcsl8tKskB6cyX4euc9cIb5vXUJfgT5cZKOML1D6doMEskefX2B45NSeGKlf
ppr7YQARWvy6K1EVGm5fQfPH/vBG/VSt3BhS6lGr8VArf77B45mBcKZjJOp/bqrWUfXQcxZ8Kcdu
GuH3XXcjQVQQPFH3GbSABZurwmO0S+vS0gKjUWQwdpnGRZNpzj2Vy4uptpU4/3FX5Wo+gQs2A9mp
HpJdKSeUaeoJuX2awQKGfU8Gwfvi5QDmWkqwxF3Nlr4oel/8hylKZhTGocBmbJ7oZUt/P9T4EblN
WgGriLxqHxDArj2KDWnlFDPJG6zbPS3a+YkuOnm/c87jbE7yXRzfYEa/mWgxxDrJwESw2RpDc82f
EysFgzwL9ZahFChEb3xnFwNtJTwG9vmuD1Kw7CyKtgDVBHwDFVd4tJ6l0+yynry6GWS1oxc01YEp
BN8MkbIoNQA30fAhMnp47iQBCBsMOs3UDC8IYwpT8EzZK9c+/lWyMI9EcDiBP9k/CUiJ7ZOtXvZM
87KhW2LFOXyfbd2cRLb1G0IyU5Zcl1P64FQbpKjrdIB3farqJwkxOiiEKMQJQKsgOg6JmIg3LREl
wxFKJtLJxDsUEyNWkJ8v9YTre+ArrgFoeIGKaTGCh+XAaJjEPQv6PuRHQ3v808E2JR+VAnGmcaZX
S6faIpfztFsa19nlR2nW7uNPG9Il//MBoGK1mCJyWGcbCTQiCL8gpadrE73ifbb0D1sWLc5LTus4
DC+ne+YV9xoEJcAeyobhNhr12A+J/rt5V2aQ+r6azYO4nQmCZ6lA1jYYPG8oOQizTIUOJd2fACDO
cuqAQQCQ7Kd2xfHga/UbrCArHQyL55ynnJ/0S6FD/OLVDclHir3J6am7comooUY3B9D+zBQsV7Uo
MwNqE9MxcSjIBqeyvaHaqvO/0KZe6mGvVHAgwOlxlPPTSYLygishJIAQDE8aCGPDaq7hy/IQq/be
Py5bz+ejE4TQFxq2kcQI+7074hEGyCoBCIKYUIAgH7rgWvshcDbyCCmNthEah3hSvVbH3w2s4wj6
tkk3GMHvA5B8x6Ze9W669aBJmD66k/bJeHHQ0lc8LR9hvbIuk92E0ObfC8hDWH+98NYe8VaO2Cb0
14Lietv5w48MpSziy/R9maHR2/PwYPmN6FfSf7YItCGJhJ0XvjR1j7S6RMEXIkzSZXUy9vhZ20Ph
53l3lZJfH9YSpBhwb0xuuLPVThosvxegOb5XdVy5UleNhIw/oqJQMRiSMMLXevYP4UzaWc8AskTy
pobc9PykSdMtt0+Du16Ix1GZURWEpxw7Euisg1csFbfwN8lcLsHYJn1HrTbojAdnOHcx3Sk2Pjen
Vl0hOFZafHtsNdEdwbBdeE67GWuGwnYj8FLls01w4P0MfcKsDBN0b/DRyRAVlmXg0XEY9ePd+LWE
2BouAfrOh12f34yGhhqkRgqVf/onrmbBdZXd5gB6oULaSuukWCUuOQ77rChJ/RREqby+imDmi909
wD80Ewr+ufv8tQFFb12JGMU7VJbUU0xeMD30rdgRxoq+ts9BVtql9slCzU5Y9JsyBi0xGTNe/0Ta
JWZ97cpKkiuL6YWgYuPAVlWwlvoJJGvPtdbj42Dxnr6+EfF3GyF6xF78/qZdWva1cRAnlheIwAXc
/+mbCYIlfpkNhwbs8HCJ/QI4ttOKFpAYW4iAI4caR1rF1MChJhtnJg3/oDTQzjZdq2xxegqliTVr
OiB6oC/sGx6pwSbDr1Rlxpst2lAe/LSOMwxNm/6xNiszl5rBKlrnVi5d8AhrN3jbxp85fpltPw9m
f7CB70u81XqU452OlBmzvCOx2n8z4KjQS+uJTWaDfqqN7PARAAPB5IioojllyWSKFyf8SGNzfgN5
RD2j+RpBMtR2DDjwyQ+2w7MC9ZIrqJsNkJjoPnbIEmu0dscDpFmEJegIjhumfigKT+h84xz6/PzJ
iZCz7U0qcObVloNz7im8lpTVvRQYeCZKbqRDwqWmEbJ8QWsy0hhnn386HIa2SyXAAM1ZU4aaWtEb
ftsdhBdyLZV3jPueryg2GkWEeFApDIveFvxMG03nqUpJ5AiQ4+hlmhdOpkH7SImunaVEz4G3W+JQ
GVC1qXc4qGR8lLQ0Cak2lay6IVQkVbHDBqbiMOL1mehv5zh43Bundg6+d+ZRK7BOmC2WazPVaX4t
ZRW8vM27rpHuxwhFOUNvBS0AG7NATNoR0nPLdKxFERYvKfOKus8XqCFYjRJhSdk9fYCyVgLvovsB
nX0wx8ubT7Cfc2e/iQ0fvch4rfVsjPst+FAUhohrQCFl7sC30ge3+ukGIi39aBeltFFd7FsHx8Ww
dgCibBN35AYpvDIDLzBUyhyZE5FY+8j0+mc8Nf0hosy7XaMcJdYkOZKUxBiSbv94MwvZc5Cdnbaq
4SLD6yRdBSGBcc9n9BrBofA5sE/rpAun+RY3H9AREdRZ+XcdMH9xnvj9LOJNv+lq6wXKKfT+phdv
GZYWwHDqUeiOMTldEhEjIuwiWWAhMzNA3uhwkohztNPreVsGLnxX/VT2iD4iKnWD2KeABCJNdU1V
tdT4Taq09iGo4ClkQ3lwIC0i924jeIsW61kCvdb6YwCvgkLcy2euu0QPr+XEdXfQTiUvfXv/Pz9k
utxdWNrk5NXpMADyx7AqexCB52/3jZ5bjwQiqCS+G4nFhVPT5xSeE/0KC+AUElGPEbyEFJ2QiDCg
DT+Cv49K9RjPCgP6py4feHWsS8w95KZIs/Vnb08OBWPe1+uZk0wNCsxnQBEI833RywA29Y2lBMdr
AP3OTEUYC6F1gKe3EFPp58EcDNrtO1c2PM0U3HoBhffRmVvrn9YjvyCba1TxEven+sMlOkZULW2Z
izUl3rOzrhKR1x6OMyItOF041OR33T4vjYLZ5HX1ZKm3CHA1mdyy7TYvzOCKZ28bOoBjCLLH2RE5
gSRaDwNEDdAHt1Q5l72PTHm59IPhnfPWbSAC8iOcU2Gu2auqS2NCOeaukMtOGvUFeW/wtbSTFUYZ
C0w7t+x9AwjHxdvC6YYLiU5tG7VVEJzbdZ+NnUlPjpwq3hCb/I2T7WuSXi9cvXAjMpyoa27wbnC1
FyYUl9NpuNj6H1f0BhhPv0D+jipTZvZY/k4qFXgR1z01XessGPLvhRNjNDvx2RtYARuinYMGwpT3
JA2ZBTiBj010y3K8OF+Fvm6RMU3ILsrKBzCccUstidGg/ZNQS/33MSlI1wy+ZoRFGPxsxTCqeRYk
gZxgYHGOrfAV2H6W17rp58Q6F5MMd6aJPqezx7kBJFT3jq41LCcXiTRsF5HOV8X3lUlHZOGQNObT
q2rr1noijQT8nRu5iTME8ghbq/k2WI1sfuwWpP5uhbfFrnGKDGE4naccQ5QvjKYSAiplK9OJ5LSf
025+DDAFL8tHgwI0ti0R725W1SppgAI8cGUf3VY9v7knI3AhK1XJjU/IxXpPwAvMUcd41VzQ9HEs
opBAsKCoqk8Tw7XvY+qqodaAIV49tax7ju1mMlsARJ01LdvflcKG1uMYfs5BsNjcqy30Ph1vt1rs
Ed/YRoHsDtM2oagxq3qtlWfIcYqp4Tt1/LaVj1uv1lMhB4+z57M5WcGqxmGupIazpOK0CmEXj+VG
kv4bkJ1Q2LEloupDCMmck2pRyKQDM5fXKVQAYwTNx+a10mNTLAcGA1QeB4C9hwZE6bCZrd9G3pjm
vWkUeelrjr51uDIoXizeZzY6VuIsAx4o2kbLwwTkixGThMxvM/fdBapb5Z1K/TCQcWvZk7Tru/nZ
VYm1fI2ijWARQRicR02fcJVoXN846FMUZFQpo5WW11qAxMPyqT+EO/Artg5ByXZaxMu1dCkU2yyQ
hPdteCqdr0OqWT4+clivrORTHZI9So/+CZSKRwqOQQBM8z8CV/wKyyaLylhfKWdKoY3hkk/RbAPT
as0e0KZibBIJeqSahkhDfviHvdBXKK0P01oFyPiLQLqqvu1YJ3bjJVnX0v9pJBWkzuhLqDGcz8XL
16lGGyulXFQ8aFdVNr0cWa9wHf4F74uFX4OMrvuY+85XZXPLOhUmx3kGZpkiQ5MLTm0ptZOEoZQl
QcnC+XUVsFwyx+E9sx2VE26NpRVpt6uY0oiUp4lLizYxV6jJ2rA8fs5PXdf3EtGVHLQfFSN/El9z
BquIzs1cZzu9kK7jbXyy4Dd9n5gYOz3dHd6zeGMTVpP3ORdaP0MJ9eOkns+PQyJD/OasyRfS2oEz
TCwrhZup0/2emZtEqF4cQ4DG/Q++n2P/BdcrMQZazXFpx8hYhUUZXkA8xvVe2X7xvJh0f9IgmCte
+8/lC3WJmQMlpqtTFm5/TpKxpQ1b1MsAX5+jahBlfDpDP8UyksMzud3L7SYuDI4Bmcligxu8rteg
hp2I6cbD4LBf7RzvtxQkQyabnK4wzdIgjluwLu4jhHHHwJDb7YnlqMWBRhDRpm16ZyK2adbk6yKD
mhC06TkxzfV8FLwqZvM+ucUyqp3prygAZbGmonpArnOVUo246e/vafFbLoHW4im8w65xZtuGAJxR
XSauHGKzUANX+7cgXUQ50AtQB/D3d2zmKQ7CdY5+e2W5kCu6lfJa6gkBn3gSTJgsT3cBAmliajkJ
YbpyTW3A7g9RWOiXiJ6vznIcOOgo5erNrzRkrzPwKaHyGWnMUtFVIf1XPzxYM2GPsz8P1MiQgHz7
yxJkk6yq/5yjSw3lETWJuZ0umlQVbcelUsr0GOfTepKvksKVb0R5pvXOsCjaNATVeMwmXirS2EgV
aF2Ta2tsvPFEvay6vno4W0lVse6tLmKXF+QmTG1p7Qw5Fi3ID79wjFZoe9cZ4yVYUcjcMLu0LbIH
voQRirS8KuL0cH7m1OohUm7O8g6BZ6/T8Rz6LxnNWp9Wh6IczhzfQJKQv3s4cJUzDQsbErEqsEu8
KXQrtjx/0rKnoZ46WUnGghYn5d8S2hs6pHjMrCSTvsOUV32RTjKIjglQJx32GmLJaLlS54NtZJnl
y9VW0oiJJ8TWenx3zQfbaO/l1FeqjsJcpdcxFzZU1qi4PHlnqXvPHmXyCObRY42GBrZxvJ45stjZ
6C5Rqq/l42V3rINHFPnQAlSXMgedca6BkfWzs+md15TbIs/rr5ueoCyK6ZcvL2g/zRh3UcaPaipR
XhG8Y2p7s8jblG7PlwErlPp2lDu++ZjjXJyr3k4aIWcJRZ61K2cJl+Hk2jdG50eM1ESzezqGS/g8
sGYvp8R/n+L5utxDViFx1TnMb0UbAc6ED74dcFEb+pE6TdMBblBkFT/LMwwVJDHhHQ1g+Yz7NxPI
j01TKGw6DeVA3+D/ODEu+fQnfX9Q2n4bBXaL+qaPptN5IPjjNgTmPu7WSajUAVCqzAJG80h+6MW/
kXXmGNmoFY2L8nSKmY21JVe0f200pVoOF4u1ZXDDpQHvQdHZbx0meBiiwUGvdzjxPQo7qeKqmfT1
uLffo2foDPdAavGW0JXOJr3USrNWLz75Uzm8maK5iXTfgBr+cvpmmgp+goYJfn24cEGjFsOh54XU
D7oevgASEID7iAftBqDQ6RZlZcDRaM5ebUVcY4pOK9/pW6LrOUqUCrn8mtsMzNdNTYZ9F2CjwNcT
xvUuhdOIp1xh7ldzIhMWn1CMWTAxL16J1GzmkaOAAzpC8/CU6uYtfp9Jr7uM6HfG1KJPPlGVxwVZ
/W/i9Be3rngJ8Y4LVi5ZPt3enPtPlo5sx6aCUnFSJGb41mQ54rCMjFUdjAnAblqCG6Eq9nigS6Bv
OUAd5UpbSbYJX50eASdt1xxy6DMrB6K4IADvLr1L6QO6iHmwKzDtdLj/EiGuG7F0MA/2ND74wUJi
UBqk99LZRw6CxRwV1SSe54gIA/XHdQiGowJGH0U6aJ+B+n1GDEWsPBxIMXa9LodBoslB3PCnOJ3z
SN7s/KW7Gy4XrJ+UN+8HSJN5BydzbB8zhpqKRNjhoh5GgS8a5FZ4ksn1nYBc6c1SlSp61E/J6UFh
9pl8vTDFliAx50GhiL+OzI7cPt9Pe1vO4dr/0vPcugn29eJ4fzsNlOB5X+7UBbKwtZrw7PvgO+6q
nk/T/8EMGAbhXJLUTP+cesKvjqVGTyul1jP+k3lke+xLneAfTX9P41DIzG40bL6LJg5rMm2B1LDu
bOYiZP9dqiphPeep/fgce3YYbzwZ/Upcg4I+K34vR7BGjUP7N5m78bsAaL/pY4kUXQI+8HsB4N9k
9nMTVZQiorvRbHWTjMIfgiJQWBt6ioX9ZFoe02RBm2g5ueiuyd8t0/Eagu/H5aowi0rHLbQWV1+v
CI6dLS77xKobr7tfmvWavJLjyMaatIyTwAbgIRY6hoRXg5TXit6wyVxgKX23XsVJajUunSsRdm+s
ZPsrztXYXZIGNLoWRo46AcEUazgHk5P0qm4MsDvGTlaERcTsl1rXrynJIYoTUAVTLiYLCStHMNs1
B7Pm++tZqPDydmduKXjaQNMLywGJizWCEGEy8xHA/dO78BKmNysYvTw9j9LPcoKkX4LwL5YsG0+A
OFaZmUJUl8OE4XovjA+MPtV/KH2VRram7dcaG2jwt7Yz0hFFcZa3HPXzhHitA/lsXM3xRHAmEiwO
tPqTHsW13Oc8nVyhNV3p+rAUuD+70Kmm5DpyAGbLUxDRSZrMUq63tY4DeCbHStjJ3h6YrEkggKJL
9FSMu1OOjriWWWO0lsfFMSvgJAglke3PNpWXx/XYdY7mdI2MQqGOLNpMboM90WNF4M5BVmzBBZ7+
Tnc3tTzS86SsDlTiHEK6XhVhwGl0cm4GSA5y7zogl7KJkn/UKwiZS31OKssZ2r9HzokFL4sq8sQ3
KrYe1Qz/tv4TcQ8BTH90NUIFEFeBp/O9vBeuenRo/IYvm8u7Rll2kXkkrhszHbYeg128pkytUPes
RxMbGIPrxzIoyhmvZPtwqiO169y9hPSerJnqd2pSasa5tUGwbrTtwHbJbS14XqMLoEu0wwUHlsif
/bUAnijrcorJ4oV0aHjo22+JDekXmk+gHnv3U7VZn2cpCl+lfzQJ4/OUDp7R+3yepZfr3NHcVZfg
oQqYTaKHu41E+utd2nnyHDmcTYnMmU90Bb1KgabwBQbkAtDWAAcMOsHsokNHSYtcXwVbTOyMsm0b
lWU5Y5/Q87O3VFerrHxpA6ZT+BOSyGhK1zUKR/2jBoLJpIFbfwZGS4irYPxTs/XCLsxoYQTlI4Kx
PMXhIUtxtl1Iac4tg9nVRcuOfBv4y0TQdqS9tZ8Ld6klt5C+zuL4w+fnwfFQtThCGsmHjf3g/2nS
91cEMRC1314ed3E0C4WWPU4ltf0p5JHdKKEF1evMP202wpGXC/D4sKgvGvlv9805Hn1MoaB2fvSd
dSwxcZlIC4dAAhtreUTCVaUKPobUZxjYBECVCcFCPHYSqJ6ogKn5usZJ6dWQc+od/8mVtD83y9Ay
ZYxT+g0joko4B69SmJKERJgCLpSY5YF2LY/Ae4w8xmPo7RGTvYN7Ryz8nig4Z0zi8VuRkByyzIJX
1gLtbSZWWjvOz6xh7TasdyMB5AzMynS9hr3vqu5Frw46qexc7pDNtL6ZiZu5bYjF9qFd96O4ogng
RwqpJ36ACEWLd/id7iftDnmkb6zz0ktgTxOrUn6LFH5suVPE4yJr/1/+Fkea2KhUm6tYdpJ+Jmye
w4NxnogeP3r1q2KaK8x65Ot1guDLSbqgaE+X+TK49/rXN7B8Tg54wl17oXTjAMx8RrkO+gYZ6wWf
KhnUFrhy+WRV/cr7KonsknOAMANF85iOpjN6vqCW1WQdGML5F6nffys/I6B/2+BTJooy3CugEB9Y
Ew9zlSWI698mF8ok5yiOtlW9wbDofG75MFWKppDUI94DG00o3j+Hwoo7YYbhI9O9IOZ7AdLtvJ1N
CaWb4K5qQd6ybU7+sRe6hxDZPLh6XmfYUkCZ+wlWQVEO+I06TCxhJOJ90Iw1guYLMgIFGtZPWmBG
I44NmL7XjTBawi5LN7o5xoAylRTBVF+zg4TcUD8B7cGlfbl66wkQZT3STJ4VKOVmiNkjtR1owBt4
naVfkvQtmibl6wZmiqsylsr4d2wYaB8Ou+SNvPGDW5BuE1wFQsn5Y8NwSv5I5caX/QuOMdlta5Gl
bY24am3XId+e4XYA9RUNlblhHdqsySpr1MxCtTArRcjNZCV/X26X2IxlVH9vN9bArtKp50THrqYb
7bEUEPQxpKm9eo9EsOm4duFWCaOTQk+HBgtU2tRv9Vv5e0LMKlMHb01wI5fBTYhm/k449w6QdHN0
Itj/9uqPoKQeCsod+IhqY9wCHRxpHj6hOlHiCV9V6cy2VgriuHlR4C5Q8yYh3DQAFRR6GWNTrKsm
PBG4RKe5CnjTY1FFrIY7UmjzdECna4jb83VX4rTTI2N1HbWH0ZfTN7XXdTiN6Bhq8rZ1YXkC3lqV
VKDzDJeLjN3F8Zz8YKjMhQqslrRgcahZ42DcQ4/rODYytD9eGSAUjJ1eKGavSyd1jlWCARQvFUtn
cvERSAf6VvMA68FgjkPQQHg5wDjt2lqPkogpHUrHlQSZ5AcWMeOVnn0V0MVxTp7xUgkm3ED5xXVi
RoP3vZchiRRu/EzepfDVoyLGLtlWMCu5VkNNZselnq4TK+46+JF1C+YGTjesfQTs/0uKxLjx/blR
8g5eZqjxNMkrF03oDCMnCjaKjN1I+A4033xWPI1vtLyyUFW7BhTbFDTifK4mf1otFcdjVqYKRdwk
d9IqnDoD/B9i/afXogtMh2kgAX/FZMjoDbioBQxFhCtHKB6spxA9WpyvVD9zgV31zhLwSTr5cDt/
z/trxbF1SMrY3oPNawew0UA+SZDtezoaJ4kluGGtDc5oSsZxWnLKDY017gadgswA9gPdGLmKUoDZ
60/cR6y8O54tXLVjA0PJ/t6dicQafsWksS02jYG8rCyHpfJjaTW9/q+IbvTKX8LFHsqXIvgn60I/
x7atuBLFKl+4gADrPoHxZsvuLMq4umyHgNJEy/HdZ5QieiVGukc3pPD6MPpFLNzC0fvapAlZleil
vP8/m8ATrH6+0de3/2Gh6GJhLr3B6+FEQpc06McHnBoC4NVTinAV4q8E75+pFOZ7Hb23XilmjYor
xmU0MCHJGw8svJo4fH2UwvS+Jelg4qT4hXCqUrFsUfVOCTjMLjpEZlxN7E2QbC6wpHHLWjIQHdPw
UJ4CtgfxW4cmit9lTI8aWRHkZS+PSccoeMvEGTGMLULZgiSem3pWlvjALW1KAu5eRoH2q2ydQ/at
xrrCH6USNNsjOPqpyK6F8ADmRrP5rK5BRiOjkt4U4UtT7UQQBYJtT6Pl3sJQpt1wh22Ggm7WuhSd
kZseQ9AgnAucPDLBZPyZqX/xG1pcHn3y1dm5VG0B0yinmcyVzV2p/j2Y6r6wY6F4JVlO4E843O8W
bNkpegZMAhDG70nZI0NtiytPbM4OJXxJ4SEvKUaNdC5fO1PgKPV74Ap1qLCn4Fe0ilocAnaHUPr4
csaa2SS2fQAUACN2oOLhrp7IcuRVfRU10PYW2UfDKnJjpvIvD3AHTbPHNasN2o1yUdeijZyBwX9f
r+16AXfOuzroh9X3gNTLuqpX2Sq3qbP+UXgS3QAavUNBYgJpSf4lGg//O6o4e8iX1LJKTNvKPJlW
dxBuFn4bRXMhQhtXPg6xjnm0cQ4X42HpO1Afe1VisOSQuR2sAmCDqzBpacMDiOjFH0KHQT7gm3LA
gJ4OHvH9JhlHj5JD6OmlZjdpdat8t30jU1nIfDe01PCRxTshswAyuIkRkoxASKKPLlIIzQ65Yp6f
a3UBL2Rp2sDtSucXdjiplwY51bJMfqtdPo2xRtCngEhPwtxoNXE5y5WRiY4fzBpZJt5cSsX4jtuf
K3I08kBJWXnDpinwh0ZMabNWo2A8qM+I1ORM23ES7NNld2IM1VqW/RbNXkSTJFp+NZTWH3Zd0NyP
tVpTjVi8rp5JRDCTmvujhc6rwNOc8Rd3I0MWBX1ZQtU/UNRaFrAgHnUGPyAGpODdc4XebEgUUEs6
7qMElE2xMIhlzLJAm84ebexmYlZHSGGSZ61A9vAm9Nz5qYlBdswOnLNwv5I1r+kToJqmM2KD/MwL
K5tAzKT92xZRu4ftqf+V9Kska2cWDYz9rcx+Rv4XSF8GJMkC9VKrRdnz5yLMF+RCYRaZ0F2fYGRk
vSZBh289uYnhytisQscJSPKbD2lHMvfpp5yZ57T0Hk+KaoJ9Vj0kHhKl/RzdGLaVQP6Wdbn4Wn5n
U0s8PNxnz0UIeYDO1lZEkEbus/wph5NMYbwYnffK7p9+dzOBYXoyWOcDp3Z/PjuBCSCN2SJXZF4Y
tJk9IHy2BZjyn8UqFNSjj6pxhJOceaqvv5iux0Kg15dPt0x7HoichDs1GccUtrn+SikLBw2Ce8n/
ecT7qy3yM2daPJVcD3fdWXScy4tCm50rrHc02mjnFP49VXBOT+OJuEsyjRDsgsWL+5l+OoEnKvKb
2JN7jDtvBc6lEBfXFECk9QUBOkl/ak9WbaW2Kf/bR30n9dlxWkxabHK6qHBbt6wM/zFYS9JQFxNl
onUSCPTptxQ1HOstyw/p/pdau6fQaFdQjdnXOQxoEdtlwWw5i/amx9+2wzvXzMMXnKEbyN9/g8lZ
Z6Uwj8lk5Zyzje0Lv0FmDwBLbo3oFdKuqGAVEoU7ng+sdF5r+tDOH5ebCNwg34d/85Lt9dy55vrI
LJxZjvqvjhLFr+n0a6npnuE9iEFxJ9JnO35yXIo+8eSvgswk3BvCqf6WKe3j2wU2D0eHHq+7NHmK
JfdvbLRYUXlhRx3Q35UX/OcDOVxhoaz8GS00cNbhWCFuYTqkc/es0slj6RJk+GNhcU+uwuaPG+I9
o2qYlKY2X82L9pGoX/kCPgSaoSzzfKEwddhyq8e7aub8+Y/Rr0s4Uw5oQEBi2mPeQktS15z1FAik
rfQO1E/Y1FFjqzEWlHFucF7qvGY35ZPqmLz1n+FHduYSjyPd61LANFml9VA2v1RUHot9yESHRVJp
wWVl5L3gm23ycVOfD4yTJP4EqDJDpD+FGq7V6hCGGevoadazprS85VPhRa+F0djFTOMXTyDl8qN/
l/SOkGewO/K8uy9nqlB6r2uT+vgpNST1R/dTMehWIp1CMbWPPfSe+68zesAoaC4TVTs3ntB7nNIk
4MqFqFVgaKSS4+uxLQCCOgp7Yvdn6YnYmAMEfsa6y7BSmDWAUpkRXARmgGTv/cqUZuSZ3MVzN4X4
WRmCICeKOa7Tx8S4S6YZun6BBoiWfJ/R7/7NWYfsQ6c7eZFAf/FnJTHwN9tx8xs27VF5opmx6rnP
VtSQQPOPFHYmRcp02roBzMcYU5e1c0+3bcN7sR4hZR7TzwMTYSO4xheayYHFlu8KlrP4hYDDYpFk
TcA0dcrJg+W1QAt9Ce2LgaNz7MmMzFLXFRFIB8u7KZaVD2A5MhWkCY8zYv/MUN4+4SW4kAw8N9Hl
ox54Innw0Piu0I8dr8LuSE3MONBkrVoMj0iHVoRmre8+PQruD/NtOuVAG0pO3xd9Gr57ImQZccVF
SrytCfae6lxfUUkYWNViT+HzHTRU201MTcpvIryJ22ivYOfa3851M2gF3f+MRWijv8vCfXEqEodZ
HYqKEu8qghhMlYmO2RLphmPnjvD3v97zavFP+DAWc2M7WwNrR5Jtxps/Kf3gPN94UOpgTAukV4P1
Hzt51FfI/9GCylswBFGuIfGRQCTtOM/l0Yg6wyWBBoyt3cVTJheGsUvtvdz44+KTtp2Kxuaf1Yvk
dE/MDRNxgltKsxCqEwDu/HJ9itSs7/BwgcjdZByaKZEy7Odbh3KPu0YrqJI7oBaS2ROAccw5xNPw
CVbVOonDxA0CVvQFU+o1BJGQIcxOAxWoeTg5eFiJFhkApQeNZMJzp3m6jLP6/J88yGWvU0S8jHOO
LYCy3MGGz0mfmRVn10XkTzxJMeJ/QzQVmaORSLvTXD85DXTRsq0/1Lhi//J3+V26a1/jKfgJ2aYP
E549TunbXkKODI44W/DdeAsgpGvnCn8BWUt0BOsmyuvUsQdA56WsIaPOLQN1GGww64WwKB4KiT/M
4jSv9k0ZiRPY2Ayk2HwShNPq4GtHBQP6H2TpPJBCf2hQI92KCjTdO+ob6BUJO3FnO1WvR+H0T8GV
2fSJRoefZ/8SYEJpNTqOu2fJWuSu5dXiTiSBYWqu+WpIdCfQxltQoGvmBV3dnEKOuYVA5C+dpBou
dAg+TVd4ZQ6+6aV/om7hOtnHWbZm/ahCa/lVgb1C+i+MmSETql1xjz7gPeKFqFAAae5GgF56WA/p
NGjqpDPGpFtUJ7e4+6AR31Tw3RrWRLiMzJcxJqwEE0dOARGH0/hnUYMalsboNl6r0UIrBj77/eWk
zOaIbcacoPwoBcx7GP7E15LMWjaFZp6hEX6aw/00wzwh4EfEUPLoTbD8Fk3PM0cbQ9ErLOBs4khX
YgVQFr9ONxNd0DAHulGoNgRYTc5npXc18oRcv3NV1P6LZRfMGoUqT9+Lh3aQmm1Dqpo1UXA5K7Or
mKOMiu8jua+vqvnvkLTJwscUL3pAQmaEpbF2AwamgVBnl5vAPDT3jGxnA6/MbsoxGZ86Ys78i1O8
Rvqz/fx2ZSH5BIa5Bo2CE6LZeoqp/W1tH+He/xiifFRlpcE06XvKB4Ad2s00aLbVozeJ1jpYcuNn
O+HvAPPIqBWz9kBiaSyrzFQlrMP6H68orts7J+0wJfLwbe9CgpL4t9LUTxoX9BrK16j90br/PWpE
6KoNJm8qb2vezig/Cy60MeMEqnSJqTUp5P+/aTzSPGP2be9eT6IIQ703OWcIHapIfM614AyDdeHQ
igvA+mz3iTPfMGO58wPSXAth9Si+7sJFsxHomy05Htq7GziOvwnLAsMsVKCvLn22IF1q8+dY1unW
JewabmhHcqvX2tnL0hw0xhxBzHzLyBF604QCh0CjoAw8tuE4021nanpAcxFj1E62IkXA51hN0ZMU
p5nYQqYNjvxhzEvqX/d5l0Td25jaFxtB1jNCWoVrmEAqgutexyj75sY7XWARmvP2d/OCoLcO6f/o
9RePoF7SJ4XuhQajJ/UHSVOIspOIZ3OJTM+nI5viawVk2AidCTPij3C/kdoxAqX1aufX2YZcQH1b
v0if6WzosebIiZZT0YNlf3R3pCvQ2QCh0z9/3goOe/L/smp/b0LgPvMrdYmsbcychykxtVkVuqY8
fTX41PMGi2bO/ULfIhCBnjxxTfa2e1HRHxditYatv+GjIDtMuAEdzGWCaZZRM8D3lxCoMAQCWx6w
3rWZMiKw+xw964lS95XxfBMfgN3SbvXlr2ZfXkehcEUvzPRiGtOw3zNOAkDsvBdS6QQg0iIliZdA
d6fTZyX9SmOeRzlhWfBGzf/DgqVkyd7ZrtUESc9fuPuxF9LqNi0IPA5iBPy3hSahokwd8nRAtt0I
7L6czLmUdUlt321aYzlyyaSYIBkqM3T8ic6soQsSAdMajzCbCywvkWpnkzFdQBFdsYXBa1N4HCSr
x1reMvgp24g6XISFIG3B71881X+KugksX857r3B9Bcp/1eMJNkGpJjqCdFff15IgcnSKlbu7ZBo7
1N/OSudbRrJ6Ptb1uflFWQaFMYTgt0V/EzPLP8L51eMKtcSnmJCDfM/s9pOWrjkK+c1xbVSh+w7Z
ZjWJUswOg9ravM3AsHKTahNv2jUi8kju2HbfyF+9Y0jVXYDj+ME+9S6FX9bl+2tjim0EKDn7Hv6q
seYBj1n6GIVHC1QpuEBmijfGikv3FR032n/+accmNiFlVoxoEI1laXcmjsfQh+TIttODuC04Q+mL
1lE5F/eqL4uYCb4T+ZHMgSSLgwAWr1Un+G6pX/ysUUKQkb+Yp3gLosOlH5ECjHZwRkIT/XfG44to
Wsr0kj0B6ekFaae/r8y+bwq+vgfV1CTcxP1nSpHcSpLRp0lmDD7cdvpzCScjRpHGAEhgiCRw8i0x
PGpMJCtF/TriNraRe/mbF4t0LJ68prHK3bg/EV+fu301QlLYswTHVV52acXvuwx4cQfUvkKovPW6
oaauoiG3wrAKMK+goAV1/YmwNXdOwLWxvcyKWKZIVyej1GlIk8sklZd9hsCXFkS8A8Ny/N9XoCgK
74TX+0t8LCfU7oOqKhzZj2ogXuS0700pPyz6KHF/oFa62nZQLFqEGAQ8ecTrUnBg3ZC/bh8CU5Qz
v42TzixPP6hZ5x2l2lHma+GXbnZOT3iZG11lYh54WkdCNzTzPean9qqLSplj1ydM+9V5lcFNvL33
LNUrVltzyeZkVFM06ihZwfHYwkOfpGv93ZQdVI4sOOn22QYoPWf9ZvE7VgZu2D3cZpsaVrQfpxjs
HhsxZEDHjvQhL/CLjDsqmwOcu8E5XTOUgExH7ESNdsUtoxMeBcEq1BY3rFQFSa/Kwrjp9lY1Qfzd
6fueBc0f0YvU8MfAdOuCno+P0TQbLIqzSFnGSfcms36lfK759p/n3TfvfMbQ/6u8DXL1tBng+rU4
px6RASmLFIR9fKqwfujd3AmZumAkLNFsA9lCuAI1cpMQ0mVNXSlpwQ0CUa+FCePtyv+08lC3IM42
UEndBX92O598SPqKRYtGDDNs1mgsG+Wqb+W+UfFbVqVTr4fnRz/dpDizZeB523B0knf2E6zcGlGO
inqoMSPeWkieL9ky9bRPtSTChDl1Bsn1KJubGMR+gUb4aDY/DSh8Zp0gr4I5MbOor/j3Wes+IWcG
dGyYB2fNh7Rv92buf5arGAYW9H9fBwhTR8idOSxF6eHBl8FqxtrnotKw/G7qdP8i6qWYoZmJHPnW
6URNa8S7VmKjW8S0QTegnvHZKtTrl3vmtbBbe6bdPx0VQ/xpiYuZWziGZf4+95DEVexfmbUUU/RZ
iz04H7cpfji7zcFh93Rw4IZTkVqWL9CcLZ5+ZDtW3Ua89ozZx4HX44QkywtCbMAaAaVGPblcjfUo
yuOhG8y0V61lLtZPnZUIfXuyDvVUCqIZI2sUEX//TuzQRAyR12bTydJz+gft4eFG0exySzoX4plN
hc4e1G2YQ6A15sTNbauKUwvbfXV/FuQTFIPt/dzP0wvTs10xsRnoZWUqEguUanVbsfZAkzik0TOK
XtDb4p1hGtiDXkZ0XLehJmnLLUCI11p6Yo6RrJqy7g2hAK4sqqCevUlgqos8YSDQQ5AvqgbFbFfY
KM+qNKl3oEXKY8nM61NsFlj7lOQ5SS3p7gEsPEGPFXWK6evpHKtvzsv8rnGWASXazgHmdMMwAxIR
M38tMCKui1jAHf+uGqokhJmjDiE0UeXDIX/8IBV3D0l4MvosoMbAZPHLtuXWpllZIR+MtxX8Gq/O
L25dtCCmDimb2n3QEYgPSaxOeh93gQi4FYeCFgSJcoMIh7LvdmFQQ+6d9wgUqAAQ142wzOr3pPFS
IdiLZ+rGzm9Qzg+Ss2vTQoCURcQqZhyvpKhumDbEz5z46lFrLveWmwITPJtw8WCa9HYzDYeK/BSo
Y1QuBmPdF6zbW1aMF52bqIXAhvOMYyWGx7EvMRVGCwDwHfdVO89PuMD6Q039SjwjHj+LFufQDJ6e
EH2c5Hw5EtG06w2fW2HIaKncX+Z2Z6jLIvDZs9BVlJe3onSYkiDRAY6Nz3Ru6e7Q24FnRwDQzofm
ZHcIU/QsGk6n0J3Fka/jBWrxNY8jMcKtheEejDFPj75v5f4FuYxoKkWL5WNsAau0/KrPA4yDSmVR
ckVFDBG/ONUkDInYVQrVXV+RDPrCUnTs+gmCeYiTg6EMrTBEhj3IGHlRfFgk2wbM+prFWhpJpt3Z
/7CXu6RSdnispuf+9TixD/8+qfSY49b/YphztgNd6cdwLDNopk1C1oHor9LCLX/ic4lvmuEtM88o
dU7r8E2w+TnzNEZbUU2clpxeCzkoKUY99YZseBl8/gmm66Y2x2tLGDv6AXX/QE+w8j530DSLanAt
CiT9lkH6V8Rg7vgEr650R7c0j/0Q/B2p6+FqvrKThF4BypJJsV21Su1itlOXys/vxMSz1gEjWaJM
jsbvXn8nQW2NkAF5bIRls+lJ8WPfS8a8VIm/Vq4CHri0o718zFXGPAW21Lqdvlzr9ZD47SM8vZ9R
c1YJ5aUX2vOQQqrDDj3rxG59ywV26fNKNzVueShkGg5pz6TFJ0xlJX+CvproLHuLnPa/qXCXOZME
bErT15+WTUFiQRhh0FnR67dptgMPqSGLtmu1XFDDrGndgaAKsmQb2+oTi1gMjQ3nYkmEquLPXaPj
Uy2flHrW/cMaAft3tsC/sIdc7LUS847uZrRRZmFkSrmKX27++8OBrCWOeaA7d/KieWpjzwfsd1VT
cFIrco/BeF76ByPmxV10u6wm4RQE2Etj7JAvBQGoyvd54t1YtRaHnILSTDd+s1zozvLCw2WSzVAW
pIg0ru548oi6+cWWB5S1IqKhfaheRYu2w4HrKUfTOeGjmTHSHxBRA2zGgJXPg9ucDvcL4N77u/HC
arhErsb/wn0nKhlC6NBD+K9Lvu4UbxXlLR6BbiHTLVBWdc6Eit88jEnfhVYOSFfIoQaWN1sdTdI2
L3Z9bngJEQ98LEQdEWzk/XpYfPE5fnac/Q5x8l0DN4pSli26AY6OsLh1EVRFBYKXkT9u83/K/viA
Z2c3PPMQ0KG39GVXqndza3KYgbucXO+XpODWHEPxs1Rk7jkpUMvagVrKQgVBkcKp+KuayI5im9e9
me+ZPXBWEN0Z2PJEGF5P1/XzXfsMnPBo/E+qTFhb8DKn9B5jsqK0Yc6EWFOfi/V69s6RWLDwUb0j
mlXVBVsIK4Qf44AlZJvNJzZwXdArTZ5oINux9pcwfSyKbTvd/72mqert8ylkjmvzdwSmiPXlRWmr
+YSjxldoU2o15lRDrbc0tfu/xsq6FdWnm2zRYC7sVu1f3sXmTE3X2R/zINnOH3nKr5TIGSbchaj3
6pz0DfRlPyezCnOrzYElOq4M2fZ4cCb85h+xRvN+PX5fwbSCrUe25NLiV5BVmNvjEl5mzeH6sOXQ
YgaCAg65hUoSd83N/dxpbWnicgoNnuEamyV852wp/QNTgKtJ7Hft78b8G/z4/qxXgPlqx13AUHFN
pLbBGIp11IMRP3x6yMr65hRFOpDM05epS676+mRzT8aNw+27ItWB6hNrH5t6J/XQI7/OA1TSKHIP
dCgf6X87K0RkJjHkAHqgg+dVyoVxaIVAkTG45ZwTdzFJuFzkpkETCqkOqKmlyvVqOtQmM3zSx/aY
jfTXQS4RwomlWNEs1WaAbd3Mjlp30w126pp1Iqwf7i25F1/z2GJPbovrzJRIjZaK+hvsK/qRSMCm
zOY1T+ma7Hl2hDM5W444eAEw0mOM32yEnTTDuB2ZNnaALIf7F3ZzaH5nY7X0l8+e+Z3PBmRzKVhr
Y2BqgnpgppH+c+AiCP4tJoH+8pKt6JwhY55fD0HTx1qCGcx8Y1KQQ0rVYp//+lnd81vDoAuRRdxF
5Y2Y3uKaRbnLX+DyZchAfDPDH0L2g68xIuYrro42x2RbD6UjSfsBylv+u1EQGHCSplt0DITKPN/E
70PPoiJjb5vJgalPrp/WE8Ep+EIKSFAi93LcnZA0qM1oORBmrZyaNg4xx/oYDgJbjTxn+xZnNZ3t
QWk8UT082xtPkd3Z96gnlBgk1kETE1GbGWgn6BBpUrfS344J+OGxqHImDr9pRxEUu3WkaDJFH61h
QI7v7Vz2PuRn7IUnUbdjSA2fnibDHK1PE1pgG+MH0hyaQsBTcnChHI3vny/mRnFFIVES25mtyr23
5nWcGy5G53LUYqR+r4/FyB4hOkJTJJVCQaLGudnUdG1lMjeUhySHkRA3j15IeRCas9GKdeTkXMVh
J3duJtXbXSx8mmag6RFkh3ewogrNmQUy4oDk7fZyqSm/Bd+cCpR2Ja0c+z78h+OsLWgxbd2m6Uf8
EIGCG3+lzd2XzhoW/v/N3gE2d/gu/ea9Dh5WNlOsbYZxAauQJGQXuT8FcGag/JvJA/yq+CyPi60q
5Kml6CFb6carQjq0VijK2CgcFz1UPEikzH/4Rp96tj6MO1dvVG0aLTVYcbI78p7BhS65rfcRPhuu
ZDUwrluXnIcZtyxeEEnA9mvlNRIOPyruLBfuza9mqJwl9+YSPvkyBXOLIqY6lOHz2fHcD1NLB9WX
TxcN3FsDCU13ZDDzCH/qo1RioBT4SnvvXMZ8oMLY7Te5H0oFtpP7SzRW1562582mRuh07KVPppXs
gLWRqWKxmzYDOjhkVDM4b8TQB+KG4dvBwseWgxgY21wLdUHh47FT8eijj28Rv3s5NyTcp3RX8qdV
M6TJGqY4teYSCM5QgA+fNf36klG1GZPK86/Qu0JGPG5XcrlglQmF3A4sGxSp9CbX/OWqZiL5b/5j
ppxeBF7RApYTn+qMPkIG56ZRhzFokdCC9w4V97He1Dokgr0APcIrJwCXbvN7VCVWlkuYaFvGFwMi
M5jNBGcLymkge0jFHF2sEpfx0QVdCtgfeJpwj54ovRCYFvL5f5kmpi2VFvamIp9/+VGCWjHx4IFR
MScsEiaQ1d+nC8gOMqrKTdpl7S5MKk+jvn3jHpfYdIXmnUQWPqj40yZOgL+aoL/wNJLAEk4snA6y
jTqXqMasvLXF//Wr+gWhkOYeYrqBPS8dg4vFJ2nnNqB3AowAXGYwXUXXWXoV3y9oygAJXAVDoePX
2NsQqByLMICM11uxEjTw0sz26pd6hwV6Sthp9BZltv9s12pPHnDDDQFFWLK/SibdGlbiPrgiqxMr
OEGYCJJDu5QVGr/EExqqI86vISa/jgweRy2QKrg0vhvVDPNnwaoKS7fn/GwY8phVBUTmp7Kev/Ub
YnmDvDMb2k7NZj5iRDm3FChCHLqielogu1Z37DmLKtxKQtB1Gbn0w+gq0v3m7ztyBjOg7UrEQyI5
S3CLhA1PtkUyvDNfU8Pq/4Y9pC2SBUi9bKbG8KM5WIVKrvfxQWVU5wdSJK9W9GoznMEbQxbK4obx
nG2pc4BgYfBOTEqMCRWepVxAAwBHe8tl6y3nyH6dsUwH5R9+z9pA2VL0KkBNRVd++T6963Invf/d
UYgWLdQRKWCldjKuhluGqSH3R19vbGe2rMCCGRohnvSD1LTtB8CNp1aEZ0yIqEYBqI+NfzPTMqUN
CHgE8a++l6b6u3EMdbX1t2BBv/JfEGH+9VCjuUgzbJYGa5dKl04dQPux861zdtbQU9ZHafyQQJca
cR4massgt5FOoI9iRkgZfIDpblhF2DvANzo1lhbv8fb39xr4lDOvnncW05QXUEU9VY6Pw9+ju5+3
0AG4rWI3QBqxN6z6y4Nn/LRZ0gKp0kBA3ypluUbiKxcm9CsNW45oWuFQP/U1rGwUqPyjrtFGMYpR
Bit711HNT7a92cEB90fWkmoVCbyWE68S3enmEXhHi75QSzNFrXwBXmss8Ju3pQheqL8kqRTxCVQX
J/IXFAZXOcAENuLW5ObgTs652lWDf744IKx0IkNfVsdwXeZWjbQcnNtvWs6yUCkZSbh7uIn5aUzS
v3XdOv/G/nOIJshHMzzscGQBiImRCkJwaOkjOx2SYEGBH+UgT8YdyV7szNqulwN5jUhQe3kmK7P7
FH8j7O1O7DlbWpYgEWGUVOKkdZWMyCKIp7dZ6JM3JQIYyjzpbVronx6MknMSoEwRuydbM07kUxIh
AZ5er/v2Jcx9OzcNCG9rRN8aaJnqWHsPLf2jI0lrKyZdbW1uWPr2CswWUXnhqjwIaKFkhb5k81UT
TJr8GQFn/s/FJhcr/6wePdCnQUZ4VI9pyyG3bLQN7R64Ghfy1SiOh1z7870TYEEUrgSg1fCGWo6h
hYWk5968ORnNUMXgLZIj57u/HKzJPDJH1DkW7j96CjvJbg/VhXmA5Q54gFIoy9ZpUCgOGj2iw+aT
zV5ViPvw2ng5rxIExS90WrHebE6BGs++XQVt6dFO7b/rjHed5C/lKPA3VvhPeXn0zIHevqLSoRo8
ggb90ZPySGwJbPJAr/q8B3tz3G3/1GiAsEgNry4xYbQuE7h1Cp7bgdnh8MZOYhSTIcJmWozrpl5z
OcGlatY9b9vbLf4CI02kiEnyNJH0QWKq2cIR55v48fTbpEhwZrUnR6nhCDThKZs7tFNByZ+Vv5sG
KBERh2jT60r4YGh6dDLatPKB6bOAlpYaUeymhQo69BJOPxNNiTh9awhzAuwATYXqrjkQ5cgESj5v
2aFgUAag4MQWBN5yG6WRm5rmG8fLIzr3Q5iLXONI5YgWjlmxNsMS5EJlP6aPGDH65Ch4O5yejk9A
brNI6BzzldATiVxnv+4A0x+/QhI5tpErmLxn8HKyVNyo5KBceEus32ksPTV21q1CP70l7TOB7Wuh
QEqfPAAejL7trKWGZAL7etTf7mox8uKuamirH2wjQwlRhyEkTDhPC+Q/47W7lnHMv1J5NGgT6Nfz
elarKVGuc/S7Mw9dXenXJNNsg3y5iX/A+fwbeda0aNKhobZR+N8JtEOLQXpyrKbmyv8ZQfV1d7KB
2rzDNtcmzmYJhHAisSIrqxy1YHvqu405ZJ2V8KoGh4bdK9UbP2nQyVwgkkb+gq6QvRlVWgbmn+GL
7qEDyxSQiaM3phsTl5mbQsmoBiPvxEP3JwGuuzWS4HzAA1UgIAMfRMe6ebVF+DhpJL32vtDO07XZ
BSy5vIE0HfJMT4SJ8fLbqO3SwOZbsPXXX5JiMIE69g3QpkYmAffywFHc+fwSCksjiQH8StrBDevS
1zwGu7CRLWIynZbJcwZnxTHQDFezw9fuPWYI+a99ZB+ikado5jrEGYKTIH3Q2DY4hPY6DH4tIf4X
V4Zt5VBE2+U4rMtX+8bDQqkqsjTJnbOce6wNAgKNv5GRSWSpWP98PDiHzVJUANAPiS6skOb0yVqo
XJKB0j3hhVVwYdD/VZjxBMX6qJZqitkmbqXXsh0vFA5OMHZIcnHUhmvX/F9i/57ENJbZOV50CCfN
l4y/B4t2MZ3Aj8QzXFsa5EUJ6HRU3Cwdbm0QOnmldYmOwyL9W1pKuBIVLmPJUUxTUYJVELog7L/M
E0geOBFQTcKIf77kTBwqubUs7QXfoAeARhiyEDTVHnWlfXTCD/uLHQd9mmwhSMHyi3GyaUXgFihx
KEF49Ivb6ZbGIH/mtAV7MTWaBHHlVVMes4O8Wgzqva+sN0irYte35OzL6Z/TaeBFb9Da9sj/Bh19
2k500CrpyShSLbrY6uDIdwv8HIiOz4EvZFlYL8D4g56E892bauXkWAmCObQ7C27wauYaA6sRUnQ+
/6GGN+MzOj16uWIi2kSkGoiVLIFn7fu+4xvmFqgEckz2rfkMw2u8XaBLNb6WmdUpGlsYYF1ro6EZ
xwFKdnXfMI4zy0lm0f+q0uvUEeFowzjOfEVHEbPAFcyvA8vA6sewH/AGONMh6e5tt8f6kuN4HmZY
eZfxsCdPTkLTZcJ6zZZF2o6Rb5Oq45UASyIo+kM8XuAvrDWLboXispUOmKVAmWj8x7/Jl5kPXMZQ
bTNSWUStdTzk7QiC2wyY7t/MOF+vl+Jh//sALpL9isjce4nhfV+6/81TlJJqU3eQzfgYwAQuOPbl
qE5nLSLO2FiIs5CZkM9yBBDYPhvCdV0fY0ePXiiP1vT952jHdhX184op5AYCc/IVEHyqYTqrhswM
RAhqXacX+tTneacGRhoJ0nG9f+D/iq+E2mg9IKCGell7T9qWXXNvAQJv6r13mGCHCnWVMn6hdeID
6WeJi4nDY81JmVJPmbyE8R6DArBC8GwiXXGHCm6hWUvqNmke42RkZPcVYHLNgBrcMShv51kshN3w
F1FNmV4YZrpPj7bxMYbO0TR8288jggeaVNgRZCPb8/hwlJcIFNbVvjoGX3pvSz8pbJTiZKeCNpm5
MeyEa/RsJe6bS9DpsIElh2r1xp8RdaQCl6pZjx0WJlZF+pOPmKJ0ZEKnSx7Rq6ZtEUXOYqPJkb1i
pl0fwK2CCrNl1m7qKpKUTZzwEgvAUxJ0WTxwLZLXJfl/N/xKxNnWbo0y4wQreefxCA5VA7lin1ti
gFaZvqqYeKpCYanZvzsmwmp/p/xuTY18J0ee9PfD2vWggbzBneH+VnaiB38oHcQX0iB+CQ/qTFSx
y7U9zf2eikuJlsOC0Hf3Y5P6b5Twfn/fOc+pgLcrz+101SaNQ+QrBkGAVEOWhM9GIit4F2fm/dxA
TuifN9oGaKt8Eaogj3Or1j9Q1EsU7E3yb4oqgIu68RSlyHAciGb8kAYBc/cabkdWheRKiyrTsw7b
16hN2PfYjU1rLLg5k9HkqIa5nTvkIcmT5rmhtBLZ/v4xGjz1GnmnJ/PcmokG1A4xPqB/S93YbUds
OkHKhNPzkTwUtG1vbEkjwC6onrWrABjZRnyDI5WOlzUTIcYN4hxSswl2zcLQo2sd64XMm8vkpWDr
3ehUpGT8AvBlqnjv56Y0p8P5WspvsGaTkbvXgT+Wu3rlAw7+uuOjcvVz6BVWpxIbWYwp5lEsRuhL
4BqlJ9vx6bbx6X9GGqdWxTGr+oVEb1F8TziIuCPOX6D37Ix9uCzhUdvLziXCmyPWSbTBVY7WN78U
xHVn25CYFmU73Wt/3qj0IkdL/8lFWfDkdX4zz+Zjhw5exkzhUE627aMJRJ/GAeVOKpdbk3nuAtxq
KPkX4GQfqMgqyuko3zpL5m+Io2D7D+U/u7irexJ/ks/CUx/VwwTogE8e97ZaBOeMpnsJVxnYvM3C
jQ8NLun022WTbvc8wb7ixHoGnZ+pMQTTuO8FL/R90OgBlqjv5XAJZwTgo4/JBoGRlB67n5hBreY6
1gmxjAIaWADWNPtaf9tdUV9o+RGCVhGTVl9Hk3Y+hXKBJj7Wh/yROZ0Q+oGnBnbD9f986TLLBHQo
nNmEQiJGbVVz6pqsjP/BRMzm5FtjypyPBgYtycWntDDiSrETN5ErTVeHBE4gTaRnTnZ/nKkThPh9
wKB14zHrEQib13n8bEBd03+NRb2a9FS0sKJvPEE6fKX13afDALlBnu6/eAfa0nO4MohC1mbpf+FX
iJ3baZ5+h5ORi1D3hgu/a0F7aVil8vCHS+uUmDV8R4cQM44fPcj1rSaBoufVDMAMvX/JOEa/TaH/
6FQ5MiBg3+b1jIzEUvqT4VNu5FoG1nIPlPGloFCA6vYhRVDI+p3TTSo81SuLg5hFeBWvZKgvhHop
LZPusuZP2dzBlrXMGeApu9slOqFWmdUWihyojIvOeFuMbhuncWZ60ysRqt5Az8ymL6rNA016tjKS
nd7mLxbuf+gYC/18T1hT/1fmIwj6NSqoeOJj6Ulb/3+VbGXWAp07INq819/gSRyr9udh16D7M0zS
B6mwhsy4bYa6tIhic2U9P5lFEuhUbqfT0PUN5z2X1bx+dnl/V/oObPYr1WkAqWtf+fFd2hMkQRU1
9/pWF4nTMZWorNhYdaNiLDd0q6I+R4QUHLu7v/mCP6XH0MI0ePcmzcoyVxqeaBTU571KEabUehRe
nXc6LjxaEGQCakYNzz6hcR4TTZ7VRd3QkVdSLPNY68YrVk8vHAjVLveLr2HYkCUR9vhvLoRIl/LU
T+ONqQHz9wa/exJdkjW/JPF0Aj8z8jBQY4/uWotuxa+ebP4K6g9/whDyYGEhK6ZxWckFPAR6O1Y9
289XcY7kmfkW17dLkI8OM9K3zqcFhOT88uKRtAyfqphYXWK39SQM2ovXy36+8tniY51Tbhb/OsSd
MX5yAWRmfb4EkIul9C0MdYDpEJXfctAws/3eCNAmDatSh0kDAabJ2txMMjMPSBs/syWl4FILvU9e
pkGPyuutiIeFxN4Ze2gfow4p0ZppPB+SKFyS0wPUBRKfHAATKYJwIZxbXC4dtpTBzOr7L2my/Gv6
/ifQ7UE3h/JlnurTpLOGTWiaWucy3oECCQ3gSZoPyRu2FAP1bx5kHRWeNexGXXBVODV1DH/oGCN3
8cYOhK8Ih4qBhChtZGt+lfu33siV3vB6OglwUWtTYvOvcbof/FkZTL1cA/p4WbiOatYXKH3meiZP
5UBdUm/RmNaL8pKXuM0fJqB6rFRym/swmOuTfi6rfePuH/rTOiHU8HIZU+AQ+K1SQ1UE8OGuONCG
AiyueSGJqR5Lt/JjMw9zMO6hXBXVY0etyf5Ims0J0Vk9WpkKKbV63C3E9w0JyX2GjRhQBRRpd8qW
lUJ6nSwQFRUL7GFzoeeQ45rTMQ5XD4dByvA9cJ0LqhqCClN4PMLk5Rl3EUcWis36cb1lHOSA3EED
/flGGQ8oFDSdxOaiXtbEA0YuUrDWaQz/XBV+DoKbV9Mt3ifFNuJ7363a3EQ3fFGT9ZHTVzmayM5e
VNQTOkmqtmCEbjL94L7OENxwXB7BVWBOd3TeMTJ76dUSDEL3q+TvtbIlGQ2sQQa3hLT+NE8cTCHG
pyP7UjK4kaDNlXD/AsgkMlfeH+XQconLi8gNVJEqhcPUa9uhaBvbi5rj9YzMNfxqYiedKHjl9bwO
YtkwC9ZvCkOmIacv9gqpFcqDfiWPGVyxoGNxzW/F8S05rEbHe0Qd4LFMHs3bKXXLefZHMsluIYie
SMP1hYJ54+An241lRU6Xfru6Om32EVkAtaMKd7jWWg96BfHO9IghP2vshYBSpeKYvDsK8Uakjf4A
2GWjXQiNa/Sf4gVHCw5uKxqfRkLdH3sQTk01dACytC/RbUYBKeYgPG/zT3qNneNJP6EE3oJx2Aw4
pO9fpOnJLQeun4RHEwHuENfdujnmyZt1MnmUi6OXW6iaZp1z0Yj4+onDH4i8+4gUQf+dn8N39kGD
B/Fpjdm7k5s5Tv4YDa8aUSpHOL+sm09GtkAboHtqfDiYsONi3JQax9nF9WZsr5vLytiKp9tt4SQ/
RzsYY8Smv6ZNV0xNgCHtSTG4OY4jq3hWJfAI6XRTc1zZwnc//747XFD0MswTPl+hr8P/Zy4FJqzp
g2w9d2g1D72Y2dc8W06rMzEDF3tFVmWJoBftKQLQdSzUITPYwqZF580vnZKzsZbisQWc/j0iZubJ
XqGLB1dF5zIbtJ4MV/cViYJ+bmqmVSySr/WwleTHGIe06SELhHvLn2IN3phmU6vWMtVvxviLcdcI
siBHLVzapBllQy8zYIggKZfpBVYjdwktO2MBruxQnLWGYHjH6MTs7Pn8yHyqD97blUMhGaJSsM8m
kWh76dJR2LDh5xsS4wDcRAnUsevBfGaTMOB0n11mRaUh9K+n9S1WBjLwc+AF6Ys+DeLW7sc7qDV2
xUGg2k16LuQbz+avEV2tTROUTyjTwkJj/vfGDpFqqJkS0sohr1EJVt78yHpHkA9FwWoWkj8cI5uk
P95oER9SIp2dYqlo1HvgB3lk2r/B1oJ+ULVtbTX9bUcfKJRiVqlS+OV98kWncY1DmjjCa9iMkRtU
3qyHoaY1wsPozSV5/rwlljIRPNX/uvwZu2yHwJcRmh7EdbKjDxJEobrO71PEHMdTUif9TKOThjIk
HtHOqqKE+kN2EkUYisEZnEg4t/vmc26sO1YoA/H+G0srOmN7JLxWZgJH2LDN0gOic5/fENuqvvbl
GH/GQzjVklmblPkiA5EYfRBdE7CT0vSz5y69xd8XCiI65xMEKlFsLrQqBeFbr7hhBLS8PyqPO3DC
yH2I6FeHExXGSc8uSawNiYl61b9sPVNzlysMUsjjRsdGP7YnAYmMedtbwrcUq2Pbg49/6auPGfut
R0UrkdXIdXRqJgxhXG1LDXxSXufeeXAQLj75ifXy3CMy8XGtAPCHlS8/TQZ8Qb5mslVX0BtItMkd
oSEaftvUBHHkKpsTNpwwlJFQ8q0SiSbbiWpTy31kMNFPep9HYnZbdDTPS5mTVgqSMIuFn6ABx5cx
jC4ZY8P7nbDFFIhq46R3SqjwtEr4DkIiHEWSZf7328hdNkMq4FudbyAyotuX3YqUkJYdsam9KWuU
lTwLX1VHnv5ELR4kbq02hVbIH4elmWVkE9BudL5oRFUGUY0voTmiUo0PLLZ79OXGe1EMe2krx7/b
TRUZUKeWqnoOnjtH/19bLf4i1fKjdElO+SqnHrxqrWLL8NcmHnhIfU2IuyRkaoWk3Eq37Y86pR9N
FhhXg+KCArpqr4a+bt7jubpPdva4iqpe/6A8PQEc934wLSTOpixeazlgs9R0Vc4fuVhDGjyJefWp
GHxgZzEBDTKc1MMDSFA/uPbOtO13gufMZHrtFTv2jJuvpK6Xic9wyTvpH3PxgWxB2tZv6UVdp4Hh
b1Wk0WNtWxoVbv38t8pZIxJ5HHv40a1QQ7OEAQjTfjONq2lz83Cr6XJKWYssLaLAQZBxfO0CP0th
hWiocG70LybjWvOnWRUE0t37IFROo6jSkbVIdzfERBRLaGK3DRkbF6k1Q9lG6aP+PeM6VMdeC5J4
l5MPspC3hxSv9whOa7kjXZIpIFrRWsVsoxQGueAjPsBv5pmOxbVkaG5cce1z8KGvaeOGjF744rJ9
PcO9WmReeV7yBuGSRBpFhLQSsSXQAuwyIk918PoyWm/zatQL3oBfc5QjWqm5GayNGNQDMSwlZ1DW
uOxaVzZE6rHitDV7TzluELbtLxGN06LbN8XOT8sYeFJ3oYAvQUfAkEsN1bfHU00uHBql8xeIw/g0
+kQ5eHLcRy3pkf1KMMaB2/MRVb2CKZYdGgmsf6iYc3d3WtegYAFyjr2EFgurSXdTIp0wUw+DZ5lM
3H4hABEfCnSITNZQ79qwEizZhwiaH7Ww4sEQcCG3YW0Lzp06wnKd+M0GQtrR0MHPPXNhmQ7ylBY9
29s3bSOiBMF6+t+pllWDpJrf0M0TQ2hsIgSixA0yi5e8YZfVrW6MudN24w1VY4dWdUlx55QQArQ3
TODCxmL2/Cf6WJ5pQ6YgAhZ5m60pz/03ZsI+vQDlU+tb61meoV1syHvR4YiKJ6WyMlf+u2EdCjJ3
jVdZUcTAtyavixMCQub+cXf0paDO/tFA/jRpJIE6wxmgfx1JQXlOU+O0iSSx1am6Vj4aA+XSbJQk
YfPXl3bHgwgCsUHWFNNBIf5LGLPW/xO3lHJA1/tX2Tch8GkUCOPPVzoX6OWo1z7GcHOM8gKHtDPz
KS3UnuG0wbjHMLAqsA6lnpKzYkI019f+oLH/okHEXqW70bqh99bWhbKXNnOEbIX7gHdCOqP2AYtw
I+TYT2U6bZiG1yvWdtk8Qou0YrMajMh7ZkI6+yMGUIII6WPpqWIRB8Yp6KxqXE/ugJtlWhr1x47h
1hi0KuKyABuymUhSMDBb6kjI2/G7X4DbCvkbCdSskAjgOhI62zpb0WaH6A8xyseWlV+jgZeJeERU
+RD1at5mgOlv/Fby562xviJe4JEKrVLFLV6rNQxTtSZfoxON5iSQ1jg1+AXRpvJnnW8IZahoLcCS
YXXkjg6zZf1ZsofjAJ8zhFh+dX+1YVQZjeDIrahepoErb0dVeIw7uyQDbY5kGSZ0GcAVGySNz8CJ
usxofMNbgvuzcd+g8cHs2OnIvth8PNRNJ+561f1n+oSpnfsZx/Z+lQ0niWr7i0EYjySs1NsxibeQ
EMQtQtIwm5oD1jRZ8eFWO6yMf+R8rytQbiad6R55qGwnpVnxvOdnSbFnK5vGOCwQ9eU4724I+O7l
kAAhSmCiFzcMPQP9wVrSnH+gaOradyL56bktfpeoe8cXPT5YeZoZfxB5IkmxkUz9m4WdioNLbejd
6CDnNT7Vf8Eo+UhEbZsKhCnTPH61eUssmEnz0yd5zIB2JtC0GpFa+j1NuMb4YTUDjjlJiieZACZw
VS60gCJCFcwp0ua7Oc5hmu5GIp7iFfvEc81rPMHJy2VrmAfUhqkpxgeD0ozqv/YcCDDnjLIjef3b
hflwpL7X3jwKP5IIRR7jGvVh8Ow1ibuGBWhTUB1mzVm5Rg94RvA+v4f7ehDmWxhetY+2XJP7r1v7
5gCbiv9jVH/xlsmBhBWMFuvox/setl3Xr+Ssp8qLrdkQjMDM1iSWwcTaAdomFYMkaYCC8i4X138a
w5XauoVAjlFT10VjthWGCGtI05Jg6awyHtLCfncgdP4RY3lgsG9+nXAYIqMbV6earwLKd/wXikxg
Hr1N0ap6mK27WWnuW6GKcalZ7Z3pz3pZ3pp0c0+jXXFDFtn47AdOv3by88v/Afb5mBDTrpb0YYR7
Hr7h1E4HV4eRuwv0+k54a8HAKzSk2vz6qbyv9fTcBwJncj1LqUm6cHFK2UbevQSDiTBMDugmetIy
oYTg8g9BAK1+UbfJUaNzCoGISGC2TeSiXlAVBuw2KL9H3nRgbicF3vtqzuzQZWKS9dPJNNmIaMDP
DTxM/yVMxqWVOcqwYsUk454GZob33uimh+0+ANLfqR5JrCNSfTs6C87V1KaJVCeHxelNlEI8a8zU
I4fzSc7/5EIrH9gBNpcut1aiQdCD2DMDBjN8wEFWj5yHniOvC4azWb8zt0XNvMFJ1+26cw4KH4Oy
cK+9nmd0Hwa9LL2xhUaObDJlIcLrVVH3P6ZLCV94uDxaijPVlVSqtRSEvaRoa3fDLuunrWrWzQbU
4vIWnpcGH/FK+679L2bIP8jUNdw1wu8pl2rhwFAyp21krwa30q7DQxZ0UlGK6A/+vo08THRpPt2T
XQ/EOjbmI/dxBP3oCTrAo38GdixgxKp/xD+SoGsqZ+HZZyDctx5izzEXAm9fhbTfGHECyOQr5aUK
IN/zL10P7sNr+D1fgTLbd7LCiiBZIGISxVdabgeMuD+glTd9QmFb3P30otGpYb8jvh9ZMj4yk7el
m2Bl3hL11ALXFWaoMI3z5czo3d5sSJGzwSAUrIz4WleZKKwUyQwU2SGFnxBZJlA3rFJVrcqTFZK8
t1c5fgGKFuHCDlcleQZlFtO4saoqUa1DsTTdmfxbwhr8rJS+tgSEohvMGckDgaIqaWz4T6jzB0gD
uKNqOnkcJIvmP5QIIBf6YSVTAakociJ2Xgc9ZY6T8yJKP8OliNBjAkENs28LcuHzrvi5pjlWTL74
dPo6VMDL6RSJH2o9QLgZIgXBEHCecRopiBdrkIOOK6g27buBsLvJp/NK/cKD3VrbR+JkEFPtgwPQ
1Rx6cgncXJSizHBvtVlw05AK3B/YuW2ls1Ew8KyrfgAljElnxVr1xN7K3rRlbtBG7SJqQwHV5Zp5
oV29U89w64aSrVCyyMaxmpwt4qwEE3BK26SjPPeLpWtRfn6Cfe5cd+jbajgg1zi2bfqvNrvVEoBk
NmkrZz8p8fbs9IGRcKzCNS402yGEbAji6LuaSTdbayekbo0Ww63nj85oIGziQB3fwrhxhkLw6Fpn
D0YA0Rck0mbN58ILgcQZzL/M9Qldl0QhPeByHtszW8WA3Yalhmq2g5oj+o/PDO/155rn6I47uQ8G
5b86G74jI45wWQIDz2VYMoGCoRn9kgrwogto9vJLPtRDjm40oHbvWquzcXnFoqii0TlLqubRA9Q8
5whZCVAeEVxwuj19qLGJnXOYZpI/a9S+PHfMfIbt+874eNbcpIfKsNmSVZHW6En3XivZJUuq1MaH
5nHpRX8z/g+p+JA3+sbnGkJYnp5F5aqU76kl/u6kPQcnzTCYzVGEf875e49TKFZMyMuXEQNtcJpY
4KrImiXtbMUQiu1sLtxQ+tWt0XW7Iny6PpSbfhmOVAq25lAvZs/X8QkqkbINqnMYZBEslLY+zM0g
u13Uf0lrptbl+lSVbBRrkPuCWQft+9gaKNODg3FtoAk2cM+eTxjgWoYpWGiC9QlZ2jT/ZsaU0wVg
LejhdCQE1DgAXz4ezJnbzpYw/kPGOvFp7onnsknWUHwssQNEbjUWmavZ2UMB/ow2vnusGSA3VI6C
mwrvDOseubyIFxtuItL+K0i5hrQLldpDhC9jYVwBMes2K28yfYMWtwHPmCNq9XHLlluaMfh8/op8
bEdoz4mKKQP4Tc9dVowLhKQndkTDxWVd6uCkLMRHwNeAYCtoPaIRXemi0nYOz1J2bIZl2QJ3vAhq
GCkmtkJFNGm4M7US8ww/G8GP73lylvyFOi3N7StSqp9/vCXDMxtLbEPMl/C0FLNh77JS/oRNqdgk
8ShOB3RuZ8mDISTlGTDSC178fTF87ikTrIHPzwn/TJgbrOzejxA099DI5NU1Sy70yDTi6DJR5K4a
t+8uR9Uo90yAXuhNUPtab7ozfArMZwu6OBJ46A5OXZdoamXbiDPnEDT8jNowL8c+x3mjpajWTjQk
S7PktfQf9XIoGMRMgU+8BmxxYBA/i/smB2YnkoTrlv5iDpj1wpoCg1b6UALS99yAc83s0u3zjx8h
D8K+zabQ63GwSUH5eUp3mEuN3NbnE8QruDExtiBDzH2vYT2jfl6zegFkJ8XlqncqCKqGGrzR69fs
YoGiMPpmv/WzYMqkuIF6ACegANCYVFmzlTAEBE8O7l6AEnOSfiWaXs0YIAxUVbXQWn3PXlPolNHv
bcoQy8sn4app1u1DqSsZIqgId9+vpz0j43bhArYkYzQjFIL5YrAS86935Ce0knAgh/At955uc500
KGo+cCyNKJfD6mCAfTqtIX5wPjr+oqhrTthPv9Pr3tuX/VPYEbvpjwqTvMoVE6yXPwstes29kCVB
6hDqxFx0Wb0z4B3WbWYJVpTMhZasIqesHCKjVuN6UiPzwujoieDMQyDqhXmv5rrBZrZOfahNOjzD
3fcJ/StkYn6R0enKF6eajKQMFvT2LMcq4zpcankXeFm5mynHoQOfZl0MfzyZz0CKLXEQZPHDC3xy
SqW7yFMspd0U7teZekoEneLHXITlwYuJA2tFO3IV3A6nUpOQaFF/8FWHF4OOJL0qiGdr9EMrgTuB
/aGDT4QE62W+K7JWKWcI7OQL44Y6MjEMx3U1YKaGk2MZtCdxKNzLACyq2GO/xrPCOvGe9odN68KQ
V07wIqxfp6F7Q4D/J8ncItK+alPsSq5uYAUBVY3NCApLTyHosml5hT2K1u4FsI26JHCtwkWnkPhZ
Vyb28aDGJBEgiiA7pOqv/lrfOW0tunTKwF1XKA/3mJVJy7HasqQJ4Pdnd4lCHN37ZZtoFMBcRuAU
x+uTmbwBc2zf1Ga6gVBCcDG7yGotwTMtnqpUezV+QS/Ngb/NcOsWrDYHC2o7kS81UpIprEs2LZZN
XBjBFZpi2MfUBMlemP68JFOWNCM/JtVI71QHiarDiHr5xalxk8Yx3b7jB1jo3Mx1CgYaq89t9nmh
hV5iPwfKTwl/aFlLcSelLWIj0McqyaFV5NGUJWc37SZtelYQUiqnm99f0fntJKqVvqXogC+mbfLH
tIVHEz7+8agBL/hiH0qw+cQqkThI1/F5YguChFWaWWwS35GHB9w+od7cZqO61B+vD4+Ptgun0yYC
7kLFz6/d0DOgwd5UPlpr1hfzbueSRrGDjEvMLF4cM/lFrtBc/iQsztyB6J1lqWGHEJ6PtngAIYMm
R5zhOiZPO9KW0t5so0l+GgnGE9XAVIOEzDTzjzdwnH8cL1e8eXSw76HPwPIlpwml2AU7cIqQBWHN
oV+krOz9o6s3FSDeDPaC+WVQQ05cTbE4QbFlUPjFh+TLVXeTUeb1cGg/bu6YRD6CkY1PKhNLG0vy
VCJVf+xwhDW0n7HR5Ynhjexb6UZz6O5BSKItXn6xwRsBachu3eSux7t+VhnADnT10ZhHzsNtRgiT
gQxq0kmgt69qcRhkT/4E5X30QCI9Zqz0P0ZFm4OR0jm9+d2mtUiZBIlHPasY6pwpCl/m8kXmuYmv
io7PVceJaR+VeJOZA/aF5Wx/hNXNK9gPfvW4Jelx0VB8voVUiVmx4UJR+0IxOJ6h88HRljAMY7Ms
xl0WenwG/qWgauVeEKo0LfEduFS/s9Eifl0yWEuqVBHg1ebynXD9Cptm901msHnxtqcU5rlYtcFF
4ow6a24Z2kFBO+nhQItkjI0VOVJfv+6yOtU1gNtCxEaB6DXXthaxLqm9IfOf5AVGkgQjeWSG4gHg
5H1qm56Wup+0heGFcnt1fr5A8lc22mxwMC+UsmAvM8CnQb6s27WPK4NQsZTgr8SuZ7v00E0dNbiy
23WHK4fBG4olbqLswwkyl8hjJcTwWRM7zWIzeiQCemKcev+9arQkOVJVyw1XqzTLiH4fI04SBTxn
5KE/VTpXjpPFwuxc5M4qEtXAr04Ihah3wglhNSicH/7PZ7Wz3Vp4WPA7vx5HjgkFrB62xsrsxOBi
dGXc6zlYUUKhySBwlsXmpv+LeQptsnOVlFdfFCiUtEy8TyzxsGuqz9V04eF+SrwH6oIFHKNZl2/p
1lQ9N5bDkJByQ98E4tQS11QFgbPk6nXh7yuQPWeY8YZOa8fOcbSwLYz6suzcB5W6xBpWzcqEnXdN
dlvtvlnHaJPmYX+/d78pu4YQGtohbRjmSSd2pd7i6CbB+R1d8XwHyptwAsuLp8yP4ax0x3od5EUm
7J6yXItbojT9lvulreUAAkPAln5P7SDduQG3/OLL/L2p3/hi0w4u7Y2jak3wSUcX5TFPjHUT7Znk
vMXa2RlEmK3JJJuO6wgnLDjttd4exFX7E+08wN+lnz/B+W5+7ZbTBr3z0Y/DaolFJwl1oBpK6GpZ
iPhC9NhDH41vXCrA+0S3WVK+0EFzG8ZcGz2X329qpvcoFQnfZIeqfNckjiwHayIj7xz96XGXwGZh
t0uSnPSOrW+eeSC1pK4uZg5tHL2fgO9Q9yQWQr5TgdvRH1JgAWxdhIYdUStGTce7GC0XG6VcMnN7
aTWD3fAnjOZqdApTM2PgS6eJ3H/kDtNxZQ02bq/vuQYKNEtcobgADw5svIcT4skCWO4BvhjW385R
MyaJBafak7Pma00eLMxkgYo0qAzv14aHIa4Wga6tCl2z/sEGxk10CdGSCf9xCIYFGpmd3rzQP4i3
4UqfN+L0+YetxRwdUV/Gy2TIOZzhFzRAOKoCGkZT12ofxvR2SCaiYFBf+AFD4jdPyAGAqgSXNgTw
SOssbtRpEIsIik596345Ik114ylnzi9Gmw4BxJmLusrGd9Rj+V23HoUMMQxi8fPWtF8khWj80iu1
PJATXIoHsZNT0SWmy9yhxQfvqDLu3+VqdqQeK05lhuVHHCOpKcEDR6+OkX+/soohSXhKISlY0OYe
J74XDmcH0CwYNOmRZmJwNWRhgT0DUbm2XRE/2iXuqG7qIMvCI8dHNwgkD/nyOI4duOl8sfFlxmDw
E+ztgbq7CO/Yp96JIPOJfhoU0aKHCkhLJzq+T8rm39PLHHmFUotpDzjXkiEobChNPVOpMo/9NSN8
SjmOPTppb6SnDFFZ77Z3Z63MbvfKXGzPq2YbqS3DczlBptXNSWOXote+YTXCwWdxtPMH5x7KNfbm
A97EO1AJu1GFLVSGcSxnOQ1/B1yBLvZX6O9MbY3indVriNlgKDki05AYpghw0imdwX2/oXQri711
zGeFKSdhH3q3MKp6XZy1WkCfLEBT6wLzymd8MFidMt+S3DD4fkBKVYx1ToCoMj9KOTDzhb0MkmAs
VcCd/+2p8DFijBzC1+H9i5+DegWIqvMEs8RYCN+wVl4TzlUXOrD9NdqycHiZ2W0e3hm1AX6ZZn9A
We4doYeZMMsNw1Geuh46+4EANgjQgcFYE+7rDX+LAj27ehHOaTOCRo6/AOE0EZ0aoZUj2UJ09OIh
aYW9hhKUXssAx5O+3DJU91gkd2Ad7S70cdjCfuuc9QTSrB2JZbsvYJxz5c8DvJOpDTVmbhJpz+qY
LR0oDIfjGNnGoKs3MhFQ1UOUWx1SGL8zMvAgyVT5vRWgraVy4NOltL7vjnfzPSkEhVwp/P6oPoRQ
jfEODN1fepcZG5IyjaeVVhaTkB7md61A4seY9y/OKEP524CVQKr6ZY8DSGCiAJ3/6ovti1YticIl
plLT+6S++J/s40Ywvyvv9vv6hfuH+QPDimPgif5Vb4AiDYjP3u58lwtPCoTbmdBwmYMwQpsvsQwL
wXYy23aeKtJ//Lm5DtO1S8jtojO6Pci6VsgBl/iUcCHnnWX83o/VvmnjbseHy6KFDGHblmZjgj8G
27W7UnipECb0Z4LWYp1/u83L7yaqhlpwGan/NM66gRWBuokoqd0n6ZUhBHiKrynb6OUBVxFpmMj/
xRv462TLpyV5VOeuDexcy6jRkCpXve6skr/RQkhcmwzb14MAII0Px4VXwG2PqYwIYwB3G7f0BJIS
xa5UapqpFfTNxEzqsMyRAfp7Lt190ws3AazXTexQEMHzwqIlbbPXREfxqzWzjHLq22PuBwqEHncT
40iSgAyCzjf50ysQRDFK9UhfRKbWDYD4fZTqlL82KTZH4aTYOIcyqriGNL/hq+2g8yNxDiVcz4lD
U1UCB7cMNYdlsAYD3+ZugYYnXgJkolvtdB3rkrUDhz+CODq4IPaF7qMZKvw8gTXnqKmzDy6Jse3B
YuCgCkMk/tIpHxMFx3igEFB8dxosEZTJvmfZz+LCErqIr/QBiDR6+E38TJdLLLN2BDC2aM911RLa
5EPSPsrPIGLX09XaGppWopWecKtnd072B9Tqe0tyn3KwtlajoHg2GjDZDxv44cJ6KrhzH4C5AqGU
0yh9ECnqdmVvUw+A8LJRJ/bu3h149R/xTN1p0tC3XsQu14Ok4IzaDAv9DXrcJCXeR/2nl5smz/5q
04XlZhMJ3zutpP9mKPyAZu8wws931tdTnBAS0+43GDuSJ/7KL6PZ2wNHv06jgbGcxcPr99v+FwNM
fDq96ElsQVNkWHunmd8aFEcUoZFyARgvfSN5sAiD+69/udBx6P6NiKZu7UCTRcmDHQVsMUWfQdx5
jKMwZ49TW5Z8Szevy5QheE2TO65auhQ/34orByeIf8JnswEbJ4nnc+ZAtJuq8nJbvJudVDFPBQ3g
pwXge+qhJH7VfJMXZQamTcjeQWL3fI+Ng6Jk6NVGPdc8mdzORIj3NNXlVBw3xvYs3qqQHHtXra8g
pJBbSANpfN/pqWpX21Y8xQ8OvJVzHxLhWdaw0AX6Mnn0CvYs49k550Ua7GHZa4skPWvYLQrsXEbf
dS43iihMrRdi4qKCXskfTD/YbWO7OJJo2Uen2KspIMQVP9G5ReMTGBo3B+lE8i95h496vNtpI7lM
5MDWcdKz+ii9jvDhNVsVgspZJ033bRwW++BcShCowcocmzrIKW5VAWJ+2Xv10CQ8lmpRBxAT1sLX
joO59uyZk6PsqcKEAyo+Zd7LnE5qWjVCbdT6b52kJ+V0Wk/KUObQjjScQwgSItX3dJyr9BQCyjwA
xGNPnuRSReMW5BhRJJI/qxZnvcFeR9d93jKEeH2AUAoR/bFHbG8WRQNAFE2dAH0hVNox0UFikj9P
DIECzy/g0a2MFWR/I9TCGnul72TJYx0JTBNUUSPjsnSO/qn0JzrMkbY9EVQbYG4o8kLkqqiVnFSV
pi+RpbwEe7AIZo4779JuflDdgdsS9PjjaBV96hP42dlbzwNfmzz8fgDW/B9OwMPdby2o0EUpFgZ6
PTP/zEC8hkg93ZSue8uHlY1JRC8nVdDEe1KftnNN2BhE5tQ+CwzQp8O87EyIYGqE4nfw5VAfOgnY
Gc7fKXLNS2UL2I0sEPmVpiLSB+nKX+GVCA1dDXhI1IBdpwJQWY1mnrM8JMXn4Lhcz5ky0vMrakdy
cSQ04izgrkY099bNaTSGgoc3o6tDwBV/vHnJ+5nEPOVUKMQ8WqSbN2t0y99Y2CDnjGUxt0sZhsTj
i5El+6mVP6yLA1HYG4mo5pDnY8rLjowRbTtys4jr9KRem7IFtjPCKHfqHcJRmpT/aD+iuTG80rsi
mtFDBhDScyo1BovjE5K8c6WD2nfxHKa5Hzw9cAZQuBhfFouYDjn8c+6aOmiV76J+OYMy8y4lHXVF
58Ntz5bX/H4/L4rAnkZBBwkOxTmQ9nvp4DhSpV2H8g6LUgt1V7Lss40PnZUrU+wCqWylK5FZyqR2
f5LBd+MqH5zVVFggqvymUA7ZwlnlC+CghxeF1+/0+xrl57wV0Gsyo4i2mYC94Xcv6+tVTYHmIXF+
B6rDa0CVwIF6w+QMVzIraVzLQVOG2u7BKlbnxRvn/cSa6nr2R29ITbp92x/p/eOJ/ept544S5MCd
pNvqjUMGx4K+3rbKby/cHI2kCcQ2HXWYWuRAMpxz/OqTLBTprCvgvXKi5vFMDjK7OwsySk6eAiZh
tg66YCYaxA4T/0uw2bfBPXkxWEOTcXUO4BtdnjS/ZRmoU+3vjRxr0RTDRAHr9BLFqVvIUqzFiSvn
+w/vDKHFbJj5wH0LDlwqO9fki17x0jnlcaGAtMga1cqlzKELtBj2ImbiydT9hyeuxgb+dQ9r8zuS
ZrFzqAC8Wx2jBcQE2hW+AJw5wq6yjW7bWaLF28x+/0k/nFIiKcHzUOvMuVPmI0Og9jGWsdSnaue4
5cTHmOPNmIeB3Kx70BWHyyN/61xa4fiAFRkOb8/FKXKnP40soPeTwXh4yFBBGxeMCoFCvD0rC087
Kd0tXYrKCS7N61u13HPId4RSkPxuEEejTB6G5qaOa3vvEtNFL+SNdpOPKASluFWr2x/qV3XKjdAe
LK1p7FZqrHO7vwXHXBgsalDAvNhdZk0iXWVw9Rd7x527QAbgjNXRj91LkXkoQu2kih4YDqHQlZCE
vmIXfhHp6QUhH0/LJXno0b9+J/3kfkpizROUnw0zMMI0rsAViXyBlJZScfZda2PaoprmWe9vAK4l
QqRXSOiLrKef/cziu4tTeinMRQZ6kooWgJwusCEaGSGVVbcQPlDiBZQ390B1FIF4iU/DGSVNfMrX
Lq9ldo+MM9tJFPvPKulFQ3E1FPJpaWJINUSlSrF5dVA92dKxkho8lSQLOSL0ceTHvy2zteyb+lHn
Io25cQar3I16ds4Rpxz4GgtHNdtJCwjv46KVp9My0vQLqIG07Xka+h2zyVUP+4I7zTgytKzEnMQA
/5RcxaY4+9egxKnEPnKkP2dy/pG9P/xwCT/N6clljEnjhipxBMPwKWndJ1cucZ8wj+J9A6Sh6RBO
dOguzD4f97RDtLLlo+23iFyNPwZMioQtvjp03C6EZJIx+lgjTsFzBq+5GRQVVtZev/dSi7BdcMfA
A6p57lWWVMB6T4Hm27fIV7ugfmG6GiC40UwC6091vYzyWKUhyN5fV1TntLWl+akrndkA3aVqMXTR
2eTNu7J2O6lgRS5XsfP6CtuIFgfdvNvv4Ex0ezMxyF49CuLGxPJOd9Ri234b3GLsvHw1Q+it4OTW
U4A+bYC8Aw6sLmVEhB9aOcMhhlleR+slPdi3bQI20fZIRIqsogbnrYfodc6GP0/b4dNcsA2GEI8n
wcJHKYAuE9A7+oTtxt714bw3+17E7q6bikuCSop314hev2DRRGhWeVSIDw5DSgPN/BIzrroCxXpg
iJkhHt0MbjuYyk7M24ll/YHNRrPYUmIakRumuvL6m8mrZjsWNzA0WJAWdlc/sRQikD4YJ2KcjoRP
N+Jc6CeJPCKLPbyGmW+GSzm6XRFiYHXC67AMd/j/h0jBzdZejCzkO6fGsK7pRyqDSAEHTBLGL3tG
2sQQwFHE56XjXMPnbfRgiYxHlUjpLZvCVPISSuhWbafgThbQHSQXJRfqezKkzCkrGbh3clZM+ERw
irDxVkG0zsOuLDX2joQPC6lUGu+/Nhskgvom1A/LlfbpALlHZ7zJQQHWjwJOs2lOKdQQkxaZI9qa
PPS+eeX+Ngmpbamz3pAAhTwjnmB39CDfVzGuevHUCHAaZIRZ8KAWjtnLGEr4XxydU2fg+iXPhVTN
tz1+ZYA0E0assqEvn7IuqufhA3EgNjdsk3RbHOb/OqNJPYV95w4ADQZ4COhkOmq4EczertD/LtCj
F7o1E4/Op9T+ANi3T46/F0ACo4uEHAjRgxMfhRfThjiNGWq0XDgLmG0ZJCKfpVHOt9euAk3vDpRc
SJR/GJbTwysa1lLZ7yfKn3KslpRD+okQTVXN6cxmQcwURdA77/XQHTrP8F20uj4EEHWMrJoqVGo5
bloTW64J+dkoz2E1R8f7OTAlOByYA16Z2Frnxi6WIo3gF7N2q47m4pO1aYnsJChYvNxZAU9xB48u
LmPCjJDmEnuB0uLH14bwWa1c69KiGnkNtFLN6CK95TpRYUpBnFW42v0hfrU8lGnDIQ+FPc1nJGNx
FenYARfNi29mCl6EVfHJQQHGJXciEf106kJWX0eRWRNkqkQnFAdYwbNnn0LHDyFPg6JmM3555lgH
2Rk9tTw8/qH7t5hsnsosGpSHy1KXMuvyriww8dT74I6/CLDH8Z+kSSvhC5kFWRpGAAcsLqjh+bvW
D4eF2rcqmW3xlPNuHeRVtgUNzw64ICD1I+o3JEpJ4voXq46QjRjsryVuegZv7UQq8V3RRA0BwIKo
urUe3MXtf3BnlvxRuS7Q5BsVbD0Q/7+UI5UTyw6KvUBOptXEgv6emlFikyNuBHh7+1GMuxzNEGkN
lslplnGMwU9Rmf9AjosRZSZT9DbsnB1Nq/1gfd9BxNdi6k+yzqV4s+IEWYjC/XW/ldPp9hmS/Eka
DGj+vJCZJFAuiQtvecRmYaKMqqmn067rkfn0CEh5SuvsEmXaDk940mQx2uYCBti7TaJ7YbIHAnYP
Pfeld2CCj51cDnTSP9P5fGDly57BIA0EtnWTfrmUOduC5TJrLtWW0mYEhcKxGpL3Gswh5pxhNMEZ
oD9aZbChpSs359cWvkRaDNb29H+DtEQzfqEwZ+O2Cxk1UbKfD9A/l8m/GF7DxgfWpH0tPDmWMB9N
AGbkHHxp0pP1J3H9LYU1jIJsQrhkPuBq0FxR1OXYOjMtOtIqikvmclP1GfXud4nte2UqRqXuKEBy
N1s9V6fUAYoGrqSfUSMs0v0Pver/CqWoc7tnGR2qcsWLmaE0ajQzCK/YDoo4TL2xONKBKs31X68A
qFgKNgh6t+ycMKnfXOsHpG+Ax8C2uR9eIxUw+UlP0HCxxYxDMzbFrkICYpPykhJlnIqgHNOLzhwY
ujNI9rbcVSHk4j0dzBm0Bo2nSHtwMQHqfPAOAoEIzA3bpFJbNFVZVIgFMD2eMz0iEphm1l04vwqz
W2EnY4HerMFHULh1NXpoYHiWjgyo24kEktNIp/E17qb9svgtZ47+aDjNU9AuPY7+5pd1bilSW6RO
8JgkDkm9fSCdMC6Nq5ViPFx0m+m1Sk3V2PJl3QJyNFJawaqRZxl1h/T/T/B95Hzt/RkDO/3cDJKg
9EO/uAs5a46w0yWWpQd10hNR4RBh6BDqlp2fBURXK3mCiFXrRts0ocLVFtgSPy905z34sEIoBUl3
YXfRoauftoLAp4j1ICHeb6KspPw+8b33x6n769g7yfrCVrreKSkgf3a3kwrYmDikELva/OVN7FGt
FBxCenTYU4lijPVKGnOhdAI728vOxvyzDlcrxyCx+zn/HYzxRkrloZj+dSkm/f2Rcqx4FwI++4qW
DieUUkZGY1DyIJpxYP5ISyqf9lEE8FVajcMyKlcd9BuIvY4vh4+2oQJTW62O6mw6Nh/ycEf8sbDA
ienRDBhaTdFrEmeOkbPexjJ6gPrMdU4R1/WRf6o5Sq59++BgLCpL2AMkYtrjOFhRf4/8DNK3ou0e
FTBG2h9usbGYaCELEIFVJzzEmQbSzVskTFe57goNyuhOqPMh+PRGF68GucXpgc8jgTVz67XrtZ8p
P3PlkxMDXpomOgjhua9ND+IXpGwfSItYJ4q3MBvm35I0g6AYGNxryJP5E1gx+fAOZxFeyad1VTZk
SMwmx3qdgv8AWA3+CqaKmwnpt6BEt4/ht5+kO638JhJ4w0rW/ZWwPPk6oecMbIlRSy/MHSnbY3rw
EAA6E5o+VjPVkJpqaMGJveb4K9P6udHgZPcVgz9Zllk0KJF6mTlohukxTYHRYQsV2I/EVwIvByJy
LKaAyIaBUZ3MmIzqWXkY+mTK4sUa/yNsoZ71V+NdM4t/SquCfunwQeY62aXTur5ibjCTwZAD3/MX
krkFzDoQOenKkwBG3f8J0pxz8Rz0iY0AHqxX1xan6H5p+dv1Ee0gLkOsv8TwcD6EhVseLXei69LI
mYdXYZc6ChkcvcooilRQL8/jmimUeSLICf6JsLZN79VOM8W0CIIVbyucW/TXtncEv9QJb0hAX3nx
ZFBUUZwFr/Vo12tymehDjcBuOCQH8XvejePCBxGSLhNMAO00AyGSvEfDUTm5YUj9YtfkKf/LUFr0
LFsl2SJZCaiUYvar5L/Z3xzHIQ/sycaUMnNIcKDuO4SPzGI4CGlCSPXA2KWuIEsglhuMT0SdEV60
I3vEpy0hFBgixawFv0aVMlVBLwUe+RM03p5d6tnG9Wes5b+xDTa27CDJ4iBIBxycuM/WivW2Z61m
lmOzcseIcHToAfphHB79iBDjQ8YuSO9clxhspOKgHyD49SWVFhqFEDWhnKeM8U/PI0ytswzSEag8
51pIn6McSOZ7hdJfmUpYNbrhnHSo3pH1w81mfMSI3vw29mhJ0K2eKk16s+c6GHegoIqZ98J6omIW
xn+5FnmU5F4AcKVcihjZ9VjHinO3+gEmvNUusCtsi6b3FD+B5dNyZdafx0cIUMFX8IQVqwUurgRd
9aVpFOkaTMMhE5xa8WCJcdZGi8QoO9PMcBL4SWyPTsbcj6jJOlUqh8MT7VAQktrqSjG7ijL+taNO
+JertjT87GCnerwB4Whh9yi81fZUJSh1TdwzJtL35CSasdLGRN/c399+0h1IJgKY1/pSXMdv5El3
q1VPTqawm+QGPzxnINbkE4hsUkbBGLqt9qtXhH6UslfpIMXCRz7IwKYNvHzPyTCKlewsxeFPFwYS
+aekpl0xb0bVF5Jq9hlhm1QDkwC/m8iJtNFAgCRwr6g+Sh73VUXfSCsfUeU36YVeS+V9b+vIOWnH
aKirlG7BlRuVqsp2CYOs9BgT6W4WTEcZQRYE8sR3wXZlVPhn1LgNX00YtDLOe0dDVHPRns5bX8AT
spgfLyymzWSHyUiqoCM1dF20oNQqj7CRewc1pUx5jc3U8CdgpLEiN7y6F5IZGrWmoh4qtPsBYuGC
QQOMLGqLPDnjqbxdiIZkQ2RXE9opohssNoUdIvLEDAf06IjwXMXU15lqsvtbJhaF2ns6ht4Nmzd2
eZGnuiTsPhWzQUUKHEdBAdUCWWNlYqvK7NTKdhCWPePjmiXVoj7SRKYnDuYUY273R8W84sw/12T2
BZIwJYFI7ts3X5uJw4KWlDqfrOx+Y+WGDR7U2/iiGISXFKd8T0m+8mzwTCCy5vUiascZBhW+ReUT
+LmieWjFAatdd0v6SxNKZMXpgPxZ22w/NOnYIxLFA0aqzmynPMbzaEYo07dKgcRbAvGIIH1vWLqH
b7VsHL6RRMiHgqrimTxwRrJKJimmP7MG2V6o0GuD+g9fAtAcU2vSVaVz+ZELxxRKOl867QUN4N7Z
tUya+03D3N5oqzE3CimmHjs1MLjKmaVJ2AjM5AZu3gOmhqZUD/2UXiy2HvRu4SGaKsPJBnBX3EBi
1Fx8B7GWfciTUxTRZ8tXnEGehGuNEQb9VwTJ+neyllY/r4jqxile8LlQOrZnIYAFD3dgGa9LTF79
AsKV+DkyvmJ2CsaIkQrTA3auMKu72nRxAUmYDubJ/l7s8MnhlRDjQ1ZbyBO2HihGB86SKqWOCAnW
LhDI6T7jEAydV2JJx8sdEZ55L9jKOlCu0B9VU2ZzZlH4RH9xm1kgX+XH+Sh4sc5eWx8iNslKbZ2p
aujPvDmnDi0YaVNv46PXb5QW3x1OWoCVkPE520ltsD3THlyyGYF3FLrblMRGAeXC6QnEtpwQ0KfG
GAGo7hxj/BMA7lI2uErYP6Y+KSKb55bv7lO+PTSMjusOC1UzvpFR1Gy7N30TQ1GpMvjSA4v7mFEM
V+RGKj73tFEkmvCM7hAJAxhIfQ89kHbdEGoIpkzXUzjILOK72ELQu0eJdd5iqZaaLJ07GlumEvXW
O1brQp+HXg55B23upk1fRVSvaHL5lRboNpntQSR3H/RAd09nNjG94xCVMJn1x0oMDS/YmDPCP0MP
hRsf4efY+mFB1BCwKtUbCd5yNnh5ic2ThFzFtSosGEojqCsXl1lx0LeuC2g4BIFyf6+k5zhdVGRS
12X3IxRfAuaqq46L0MN8OA1JS134Ddoi/8GgHHIMwKVdmJEvqEhQ3K94LLUxROE8PMP8E9Ljz3PK
oChdJXKutyg3ORfZaZ27gSWg1n7jZ7hHsQDb8m8/DJcvA/hA7USW5xBlZ4KPqQ7KFgCCpGm0Yutf
VgqxQsC7yEBrHc1gvv4CjQueQXPFwXv54SAwe88kUG0SIlg9ldfjW/vOwY5dxWt0EqRKUCpD7jsi
U0pfGidsqjVK7qDXapaJLdfdcWjMQe6q2AqQDfdiUqbPlLEdGtB6dEN8sSrMtGthZ/xGtRs+lgNk
mdsC+h9ONzc9EsyJnFiHo5hhErlpl4+UqJvzB8h545JJLrQ+37KPh0y+Sathe6LmyK3wCA1KgfOq
8+ggjL2W4uy0sai0ApzG1maiVx4rKy9RSNksBCovk8ZsAV9FeymAoU1VyBJa6fhDmX0FEZIuN2b6
2NVL6nHI1e7k/oTtmHnvq2tIx1i95S8jQyugsMdtP0mXgeqknmEQJQ82PusX6DxdAlw7Iq/dJsMr
ssJXViryZ1LKtijm5gC9wYc2iIzHJh++OqZBxw8EftYiYNt5G6DLufTV6qVeJrCOOZcnMGHSat2l
uDgwLwnGmBGYSPMrvr6i/0HaSxx9DNA0FMzrvSmQ3/PIk5DbUtdzDLnURTTIifrNmhb+AK1byNaw
9tRM24OViSAab35Yx0nhOAF6XqA+/VdOj9v8zmNdtMWx71F8vAOvG1jZRXVHh/hfR+QQjUh1z73x
yavx/4tX5OUmZxLrUej1jEicMqmDdTRufsuJV3ttbQXfAW+CLRY7RlxqIKrPFRa/mFOvzq0/2ST5
9HX9RQ8y/Fp0ACLMtTakc7W2y+ML6LIV7yU1nj41WvCXWOZP6UkeFFH7CX4V77P13pNtglWbpevr
7AoBVN0EUJ2XGhfJ3+6NC1THAhGJp0vPr2tLF5w1J4ADbI0AujMTNGyM2YImw6yZ1hjQ4YqUCYnn
dNxcL3szMIXwIZV6Ra48WNLEGNVTKf75/39BjppSnGkDXwOowjwy7bR3ELbhVlAtSrb78qzNPp6y
WcJfwAGaMqjzgApSXtm2w7dEdcsng3pztFYLiesorfYGG4Ix2nTplHknW0F9Z3A+K4SGezKD8t7r
5KG1DKjonsSC0h5/2S4sigen0mADRSvxqUEP4VyKb/teC8r874yBdmzJ5ewrt2uIlby7iJhyFYz1
ETNuMkpkLyrpSCm8UA++cwsJqbt4z1YzVstqdSgKmTZq5SmDWRxE3Esg7GFB9GknYK5aBKNk/EEQ
cULYA8cv+bdJbSzCy5PtFkIoIgAdf0eFEtgvFvlo8vGyCFXIF8YAWYilMP4smDkqOdPMzkQ6eZtQ
zTtSJ4REqiYbVayyShLp9RDuUjiMFxJne8HIWfIbDDygBSisMoW/c+3a2Ks/PQbO1rGCCpAI5EX4
YqJ8mmcAw6wZOa4jfExo4imk744Mp59b0oPTCNqYZXaTc36LfCkQOoX/t0F9rzcNKTcYJf94vNqU
NMNVELc3q+c3xEuNe1J1EnPJ+exN+ZMlDAbwzC4/VRH1ExS2lLd/hAFaDH2YmsjCMxiGo7pndmjq
ERI6bw5ZaJ3aU2e6AsApGW7l+iXem0/hDU/PpbfmV+B7m8XjYFssEYlfa/ISwMlny/GF41vqp3oA
zB2e+BBz9yyHM0NdiQltgJB89KXt0RbMtOsANxS5bQh4AUTFhoxv1IOQU5bXNbgc7C1e85tNPhlt
qzMB/IvNcnTkeQuOSk+mr4XZkGAQnWUBqmyZZ2UiEOKsUQQtLm+Y7sigM4BdZ8WY2wSb1QQ3EslO
vrRNRhcxX61ulcUM3WjQjQCktPfNp9pDBBAqMnNLZLr1QDy3ENuyk7AIhcGH8rxZxNkTjs8qguxO
P/RNyAJ46yhcTqsfJWK/g78hYuiA65rHYWawH0LwkTBJbvmEadrAX/l0ZiUMS3NY797Z4v1hcyut
HDMh76rarn8cqhvkOcDtbSohy5y9rG+rasDFZrdH7MUyyQ0yngYM1K8BOL1fk3jf7eP8jun8POm2
6xOdOfNSDRBehrNptnGXPzN5RlvAJM+aY0nlllDU/ylI1SG+HhBZv3a4Ph9K4s33Y4C/AZuBHTvl
H2HqloxCv0hevM4u5URh65rpXwzo6JGg9ut6NNM1Yu3c6fwy27NAB16cE2/CFBZSkP30kUX0w56i
KyJ97p7BjgWnmOJxSfy7ugR7Hr5cGTiFd4G1Sh6VglEqkeztzCv7CQrZi3Xj+pkvMNfUasXfpOLd
SMgHMVej+jEkqyqpte3IJ20dkNqoP55phWwpLV0sNzjtePTdGGgNXCq0hM+EVHR48p85QKsTQykU
t4lMtO+kMf58YcKHW/3gJNhnRnP/Zh68E8gXuH5nWTxWbKUtd+yYDO0s5EPGcoE61tVSogXhQVI2
MpJBhOdXxcdpbZ2OyfglESlulcPLXfL9WQrYq2uMHovwuV1KkEa9QJM9SFNnv3BZLeVKVN+CFTDJ
1j5GUos0tET8bRSnotGFS+3Ks6U/H/OFqfqK6LdPxwG/22tsIn5Mh+4YMtsCy+RF94B3vO4SqGLV
+7Exi5hIkjet6aiG7GpIu9loajR2tbLyoWoEeXjbnwpJlfN9fwklfaqRHROF7LonZEolhPWjcIdH
oHLF3JLAYS9AfMgucZlT6zbnIUeOpmRsvs3/YKfaFhKSwYZwfsiAhJWI8E2qvXqem2hAFpHhuMWc
A4nkF1IDCT+/2qotAMG++Ekxp8VENVXrrYu4zYwc2/+LRAwIGvLvbMIpi1dusm/HkQZ03AAIs3DY
YN1iZlkAG2nomVQ9Ak1ODalMRWOS9iYyhzcDXp/TES94dFlSp9zyQgLgLAWNznoOcwvZTBQMHjjI
vbe+tyDWdty1LUD6el0onrzmU7PGhZseciK0Ajkn1JyWwGMQaq1eYb/L6jR2l0wHl7Gr9cVHWly5
YHs9nBne4ra9Fe5232WUHb0JIa+zQZJ2+1jzhPwFp9yHbufOIW9Rb9h1mf+sO0f2hrO3pjsTuMEL
yj4xPNEpOqOGTr+6c6zIXLX/qsJNmqvr5pw0IQgaEuuBIGsW4Z1D2K7g2g9F2DhRnQY3VpuS9vlO
RU2a0MGPEUpZD0iC7rF/Bq5tSLKKE4dbemewzb1p3e1BADvrjPHy67ajIJDlVftJrm/WZTkdImAm
fKskyXtHvDT0IXM6x1P1MdOspnx4Eg67DbZTHxAE5YpRgxMwhEpfISoxpzJ3VgqFVMdIUs0acmVG
9e9kYV16BHGI/P60/uiczm4jbgnJALRBdSzNvKkDBkafYIBMcwqSVp9ttWhb8l0zen/doXLYiBgn
nArKGS5vki5b4uEy2EjTehfu1/45vPsTUu7mHv+XPoQLfJ4BD1LjE7ATZOLrsPyfJjsn11W4QsHw
bL0PxhfAQ65YXvFlRTCrIrw8uKmjgB5O1Wbwrke6MWTwFZtX9lhEo3FulrOwsQdZRwDUt3unICbw
4bhrnfanTJDz3+boSstsoYxEKSlJbkZoxqCXNwLbloihPwVdDbZXn/dV5VDG0ACV0LEzg/Hy2ZI6
585Fi6Q453kqKaI3witLTLAnV4IG0XrRGH6O/wBlm3rYpgElsMRPQGRS8Jc1LVlY2RBKOEtYkaxm
754Gu/yPgNNQ1jSaFpO27gKfEyxwlIKYE68oK/JwV6TKridvI7t7h4UahRatvq69GR1peSpZrQM5
oJaY1KKdsZBaRn3HpJ9k+6F+1j6jk+SKRPDy0oyKt0fpq7BWz6guBfjhoIYQnuyn9PXnTLLx//y7
qlZMBGLCQoV8tkhSIUUFg6eFB8kPnlRakbJuFzdSdRqA4Hi7ZZhgYAKLn15A4rkUEYHdOpgygia4
/Oukcqiwilpc/PogBumZrZ5kO/U2/g9yi5Tomoxo+lGZFGVVypzkwzfenwKNWENtZ/bYBgEcKNuT
vhroJJJ9MMSm4Z+5gYuvqOObKJA/Y7c2ZPISeZQcHXgPKXwUqYV3sWs5vwoGsDWdZsX8myN7QfUZ
uSl6y1RoKoSNtepzej9P5CulyGSMoBALxzocMDKy0/CxO2fQ7ew86Nbli0mc7u5SLMwBgG3fcGa0
Bn08XJbyHSd24MPnVV2ncro4fO49Q3bj4o5XzPz9t5Erf5Rr1IysPgKw7V5JhxjBUzArteD+nyW8
BqKobyxkPvL1IC68WARmvUWhLQnH9NAmCK5P7Ahf4nsGJzuo4tZ3ePVFUsm02dAW98Lyt/G/x8tR
D3n1OBEHNvSut8HEN9JrQGZMthDWczI5r6eMCACENhGrVCObboLVHKjx3lQMxAhsqM56nO9mv4A+
Jx6fncgO0M1ON0nKnkVnbBfCXBU+bo/XAikIh1XKsD1T3sgn5TmE7E61DNBIprukCWLfXzmoawrU
Nc925QR3gMw1ePTQWbPZ0jgZbxhZEi+V3CMEo7ebCIrerVp2TKA3DW1usnxeXCEaUFIRWpy/SV+R
Mri6JiWVNVWnsCeInfBQ4BOI9DihwshNWt79+Qngu6vA5VSSGiBpEhbP+9owkpVYMvkcSOGO8cvD
o8La1itTJbaKmuwDM5+JPC2jtI+gtFoNXYYA3tB9+0k8YNDNLxrcsngq7wlHgmi49hes5OlRuYMM
K7RDhDVWsY2gW7LBriEgvHE2q/+sOUutDXT8wnTV8/y6f9DrLUj2m8cOu7nqJbHDoQRRlnNR2tpd
eE5UXE9kYopq/N/6YPNmGXjXYD4uB/og8Y7GPl+cJTUaSH7NYQOq3wGRHsXdmg6MPSOk8wC49Mp0
Coxv0z7E5+c2kPeCta7oZ1/Ow0lOy/eGv7R0yJBBdCwEG3Yq8W+VjANDIw5M4dAlnP0naSWpp0WU
ioQC41VaGvSGoPlQFfcjbXYLwqVO1J/GIDOAeYFASSczsv4bvRJ+3DYBt1hQABJuGN2r1toEPdyh
wPTwh6KOV6bfzAyUYxC+IlnoS0xyqoMpMTD0V6XUbzPFFhFHjbVUOnX5jTygzHOJNIrrOwt43jmk
VB/SQn2ozD02ceqohou9/duOc8oWZVfFfipGxppz2xr/3ln8ry9xeckq7yeJ0pC7UkHhzOPub4Ux
2u9CkpPq+NiFgPB2QCYA4jHJAkk1dmaRC4/XinHn8eFHCmHC+krgUru4lkEYaO+fiqoTsicB4qyB
7kuvIle5QUfzp42DBrrv4rk7gK9BLsiq+dgvT+WBygDcJOrR4cKaVVj0Rpc8dHtQCj/7puF/b5ls
To7tpHosHhyaZPiwywoEbpyZLEEplrYGlzUoxZo1Evv4U3y1jWdP6UcWR256La6vO5W+rV6n9Afr
vW6EKZ8lcL6NHAK4p/tna0V9tKuM11tMG8Zmz8oamhks0ucp85d60RU+Xj1P6QU9Wir03QUMbLGP
fD/NjDRwDDqtkXqAhX2e+r4jozFBECxaYXf251ZZpW995zvoeVrbeskxXYHdQ9Uo2kHwev6KKelW
ga5IeTH3g0GfPLzW19yiXCGfTA/Ic9prhvfx+eayIQwPipGoFESU0VoRKKbAkNLsbJ4eR3/lKW25
D7jwfRUeZKcVXNh4FxZKim0axsct+rY2DactQkN3dc4Ewdx4K2bzCba3hoYXfLQa7XEQo9gbQdHU
qZMaUWPJW0f94vfe7vrUO5d24fFMegWEPoA0R/ZY5gEZcaDog/CssBIfayQmwkVjW1QzR1cyqskB
h9Uop5jUCqFv/PmNDapcGk6JiFzhyRSPzH3LN8ztL1xy5kyk/ICyTugRFiV+5vZ9sLK5XnbYhe7I
hJOISMLPsrNyxr+e5AQcd/IciXCBCXpm4C8rQFzc0PRqFHEsTsbUmSeXxPXAknwWAM1sPFCK2fE7
viImJ4H5UaDrvEtoBWFoyvxFvQNLfU2b6Sa01xAVjyozKiGRaurdrR8IUN8KaE0cX2xe5mRj2TFW
vYLPwfR+JUw165OjHMEesmUIdQN7JnYWuGzQiRwprRoyn0jVB4O+N/0KJtcIBjXKc/t6Hd/wpAHQ
GaXjRicbJedwK6dELJy8dFtQq9TqXzsYtvlYawu2TEMPo80xpjdlrpW4bj0rerCVLMHmOloj9c+e
UbM1bLzwsE90L4ghdI1rb7Ov1vDjEoMhsHja2EptZv+uIOz4bPeHbmQ0jT4hTqNVLAI7U4u3Q3kk
iNP7DxoqTT9t1oAFh4eh4NqkW7Ommv6E4BD4xJYKeWFanXgbFp2yH3Kz4nYf9YhZKb9ROD4I+/vV
x/Em9IwnoH21IKQB0RneOLXx0vZ+MSrv4skXgVEZ5EbbVwt3etJHI5dKtCgsVmxj0EQTDoy8HPja
yDeOL6jVX5rtTgWLNnhvHxH3TQorfGgLqTl6mtgcUvsiAL/lKUhypqooMNGweSWKGQaJTskEUQIk
eFsNpjdtlsmo8Iy3HZMBWxpmZsfv85gu8HtubRdvc/KQSMdBR0PLiPB/EwWda/yYKdzkPd0dGWlV
T3iJJTcDRvgS4fiDoEZWNbIMaWRSjKPSGjPV1x32pbXCZ4/VgYFFpFrKIGul797m3yCCecoAb/Vu
JJe4FW9B4WX9pNPsInsEIkDFJU0/CVwlgEWFyqGU/30ayTACi9eH09Hp9w9U1zUfNkTFBg1wcS6M
0Hl0uUM3sQ/4IvCS0EaTQZ00fK5gbbeWsC0+q6O8NPGJ7UUOm2rzSxoqVpjuqT6saem9dhHrKmMm
SJaJ02CSg0Xpry1x4Cyjd7zf+UXwGcHL3oAQSxfbnhGtqfh8HTyava2r6B4dOCCXQlwzVOeF3l0L
XKu91WHTyfmy/p55z7bh7v5hiH4pUJHjFM4jFoDztzVC4hv+Vu9+BbwpQQZcJQnXWbo2Zz9Zyg3K
PjP9YpyKgqvl9tKdKheu39z4zNwNMhXCgLXrXzHCafa6AvYRXCFx5y/jXe04R4Q0+Uj+I9/WmQAm
pdHT/bIs6tfXGFAEbhQP7xP4iB6kMaynP4hBZIHv+0bSU9zHt27+Cqpl52tLlCdErHT4Z4bLdqeX
C0BpyHGvXJ1zBvDKnwAHLg3uocb5rJxCqhGg1mplxEw68FdQKguMwCgyY88EmWuNm//KqaeoF6jr
Jx/Q1dZJ5K3bOzRdNhV4nrDTLQyeWOv1cEiGYksbu5yvgssQiIOAqVAf5yeYtUa0DQPGcUnPTfLo
0JNbl89+9SJGF4w66kHtbDS8OzWRgmx9+FDEa1BNt/To/oQ8haxPRc+w5dxvnqBfO2UHhqLBai43
fpLKraAcnyjguK0awvLgEm1Nd60rUzbg+i4nb21v0nM3FuEI3F3K5pMxB3hpel9DrpJpxGAb/E7H
9vIp4nHcEXsCBiq//8RnkXmnnzI9NDrZmrJ3r+Y0Bf1vibdiEP4EyZaHVtjOF0/OzcAMUb+/DAGg
mUgzTlX/ORRaeDWe1zN+RItgT0ClLqVvmu/o1y+Oubv7C420K7I8z5RALT47s9+U6HMh3+bwsi9O
r0eVHF9va19ywqgONmHEljD9ZIqDnJjkF8KUBelqoxOjNNEvgIaK704IV3w86eACTy2Cj+yw2TbO
0nh0+1mJZq9AhkPu7UBkyqKSGG4lHr0eU6Ufh+m4UVIvKLIww61vXG5uSJiHp/Z82/HuCB7OwFG1
Hx8EoR8CQFedv6neUo/NCMRE8tZgUtaZRBOsbr9HCTofKSPpxF0rvnGarUY/T2cj+5K2mTIV2Bja
85rS7K+jp58UD9r/Lhm7fGnvS8rRp3mzT3YX8nNxtQ8NmZR1Bjhuu2/eZyXRwAVFRfuHTogv1vPA
xpqyGCsV7wdj9wkatmD7/WGcvIWCpRZmNee56S5PUmL7gSCUZGU1ZP5Ap0uKoGpI/uUmIqou0pQX
ZiGtRY1ooVcwXuwGOKWrqI9u+DLl2wPhaa0OAd+aqjwVgstBjfK+1V1N1mmsSxb24I0mL5a5e6RU
dnwkMWWqEynWCHH1VB0xA8UNXqmCXoAW3wSo7hA9dmEqUrloZ/K2qrl0ydLBZyRohYVLezvGA7nS
MPodOm80pIUfekPWU0w0j/HNJCVuejrY+7hvSiwH3clmu1C/UTYrcHNPtADv6JDv/35JocM0NE4r
mdLq71gHCQv6oC/EtZKplXKeFF1x5K5outLywNlk2aMJuYEIgCYKzFVIOObc91/7v9PLdpg7DPRL
mlNb+io8J4kSmzYzVwMFTVVqTL1k/VmMYc8Gfq3g2luOPHZYbz7d2wo3Xjrk3S9c+KE9WloHwmYf
BvqxGMJb4iaqxfANWfNVvu0he8vBxbVkSy+A5Uc6EmRxuyVT+k0zIReesIX+a1aEpwhYzV6DzQ+V
MeWWhifDs6Z0ZUDmcNaJKRnY9p4Cptz0XLmXoYgR7sUUZIUWFH9tFR5mtxdDW2neNf//NTZy4Gy7
JpS+Ax32Ns89A+pZdTzMjmWhn/dISq8SmswxHPOW4YDTIdYq2V0LBmv27u+MtM2AJHt1bDKcSfV1
pkefnIr008rF3Xj1mQhChonYuxUNFC0VFLRjL3uYqZwJtYvgpyvAGKEal23e61Cw2c80DlF4d5Ia
CPh75eKQkVCYAN/faHE03hdtO8QEzAbAiJqig/qUj1pO8KWTM0IjSqel0fgXnf6KVHXqmiILBrG6
W7jdvu25On3Z5aWo7M70ssyb7Ss4V4VrkvjjH1T7Y6NH0yhatupRBXyJimgwC57Q5I2qzK+yrXTz
VCAf/z1JpNNIA+jSbcikTBhOqLZhfCG703J/+hLyOqnrV48wXgfVFte8h45rQissJ+BaDNIU4EGz
3iukl14ro1MWcOOguc0sqyCxrRzTpVp9QZR+5ognALCZ+tm/trRgUOTeD4Q5SXwDRCZCqGuWU0z3
8rH9+NRYuR1RVos60z0/hJxGGBpWKQL1iscII8iIyL+1oARR9iOu08tcqHDAOTgyjt6EIDTgZOaP
zlvH/fphfVSDXNoLP/73SHXVJ4RGxuDSLTlvcBG58MrpJb3P7iMShslBEZdZkZzp4x4wjSprLmKV
SaU5x/iPqJXd6VbEDn3wsLQQb120oAtPGaL2eNdf29odoDIPerp7OkodmG36fNo+H2RDfw49Dh//
9rm3+sRmhpltOSc3EZYNRt4RckS5da+ZmflcyGLyyGEvvCXpkUPV8c2bQ2FUY5uu/ZObnsPRfSvh
XOCKRzJYS8UwmvuaNjKaclb92Hr9Imxfs1Ym5Wslp8kJVVDXZpQEMNghQQAWcFyOyJIRhxABV/jb
tUiBC8TwCD5NGNwu+hzw965yraHKui9YPYW839ZL+fif8h2JKckdEcGzJjTH1PjzZf1DXPAe1ljf
Z7rkm35vOsJoQgMGki4Ts37h9LD847a4z+lsjGrzRdkErdb1GzvqEBFuqu7VpD61TvEgzrphMzvr
gUhQjsCgM4u3J5avZEOXvg0S6TI9dM1le1mPYq2eDX5x+AAef0AZdyFUmmYvIqHFUWBlSOv+Y2nS
n3Xq1IF8Mj2qxYlyidxYoIoR9LZEmrd7ecZ0XdYYNgKu0+06VQTakRn8Kh3C3oFexyY6N1q9D7Ec
De0GSQcUhJWA2fC/H4mZamECwXhesPwQGx9GzDPBBzP1Ec48wy+yBdghVolcSkX/xOEt/odt8NQc
fHIGjX8u3zN6O2fl4OTIQXF5Ib0R1r1GncmDprixY84/YxJra2IBNDB08w0YkapZ09pDHwQlNPT8
5T6ICHuAxUGJivE6awvaJtWwg5BVH8CiPnDlc9gZP3P4I41yF4HS3wPszxzrW7NDByxKm2fHn41v
EH4rLkPlah83v9xFkNM2fT4X8jsi12BaXF4VLXC6G0UFXkV/LdlaP8iSbi9Llq7Yxrr4+323oMzg
R5o4Mbb0caBjw5VTTwiVnLpY+CrC5mdF1M2yYKdQJLKvoDTZwRua2GOShmC8MUwZ6viVdj+eF/Ow
IfWQUBu5tO2b1jJpfj55wqgCSa/iWaXnOmVVbohw+PBKPd2NUzj+5xrA1Qj+0kuE12FXXd2xXZPk
tWHexLK93P50uMzMjcyYa9uJXzGbdNYVSq0UICqlfxxhHWMVp/gLxSKQZcAbpPnq5iREc6iAyNAH
dEihSY2aPRVZpa9eECp6R61wXu62RJbpxlZQ4CrDDfF5YooDTKyGGGNfg95sF939Xd8bYxpUCgNk
9k3nUL6oVT+SzJBmWuy7MohT/DMOQDcEmq0Ai6RlQ1hwTXBBrLgp2auiMir7PdnBdL4IClQBmyb7
mfC0AqR08kxpE8VV4MEl0huHJYALJJHUipua1iR8qNQqj6yZwP2/Vg3eOp9ZpNSN0srJrsr/jomz
Ucn5jF6DAtMf9yE4Y7TBYR4XjP9goXrnLFbKWv9CslWsxw6sVMq66YoVcrjR7Jl2mguCE9PFigLv
7Lo0sizNFrYDre41za1RiOLOlSuwIxueYsRKKS8XzkODh+37wMQ/YTpb7qDqad0n+zqx1olVRact
6/cn8wqpeBshGlRx7YUmI8iiMsR1M+gXy0B9nLmWGxaErK+h8RVvnshAEE1sNxUpnRKFyl8uqMyz
STmCKObrocu3XTUe1u+eDeodZDGrDXma/ZVhHhLmaFVXoQ0DnOicSIJ/6AAnweLfZPDZ1Z0IktTm
d0aM26FaCsX7gAOI9uRBdByV3ij/7I5uGh1duRMVruGY5SMoIZnNWZDm4YAB+s3FR6xkbn866usg
ReUWqTt9MFv5CVudGqCnVVcQ/QLLf5nO4KwBlD192VARGDq939zvfPG9QoQj7IckYi5pJRcB338O
ib1HvOjiK0qWMAwDLMhZL/822nurKggQCkpyZvzqJLJD9iIAS3oAD3PGltReES2W7mfCdTbfJN9z
szX0j4pj9xBvdej0fO01VsCS/eRW3LMEcBLGAawEmq1GPDUz2oTltnXrlgZuFvsW/NfzAk4sOy/C
IT9BXTI4hoCdVFySIWFjqBnbcJZFrYKxoEwigxEM7KyWcA6ZcK68Lk7mJxQolF1T858jWXsdb89l
2HS4G7rn7gy3GEn6tPuUDWr8k4OJGXrPXqSa3UhyAdDP6CyoXO4dh8w7n2sdnUexqGko7eQ5wdGN
YRM0kYN1bxM5/k9/uCe6YM/NxPC5O4QX7sHF643GHftogH0kiD5LR/u6ukY1Gf6Sq0i9rcH04wyS
Cii1kLgq/i3q3NsSKY7sEL08zkema82firde0CEJn6MNW/PwUnDqJbdVcldSrqk7mbTmMdAhB0Gi
jYuLZri/BGWhCSAA+1/eCVyli/FmZVjX/BbtAwgN/89JJ8M7VvpwIk8eGwpWM+jRG9gwOrKv7RF3
QW6yE39OgLSs9qTbD0xpEv7ISXwYlquLr16tEWIGFTPssHY86T8tlQl597NQl7ADZK/AutoSmSTa
YSIgyLmDVxAnjnJerPEs3KPKh0mdpIJ0fvQaDAqNuxXrnOdE3bXwVwiRGXy5V1I9px1V9wQBAA5D
xKgwOed/SfO8KoFL67qJ/O+1DrGGAx1/MXT2IdK9GC0ZI2RoRy3xmgug1aGqkZogYKL5RVPNii65
MsusRUNlfhN757gElDrG5XqgK0VYQJI8CP55Ll8imqddqh92sgO1l7dXIJzJ9cRrzH0EnLacA45m
WckqaWSsStYQ13xgeIte6Dvqr1FeVJNPZII3DQURJX2qnId9FNFOklfr6wyhyqzm+VP79+/2JX4g
qZxRq9OURQ3R6/y8286par3qo2XznXFsWLIe7GCdkXMzd4NK2B295MWmRGdtpF8tmWySdlgMDYG3
mz4S4+dGJFRNmC6Y55NtI6a3634h296Id1awmiQrB1ycrDqTiIHDQIebubbaMKZcOpcPX042IBY7
0oanYtXpc/q60fHVAkr9G/vZAOs0lC6WA4R423dIVqFX8Yj22LMpk85SBk4V9cOQCz5MvoOtlPMr
Q5JkYfBS86U2lFICzqYlq13Qt1Vsf49o36CSGoV2kO67VEnHtv9xAqWzSTv+hW7MRpm/o69wX4GW
aRbvIs7WS2t63Xx+nUR0cVmEbUAU2u0Ndt0OxRa8FPUF+l20QbV76TH59cgC9ZSwmt17PI0+GGGu
hbnt2DvJNI/ZF8B5kVpBO+ta7Rl66pTp0TxhWZDD5flstjFF4Mu8sCKzxKXHH38tvtDnHAMDi3oI
JFefFrvKDRRj/5Kk1dmoniJ0QyKTu5w8eqIW8eQIfxrtJw7gbzvZCenKjl1sK3lIF0H++Lf4lS07
RRKsxtmPbu6nURco1fraixKl24JX/bg9/svlHoFmv+HbJ2OlDdGSPfet4x1bZjFR3MOIDPsOGvnT
5z3ChhksjkyT4otqNLBByXgBdEleBoAXGCslN2dJZfN1OvYlvk49Yciyq34NeyM5QNy3MmQb+YDg
U0FJBjxZEtk/jrH9+RyPKyk2yOQ/+TN5BDRA23FxWNpjGktevxtWNKu32p0+Xm6jv9k1SGu74GBy
tB9LjVL97cXHnmPS7O7ghIOng7ZGWOlBbslCgyXpvUynDkcwoqjPvt6H3dWaCr4Wmdyz3gS9/Ap1
58Rpj9wBkEYQsxxw2QR0pbyljv4AvKnV3hsmN6eY92BH4OWmHdH9Z00Xp8WZUoOcYZM68jZGfLPr
JZ8TfmNU6FXcQghm/4t085n92bUg9j5k6pbwvhd8fcw6c+OinXJi1y1sNdg5BusElFQF8/hg8YNI
mer1nZE8oj3O72+QTHfTb/qwfXXdWQQS7lGrHxNMfs//hkaaMUMi40fEws6b8HK1zfBBMNiX9ALc
GHQW+fyl1bWZWZJPngnELbdQ70ltOVOevOu0HInFuFYiDMnK1JkdrbnxnMYcWjIGeU71Zvebq3Ov
bocj5Mb3xxzsLbmW9VV4w7qJpTJzC15TK4WOkzLhLowHeg2Tse6F6XZHSMfRQPqy6kd6U6WkfQPb
9YddyG37Cxc2hENVpXia23BaVpcYOQs9myUjyTQ6AmfYYNu+jln3ecJOWEqvRcQvbHd133AoOtXF
LRbkUG6Pa9NhRI5RD3B/l9jk7YKgTRY8LUzaKPZJm4OWwarYxGn7Erz61vIru9U63FnOlrROd/gq
FwcImszE0xWd0Jvm0pXV7NGaDDRSOUJy8rndUfj+TQH4C3Mfv8+qZHGxARPC/YZ4Mc03n6AAkkSh
REwVLhFONsg1HcYuNBhTxZfUstVUCYSn++pu/kpNvertkUQc8ISiWGLaQ8wjYRlHSxB9ATcY12tx
xAp6PcLGajVqKIj0dtUQazd4z+d5xKpx/DEtuQUxv6ctD4Rpm3b9AYsygiii3+ZDEHe+GRkAtV/o
RnqaJm82N3Uy+mgqwU5qsqERAbJYVgtPZDXCaHQ9jafa1ZXPSfn3CnpyBsAkp6G+tT6U5j8WPdvK
JAalKkwwbnocnE9LUC0l6m/H3UhpZuI40raHWZSFYH7sLkJtuVnnQ0PzXpAqdL5VUM0FMREZhb4n
l/RV7EYRsUI7A7O/n+ejcCYNcjvbKg1vqv7zuL0WowX/UHcUT8UlDn9yVgvmqhRYoRxrSXqCHnts
CAN+Xy6K346SltQU9V8I1415tmVSXspT9+WYQ/d04swgNIsR4DJlVbNX7l2NZyVxlAwRW4hU1PkX
AJL8yFn1kIQAoIy0wbbWAQ0TezuaI77D6l6a4SpprisePjAgoi1j0ZEBpJzwX0M1Lq+EJ84aRlw2
asiUblhIEVRxB1AD1nymHPfCVj0b8qjZGOdTZHQG1N3+pHfAkCKB52Cv9Psi+Ox2s0qifN0VbiXH
YlOfI98IDt3X5Aol5LMOsYLvO48INx9BdUyIG8osNRrZS3hnjFSHdWXB6yxR0CCYkK0O2J0o9HFX
8LmUI0pjL6Z0vSnGNhh7SWr0bHw9O9kSfNQKsSNVWY1ZBl3+fxEQIRyEy8hOlCecOJ2g1wGmh0le
oqA4l2Z0mz4MUdxTPPAF1qNyGTXNvSbAkceH4IT3llvq2oskQ7ZxOHNbEmxaEGyA40M87Uw3v1Bd
YklhxWoOL6dzIZzJXAcxdu63YnFyW66LIl/2t7X5UAcPeppFMCPy02/PJMrkgXQhP5GZqVH+AswR
4mkd1KZoesEuFsKAin+6ZEdUzPXCnEeU00lNIaEYGMpLbTk3NY4DzbWXrShy3giQ6rGqMnyzihpi
JG4FSqc6F7Si9TE5XmaFQzXbqx9kpOLv/qqcRgCY4PKIx7KZAUajMPm6/8J9+WIS9qJR9BuoCnP/
XooGKXWdQjOuJ+8u/K7ex4SqWOaY/SSJ1bagSG7LE7Fp0C2TMm2DvZy8SG2BvYhNKqC3xdph6MO+
2iPLJu2EvqKUBma8YCQXw28fGE6QAaEu3gUPJKOkpDen+9B7NoAcvSxWkXooZnk/K+YB89qbxaoQ
eIkil7/2bAmf//zQN1dtE6TK/MOQ90Lo1R8Xqpdkyz/irdEet6u/Wp1xCJw0q0jcMTQdi1EK9B9D
CZZYDpFTGJUIii7gTIHqwMCok3soW1ZFRhEkMTu67uLThxHn4tw9VkdjyIwd1VvUqO+TwRJqq8Zt
CJH+C43HH2zV3L5HRqQxEUZcHe5hfjDgn7qoE0kB+Ts+OyHjPaiSWefie44KYY8jKz/0x3B0Ikgn
7xACPXieRZD1B2pFNTVbriA/vODX9Bby3/nvGQDUJRWQ32gRl64JVRukTD0bpmJIW+eoR6SmgYgX
DmFlmaFSEhOsgT4lm9hX3ChyjVefAch6bxqwV5LWgzW11AU/LdSmId6G360+3nn38CrN31aXvttw
5A0hNS9yZwKXHBGCdkwgfM2rll4M82cj6QOD+MF0jCWpJtVswQxhZhNGSpdNJ7ShKoejGHSPFejw
F8wh6OfE48LJEab44wM95BGU41suON168tedzS0krDq1nkk5RlVeTFWRV8+o4P0L+bnmmTC84a8w
gtkKMqZu/GcsJEfHg3Cw33+ZOr+BLOAqroHUETM3+AVxgG+T5/7p8onk2YGr0BsZX67hiElz/38X
WwsMIZtcRXzfl5FAYZxNaHDXPjSEOu4s2rvX2GAEmPpQpbJxQvHYjmGlSfs8afmMjiC2QiKgvgen
x/aGDlbgmO9P2PsxOqgE138r0pGXV3OL7QTOwoXIw0ut89FL9IP/sQieMU94Nq0uq7od2iciMA3L
859tC8+CndADXZzrNKaKNyXGwJ360sxn3coBEZW1Sq8TEK6R7Y+ZfTP7CkJ3WK9ZqGKGiqlrPl1M
wiY4sekExB0xFVLt8egH9m/wKMHbFA1AAq4UKap7KWIqqGej0cKdLS4zbVtqezrH/w1mSuo+PMMZ
zS2qnmGg++v83Dn15cYvZGe5bKwBSdb+2tTOzGpPs9jH8NNOvlRrsVmmhtLl6DRQsp+N2FfZhkqd
pCYXCSdrPGxhON5XIwrjjFzIWDvqY1bzHMDljtc4E1cPwuW5k1k1ZtrHTHXDRAlq5gHHbDnYbCv+
MQI3ORXXGLulB0xWQHGsK+qnogB+24HQLwprsfbyJCgKrr9SL34EJR1gaCkJStTGpii+HLlyzMpb
9lzMtu+uN5v49gVT7kd2p5TZCkrKe447EnXvg9z3HMXQYq8/wjpC8RiiWAqWbipi/bgcnr+w03hX
HWePNkdVcnPJ9jb6FNuJsDGCG/ZcxO+/nJv4P1sB8lhWjaTIP4hIWP9ImCxlL2TSsLCeetzUyF/f
vO/wd8EWY0fyOTpjcyt4X7hdynZZNBOcyyIpJZo/1mMRCll7mclbK7WrXwxoLe3cKeBnfvwwbg//
ATK4qbfpIe3dxqGUccDfSYKAkK138+cdT6nk9avQJcBY8wQDlfWsRVlfLBWm3nvKzxBIgGXEjxGi
HU16KKzIYkqi4r/s7lSsNcikceXvDlOAM4l3qY1po63QuwoCLEAQ9eCG4pSZn5LXvPeJ+SvsPiJa
2ggr90cVJNBUgQU6mmCjHkF9CmIGEceqxJnn6IAJhfgz37yZfRDdKyEuXD4du2prADN8ETXCobSm
KSY0xfmEw4mKkW3Gn3c6tr61/fEPP4DPiNoRRTiIVUPPKrDOw1iY7VRoNLqavTl394L9w/mfsUqZ
X+PfburNWH0qtmhwFiNnkq/FQrFGPtLIjSRS92DKtHR8kr9Czw3XNljARQw3x/wCnqyrz0aaX1sC
L1yDvZQbyAoh9D9vAG1bW/LxIQq5o3u8RmaX/IW6NjBRnw8yNpW11twDyndqiwTi/zLyIa5qm923
JbKYvnN45zno6e2f+pSHIFAfkWTNBBlN4oHINYFNLQCjvipOM6V7Y+WkVuYh2lnFXeKHasHwMheo
kW+e9PnbKvR7bTT25r+m9fn2NXiDr0IEp+bKBm88kfBxD7z5E/Bly43I5qEu3KeIPmInoV4WY002
NlT1Nm9POvN9sAHkUdLQ5xWz1b8pno5/451mSOpMH710tqyOcAVuKv/aCAsfQc+esHqzV5geDo1/
/0/XB/SZohAvY5VuzdNdk7ta4ZI8bjdUM5l215zGMCZvTrmh6/gTHEUEoy0I0c2zq77U/YtLQsCL
BQO3TRN52ZvIxLKxszpHN9dDQNEQiF7AaoV/AzG3GC4v9d9aN/rNP56TBba8L3Idx5v6HYfIO++v
PdNdDTaj1/IhtskuF5UnRUtZE/MHqpbuTsJFq3Be8cG6hyOB82728ctaAnJ7zwuoYQh38L3B2IqL
3l1z2wVtCiI0YMyk2qG8fhpPj7xjSDpjrikN6V7pMsnCNmhIFu3ELoe3t7E9PB+5mv+EzZKBFeJb
OcujLT/0yA++xT85az+NHQlQwpLt2TXPVMQKnnOvmc7wacwb+p0Z6t7E7EAWAwKluEWH9LvqiavI
LeRu2MXwNaVnYqqvku0/O6U00UWXRknC4x7MqDA4fG983g55lZqiP53+52P2pEqsWN09Vwjac9i0
GxvuQuhCBBwgZIUGsHnmGmiDqoUzkPP9so9l+PXPSR14efyvuHAd6b/t1vhvnF/uy3iPAClxGnjy
JttWrYtNNFLaYnjKJXTIp45EOGtkK52c7h5juk5yf1axEvA8R5ZINbL8y2u2Akmwqh5iSO/aMQAP
+PTwuONcY0Rw+CupcW5nTLA8IXSAJmGx5sp0+OTeuX2TkpC8KkSZWg3OntI3fJihliIJE1ah2POY
lz2qx8r8OG431ZMDdpnfLgAzbFilAyIs8DaoRtnSoo6pMuZgT3M0ucRRaNuFQzb/tO4/H8UYLYnD
/eqW+iHeta4U9571AC3mp0rwVQWh1t7QsUYP8kWGcwzc/ZguwdJdffJT0I1vV60zuN4Doi1MbOYa
m5W/SFlLCPoA7flni7LxuVu4dlX27Lb51ZVfdSw2HkQONOGy4I5XoF19PhqfCMyHIyiee52w1jZq
vS6yBDPExMjdk46CbBnL0SI8EpabRq/FOdScFV3eyUVv2+fhMVzQSUXVsGZ9NFtk7ysPIYK5MjLj
z+610B1iGvN7C0DtQBtWFJf8v0JOiaTmi+qdZ9uuurYnRhFqixcv6+VIldNoD7/v7mREEViPGAiP
B8WLqusseXa5Eadr5NwjrnJtxfQuifxRFSiDwfCSxJCFZDPc6KjAEW6vUaaVH+t2MxP8Trtaezxt
/27WJE3cIua9U/DRPGOtqiQEZ8FVk1q2b+4bbylLDnyzKr1GISrVNDrXAjDFqGmvhNVg5VUVu+Be
+cqPXtZq0NHe6OVlXEXojP0asuO1TmgpBjfYlOdLwla3fbT7MJ76yu3CX3VBt1g6zYzglFeU+cr1
VqiI7VUj/IwwOooc3wl6EeCF8bRRuD24fHmcpj+v5CIp8G+se8ynAKc2qXB5APkB6rvGAM08dviU
Lj/bv+gHga+YIA2+6c7oalT7IJgHC+O1w2fOBvx1n8jThKwzxZ8g4Am8OzpUyxF/ppXySc/laj66
PyrNA+YgYyw7/eUktWRoqbdWJwqFUnpStKSHScIFkoSv/r/KWHWPr4RypyITKnv2s8QPPcu5Ev88
1V8pzbrip34dfFO90ZRRhbEQyzng/M6rpZrTc2OatDuxn6PtCB0DTGt0i1E3pfuT4xHhGubs55SP
AqRmhAyCn5F2Idl/DZzE/U/uQMgCx+jo4XB8mBy3ZO6XM8PGxtEhcrR4PbBJe2mFk6x6OhpH1/fU
frX3F4LfQbUUW08XTSsh5YyfaNAVDNcE1N3B1R9uyTZCYxKu4o6JiqtwEwMPt57hau+Yim2/f0lW
DyljI3hbxVFnvoICYDMISKt/dHaejUttZbDbhE7gn2sq8r3QK2g37T05z1/UcRThl2p9K/WIY5Xr
IGo25aUhPMM983oj3MraMsu5ube5Wcd0fnZyPEVTtdNbzFTCNr+QeRkQlDGk0QFQ2gXciwxUeOyQ
eTtJwbCDsc6winMf7bu3bSSg2bnjfJogWIcN4U1ABGer05A/PEbKdcbshLKYp3K2qacF8AxYCCV2
tQTd8IlQmIrVY8VVzDEbGvwe4RLsKwZ4BFCEWHhZEUmY/isHcXy67e+5rR4cvsJXuXeoTPx7+Ta9
pyttyugikk6Z7ijAEyE3y5kVpXWug4FwZda1EH2eHCoYuJv/o9n25DzsqhXuAQl+PYLwFW2QeRe8
TCUq01dENRuhOYv25ikCylYZDqqpWkbHntcxdQEBQNz7cAJOE7VT3nTSC0YaAvmNi+dSh3MEZ3RU
tfHxt8R9/4qWXRL6EyCnqbs5ZpTGX8WE2WlVnKyfAM0cibSg9F6efY1CMaPhK3qzMBYZYB0X86Zz
QBTSJBehiRoZP2fN0U2H3eOWNGlKG1ojJa7J8S8lrAoQjSjAazf2gdWAdsls4bUwvMmOpr6C3OCi
5GoM6pF+AOhqIp47bZ2O4R5X8bzi2C+n0ZiQnKSj8mvOaf02EbE2rdcposZG7S6WLd6ivxi7jM7B
oQ1WRblNgNP7bfUeg8bnBZFiDyluDV2ouzhtynKrMsm00KDHricJqjbPOIbCg7oQG/9Laoxr9qLQ
ocvc5S74G8U4Z+SvqA6cL+s+jjd637xudDZZEcfuH+Zd8Xvk7fCh7Jtop8mfeKGhoN9D7tVnW8hy
5fj8N1/nUueXB8zuo/nTwaL/t1qrUD2iBkwVgUS6QvXPaa4Pysd549vblob8kSMUiqUk4liOd+Ai
4D7jqKeX5NQzlp271m2mxM0daIn9Ed6BDRqOp0ZNfn+NAhV6l9bCyz2cMeMNEX1lDnw/I+0jI35K
FMVIwY5l7vesmDplnrI/Q+GwXHRQiOZavUEZ0DJBCx/tYqKUyxAL1+DlUJmtVZIY+NYS1j/kAT1t
DevxILp3n2kt2AYMZo9xGP3SJnJmOEbxspLmU9yfqMeA+j32PPMzANI3XHfnSIWaH482sCkz5RIx
vorMonKXtNvnFZm/1PqrgjZZqHHZMXmehUg4ZS4+sO4gWckEIBMcwP8C68SYMwH2/wfhgaqdPIrQ
boR7+U3wtUYUh8xNmxrndKEoyIOJXdx9oX5YDw67bRv8ytJDWEGTV9Tw5w6OIaMS4kc+Ea7S6Bck
ZW24DfqRylyqK74soqesr3kWj5Kl5q8vEiiGaUkvyLN1y8oBpC9v8tkpQ986h7hIhNjbZyttdjE/
HPYGbSh+jKPx9rUV2GKh7J995T9I1fcj3veMgwUOFeLiOYDD/DahyCdPXeSK9hCeNCPGQMqTDiVm
51/V9Ct13nriZ/+Y4gEmEpp+4vfkYd70rmgN3SLp/rb0wtBoucxeJYIZPDwYT1uRBD0ydOge6Um9
hq4sRsxVydnjJ3YddIG0TgvMMMTI53sW/xxo9qU7HNN08d9dv38Wiic5JUp3/GVBszLDdq6SeIEt
cB8oOOoZW40N8btHLqT48pc9SehnKAhB11srWZUPuhJSRG48jYn+Hy37Ut/7XwWHrf3/Y+tJccCJ
/FRF6GMe66jO52RdWlb3FXK5JNoBtrCYBfg3MRDi/ZtbiNz3mfrRqTaS0SzQkHMJkiXRHGXIEhWK
syH6JInq/jT3XfppOM2EfztoN6n4lD33eJrxNCNnLCI8zKk6xlfWbWecy9g+KTAM31JNY5UDKjv1
n8UDWbh/vEcY1WXxcPvWjPB56h9DMoul+gYJnXvzIn0WQIHDal+MrN52D60QyUGE2sdeANcbaETr
EQaFGliV3azBoR8DkWVli1+yBxlZHmRFTNhNMjzogj1D9MGj0y50jqEvs7Oc4AOtJVJN+zL0pG26
ns1iYiNfrwvqh62s9pkYM3GyLJBft2i5aO4WygPajE4sw/OR9TKABXPuwPOjojSMhLhwwm5hnF9f
gSWPbCC0zrx9KbbKgFFsa0TcuN657pVAHd9phBrgBiDjVv5we6mrHZULvlniH5RLD61txuM5iNVy
0NfnfLc/FQgrN7a2UBJC8i7VWB3G63CoY9wGXfR0eCDw6aRXabbR2iTVqO+/uOhiwTLJYoVBmTVB
KIsmysCGb7xl4mlV1cCqY++RM8ihr2eSId7r/ToiS9DV/L7c4cgkF+9pYI1T0QPI1qQHDjW5IpOP
qIP1qsQUhwMtUPU4YTfjFMsxH5+YSPy27azkrHtubPi+C4QG4220wWMFtEF6SGEpl4X4nq7chFBk
w0IdYEm1A7W6YDqe9eR7baSSTlaS6la/1Z/j9/WouvbSDy9PkfQSufDf1SPVRRPYFmLPoq+YNC+G
2Yu693zbJU8s4Ca9O7ICfGxTDiqFqwGlEM+NtQvCv3wIu9713TyclGnQJ/8V3P1ExKKQ790276Sb
fGAxqNr/DXi1soY6CsiJ4LFrzgVJoD7m5j8X8W/ptCrhGDWkYsAv3VXoWb1IiMQ24bTaKxHF9A+f
1RrMqrQB4sr7NRW4CiC7DdonlQ+GpC86y/OHJ8/Vf6IxW8Elcji8HDORv+xAgkdalK5PN7luF6LH
N5wXTZLIMbeq2u0hAdtpQVch2LCRfbF1XA+9ehCKYDKWhQBJIS9yzDLT5Lb33SIqDC6kLWcboANx
IWpnNOLG033EvqNdAOFwvf2Lp4xgH4VkHKdikHonpO6VEWioO5h58SW/Aai/DL0BSQ7n86zYj0um
klfh7QQDkD3G++tlHeSL7DOLS8F9z4Xp4CwFKtcB87aN5Qixo7axsSdxMekNP7qQo8EGVmeyl4TD
RTCFYBGrUea/UE0G+v/B0eu/8P0RRxGklyN/KHeZCJoxaSS1SXvc2Zu9w5qDO7jnT0gGj67DfJfu
niqVp0CQe+6RMgB0DYThJvsBBtoV99uXhI4sahhEZhN8AAzkMffTcd+aaAfBQuho3nxm+drQG0rl
2LXbXBiAO9+dMqAR7ZJh0eR9Ntty+sqwX1eeUVrXLKPgL0Jv/IlUHb6sPCfJtDFGjcs5eMeL2LHN
Haha42YGyW+l/s7XA1VhwNOR13Z9M6RWfF7lDVkHd9t+TEFiZ1wFEiy5G/ire2u+Oy8+RRdKsrtI
QvqGX8mWfAqYkQC5QGmF4AfHrd3U+eX7bSflLicaAsL3kjFCKuoyNX0BCqvXW2c4aRfrSuMs9E3K
ogBpDzpN60Q4yRtoddPr3wn/NbMgVAye/K8I0DZbz2FzKp0LWsxBAywYKNzUWKWRqsT1M+cpI7Y2
faj0mYIrGDq44NwUPe/Eia+v3PslkxC9HwmiHLx8tQYQIhDnyD/jpfIewzwMgOv1gOaGgzTWFiAg
6x5JgzEFY9UDOgtgAnGQ91ouNLmSeyG9PH1QoyDrMeMjObbZ03uCs3xae9z6ptmktfVf0MNa8zPy
vZxZnwsZw313alhYUmv8XNOFEYLHPhWxmLIjc/eig+uVJUtwxAIuXZHwKwYD8byH6dXNiyHYpU5f
4wofr8NuBUl5P2RQeKcm6vGaGdtkzHIIxBMWNZ7xAKdQoC/vVDbA2SqCMjKdgMzMrZCc137ndFwo
y6/Pwi2+nZVCuPSST4f8GcUzLx28n4pdekQEQXz6MoHfskk/bUbPkQS/wYRwLGZmKhYmPXcZgn4Z
4Ll9WAWMZgLQlD47Hs0VczMmCGT3vYfZjU+iBOePu0ydIIo7BdUDZAq+j90dAayIRL8aU4sfKXIf
T2ayNNYFGVhgx+YvgFX792+Gk6oOIH/++IZMp5vfeB93dVx7fqMFE3Q/Vtv25b1XQDo8jIDKKMFq
+PRUxa3Kdf+FOlC+xAWi+NXHZWkfOJ/dfVdRGegPoIdgGFC77YpleUfGn3Agw9IErtG53lsH01ht
+/0rtiaeM7IAvD5L02b64CadhS0WtLZxX+HWty8o9vcGi9Khh1LXViPsj7bW3evtl0g9fk3X72k6
3VItjDvLZWjpaTQ35PIYYYf286kBFaY/kkzGoxisSI24O5z74tBvpyLz+DEMxBs16hW3QuK/+B6n
lo2hGJRB9jN4eT57Lo1GZRDJHT3LQ9Jxr5CCZywvl86DdwR0tLOZx6xCBehgU1UjR2Tpi3Wy7ajA
nbYLVXhGxNxoEU0sW/cykqkDkcy6czGgPJqnU93hArFzvgQIZsPs4Ps1sr47vxPmOJqE99DexHwg
dOp/fgV6YTsRQ/I7955X4jrfimQoluzACqPSaIuWgk7x6p1xB9LFvZO2YVCmOeZu9bqezpvHEyz/
8IT+4upc077xek4FJX8MAMpdkNvOd8dHaZNIOAXzdWHvtJFB9ESlam6X/dxW/5RJXafenoXDxqw/
xMoxNOXFZaEP8TDpYg7e/hlEehtlq3oxjhwz/nyGVO71ov9nd5REtXy+4tLXLu9UPxIKcsjdVqv0
GwG9KqIvgTIlWL+w3bBC4y3bKJuOmkNI9I/hCIMrUsLo0lax4HmqDqVFFrvLBvAzexCi+/2girwm
e9OH6IDf17/V6K5R3ABHFCJG160uFJN4W98M5TPg9SW7pNC5DrK7B21GHFt67szi3xU3SPvoqbUT
+SsvxWSxMk56/AHafZItcA0yRV1kWTb8+hgs+CXTAq+dTeEhhBnkFxdMy5HCW9GTSlSVy7lWWo90
TY27PClldNgzOkx+s5ppmMF18iycfFOHH1vqCls9txfSXl4RERm0ylNWE6tUWm0ASQ4IRhWGgFoo
m77xwF0BMK0mIX52xlnDxdO3e5Z//TLjZSK3tq45hJCaqiXtVdoeQ8x+JpYCikzX463AGPCz6qZt
AFCrcPhynr8HYFFHQ3ImV32df0mUJAyJuxBlF1kfFS95WklTNCMvKH5d971LC3USAt053z8+BGD5
/1cBagxV6MdqEtXf9/9+DPoJhlGqTgy823ax2Y58YrKCCjx7UMVUbgKlwD6wBcrZn1QoqTjF5GvK
lZ1FwTa6O1WSThGO3R0kchmyfsL7kNfp6PECkQRHLbxu8gno/ZbeZ7EjUDCIEePCxMM3XTIuaF4f
mnY605HhIOfb0j3HboMVcgCQdO1ZRH545n8YebUFu2eEAdo+6dWsV7fiEZEvyHI18QWC16y5BG7O
BO/0iqTR2pDscJmpo3j1O3nUTnyOpfdkvJcKerGQ+WdXbc7KmMx47GuzxoiAaRHJG6umywnmK5Zp
yk96Qi7C4f6wXebALqnsHqW9fBCvtHpOmmbfwu0MmJTAm7kO9jKd63XFY0XdsrS1M0zO8PSAFoxd
yY8CfqOPxAJ6pCD52P14rZMLDLXDmB+0dnLKWoW/mEOgoDNIZ2QT0YW66LGZnTjKE1kSYxp/fe5V
dWjpoxYlcRH8N9QBjHWei4vgeDdabNzbpuJhNDXYiGV6X6OGDvCu3LAaC+3frKSqpZX32rJX0AIB
H+2C5rfsgzTw/dLfTcOfK/zI0kcq9IZYc/BxMvBX2rIm5oqvRGuxkyzUztOS5zaqPkCgPy8vZYZS
O3l79SrqqLz5vzytmNRyT4fS+COvjykqvpiG36clIFyIzOartnkUc+91D43brmclMBUszQTvQ8XK
RdhVvIq4qbOq5ZnjoQyAkY56jolHyb2eWOlQM3VqAhEs6CXbyb3/psnhorzHrAzjxtmjLwQ2CWji
9AQZjwFNIG0H8OsP9VATaVLJFGfLmXeZWJ+TToIs+lORqv1YW0vC+Uc5hCSBife252LmwLxXueHj
JCQPz1Z8srurPY+StZC9zKeYG0sFirzGIcGDhZTvjBdN7C7VxZtgUDarxMAgjOeI55gzhOwXIm15
ssuLOrQQ2OSrnQqARWtVD640e451LfPzWBpHWt2SSqKtwZfGNELvu8996osM8n1nsXO8ww4v4Gmi
4nr+Yiu+zT7UF/N37hpfFbT8BUrHdgEZUVb4yINBJ0CHTTnC9M4UYL/nCGww6/GhYEVF89qYVtp3
6kwoDzRHhHyaDlkrAo74QGg8ys662MPlhjFM/EaixKrLeNBomathF4HfUUWaDuqd5gHgT3Eqz2KM
JES29mgcFCvPeSB7MXyrHvoRZPytuoIYxG/1cdHQ2JgvEt/6u+lTfAL8WslJHAZBXu5hlcb/o7H+
cfmRRcvu2V7a3wi3dWDEukQmdWWBum+fGiLCeeeAg4lSSYzIjyaRUohfN4VTe4QJxxSkENDqjdMe
2TdfWTOjXRHsqZmppIGj0k/+xu55IDEwN98aECz6fOU2GDGrVBrpGCTeKTBNi4ZY79VTT3f4In41
tckZTGV0xtWuO8AqCnHkEHkmF5GZN7XZZI/ezOFFqJRRRq8koviPIL9qgMw1fUHOrLQmY5+Vn84N
iUMJgZr1GqTKAYcNAp4GFN1ybjf9XjEVS0az1C3N+0Wo+h+j7CGarGLsA82dP+dF47uHKnd2VNHz
HKqZpzrV5procuLYUKBRyEbkwx5uIUFBn0PfjxLdXGKivnxGDJ1DuwYRVW4ibh+JTfY1q1I7qk/t
Z83tygAo9oNiMBpjeU82uKGFeG42RkSogR14/sTh8puQPGRMG/F0VX7vZpkr4+mBZhFPOwvt7l72
5opZwQZG4DQQF/csw9WXbcGHVvCN6xPjKDBmrJd7IyMi+bptyhwe3I1F+KM/qff2ooYleBN/nUHG
I2MA2IXRHFxKjR2eSVYoftTihWhMzoI1OE+id0o97KeczMYXgqG05VJtYtSngD/kOD214vRaqfve
u8EypCqqXgAdejv+ASXNHdfTKPeiaxwEAJikdbRu181M88iKz4nn1nG7YblgWe4K4hS0PWmVbnWU
L78Pr1vwunLtHNaXgs7TF/f6Lk60iKCzMPsdgQIpD91/yOqR+JstKuv2KSS2YevxcpM/FygX7FYG
GRTwM0166XuOmUFdq8xy+N+PDgDxq9bP0nq7SnpRygPzkNhm1Bpk7TJnnmwAqVdqntqYvW+vzVRm
xE0+vf66jg2NT5U6L5EbqOqU7564EcuB5brQ9sNIFI7zdR+tHnkFw4/3byHBrPlZoAo/I6R1kBgR
3m53Hy/2Go5Wapp9BdaIiNAGw5Xruvu44uqUbsCyyvuylePxX64rEQG7mCKJUAu0fiwp7Prwe2bZ
0fjFIvo00b2drlF3b++DiDqL4NOSR+WpyuzTWTi4TIv+YerItCVmKedG3W8+Dcc8rUNMWYH3x/Mz
ZSADDGq1QV/vAz7VrDRaNLlq7RYla8KDY9hM4UgUBB7oe9c1QJJW38jwEM1oh4S5aSfliLpAzLCn
S3Z/UUkL/1l57TmhnCZXGhOtxzP11Qusa7c27U4Zt1Pg0rLEPsovz6XIv7xRREfdRBuD9OF+FCJN
7KPQz/bWon/ZMz03y3ZiFkejbIUVdjWVUHppNpTQ5l+WbfjPZX4wFzVMaOs/utIs24CquUZCJwr+
Ew2x00xY9Cy/828EejBFJYm/PphDgsw1nAzu/hePaAozOikcxtaxx7C+/zZ6+omIDM6vOhO8KqAw
0fDum5JJJ3RIatJHB5/BSLt8/UpO58vuK84i0uaLAoSYJ3HkHi3x03ZIDix5SCMEcYpA0VxGQFw/
yFZ0emuiFEjicqFKDByVnUvXUNqktWJ0PkMghc95g6godfWQEdNICHWMqT2lqV6d7xXpM0pDKhWn
9CpC0ojrygKfkYk1NklrzU+IPn7+p3wLUzvdf6f4jcR031jsjLgaEJgceQedUdRrgRjmc80G71YM
RlCDMGL1fa+dSlRXcya5OjTmwKqgL+rOAa/RJxzk1hGjPvUAovdKuX8dnGO1zF6tYkFT6p/opuTw
qYhk73pkVSa+TBqAqQ3JmWG2U/iUzi//zzM2K1cOAwjxkpOmlPVbEIMSbGsL5+J1LWhPvSpU/Hif
waUqOggSTEXmX8kLtegmFpc9PWnA9sCamrJX+8Nb4odQPGqaBc8uGXbU1Vig9ud7W9+bOqxaZzaz
F3t7DsViKTVKZwA0YhiX/8HPhI5fZDXPBG7gISf9yd3J/u3klWn+Dmb3OI4E26ZWlXg2OOylF8VW
8o7xLX3T2SC0Tss759N+eCtTutUfyO72QGTsjk0DLjnz+dbTSCsImWIDNl3cnY5NTbCvjXnppOi7
z7E9aF1z7v7mSBK+md2clkAKQLLBlBTGoGvOZC0spftOuNZ+BFfcubBcwIs+hgYxmgyPjSrxoXw9
dgxpn8eIPgyL09sWv2wisywx0DbyhG4T/FTbi404Cnj9OVCWQQYHSXou5hMaM2TEwbL38LLGmyjc
meDEJTG4ueeZ3Ky85TxWJEtDChleG4iJVk9a1xyvH2gmkn9kA9mwCrAaXXc2zeZJc8/+YqQbaJeL
pq743Z2+mrlewFR6IemfNFFaYM9/rlAEIz8gr7zvkOxU5jlhlgUcXQolPv3RL+NeELOC04D5Zr8/
LXQ5+0G7W7BHLdz45WdZqAhJ7RQb2xQQraxRWECnMOSY1whvYKyQWOuI1MS6WfKCUW74GhCj/b9a
NLaBx8fXJGMqeiFi5Nz0Tak5UGXmxFETBioMGpia49kP3hZGJfgM3V+X6xM/3AASjlZrhhLfAf9d
XttIbeL112+Z2ihcBlhEyOHsrgsrHGM5G7WfZRs9FahKJ2yI3sXGtQQnK392QHYmbfDB+yTztS2E
EKlCfao3q7fktR1FnRYblJbF2EJ0XHWyMqxqDjtMr+JZOIE1JC9+je66NVbX6kZuwvjq/s/3K76w
kgMuvZ8bDxzsxlmtpLPL3xAnqjjePQadIUFdV0n3earbh/pMmg2Ay1SOgjOc8FlPrnadKfE6mrN5
JSdtw3wX12tJESbkfL0vrsOkohk3N4GTOL8tF0cJ110XAwp3pdZ/o3loqbshBdvUAmGv3DzP04sy
9x+XBGf4rlZ2TZx4WK5VIU7+FVvyEDgYTdXTQfgue5QpTywdHBDwnXWfDVkitRU8CunSuKzP3JPO
Wg2GDlemBfJmOSQnAn6G9M99lksirkyZc6SWN+RcLg080ULxTOnzFTj/oQz8nJCqKGAxBWKXtukH
VKB5RyPnRDvDdYtN/QYFzK3WscC4vH9JT0WZCla6kQMK3R+IcejtD219+EhSE5/Hf/Lk5RC9CDpq
8ijFP3QJSGCvrSnIbeHtnsAnj8RR8QBnP/z8fhw/h7NADglosleScmd3qqzM3KVYd30SzdE1MeCb
A0V8itF7ZR7adJ406ah8AmK9uPn9cwh99Ewhad96+VLi2xS0qRjG3OlZxHT64Q1HfWk2v7Xr/tlx
66Y85qJMMVBpk3v6nXgKiZxURp2KYy4RycdsyRFcim2D/izycxXkrF4Qzv9xwfGsFk/HI4w6e853
n3HijOOkH5K6r60rwY5kHWmP8QIsDKRPZyiCmA6w+m97kV6rRkkFlm0sJQeXtgOZVNXnyASpHY+O
r3UPdw6BJCDKTOUIJqDH955cqmOJGXqRB9Sg5g899EcQB59LYaOi0N/MNJXySdYHrpgN1aoJFONi
10Ogx05mvZNoq6eAIfPZUJuKxYMPvskdBOWgruZYDqGar6673pHuJ+LGlssJGFSPIWPr1z3nrtPq
q2worMOc9R4vn8sDZqxpVjYUZ2CldO77Uwl/ScmFIGvJ72NcPXjXtiizGn7osCCzjwVYVdQobh/Z
8RXXuo89EVaXtNy/+mGyCACMYw3UIVSpKcUBHOUyprQZKUcJqJ5C/hfni+m9aMUXo94EaYjFCoan
Wa2Z0cbAQKfF/gXEjuplXTKA923esEUxPu31zIT+vKVPflgFYEZOcs4Ed2dN0HkTNtPxIAIKIIMj
u0d0GEUvTVywW7kP0bZfhL22eGPDfJ0uwSbRddxtvI4A5KFAGxWf65iokPEH7lmxRU8FLsfndVVJ
BDmVh0GBJGxe9wt4DHelojYXAUaIBADxh8yseee4gJjImKHMpCv1ihhh9pQyxFbuOCmDM7BrfE0U
JLWHbMghT1ClehZG1NYOjnKUqXtvLcVshfcr4jBdEsDgJgjjc8aglgIQYs2V+syQm43xePGABdjN
JKcuy7RTOxMZEcA4QQJQIz5qLqzlE7Ig8mal+aUEbKy7NORZ/3m2L2I5hwZKpkWfbMbZuhEiZo1o
QEWGWl6ApBsSPKgP1QCLLVq3WJ57fV/90ZIFchRVxrx9HcR8fMlSkvr1QDkgDRsIGB8ZC70rqxwy
bGkyfzO+tU0LTiJEFau2Awx9DGK58OdlAv/q6IbdCjKP8A21QUgC3piu89pS6NAMZunMNSZKPxnJ
ueFbLIFUzJiDKZ9J/QJ7+XgWcedi+dpwORW08hsx8ReLMetb/uhYmJlupioqA3Rp3DYi/7unmQrF
+AhHD8qb8bBXpTTRdch5n3RLhvarv2N7FWQVpPo23yNf50GovS8GQ9GIs5EbDUr7KFNf1cfDjDiN
6mALAdMx8L1lmHVyS2kDaUj2KNxB0ZlogSR4KEPI/ZLSEs5GlckAaWiH4Wx+s2BgqRR66B9Mf2+A
a2RZdkVbpulfwkbT67r+VOIAJh42jYP/dKfGKN6nkOX4FT600XeloKWyLTLI4Tg9Ts11zf6izVVu
348krp3Ppzk011MQtHPyTmssuo8e5qOPPZMc53uhn9GVH+P/+nM12HqpjhxZjk7G9RHqUOz3luWz
oClB0O0pN2I5ly8rkyVF5fxl8aV+GtdnhI8m3k5LaXOQCuZvxFAiNdv2y46Vf+hPg/k1UzVaTxXA
5J/ROL9B4mBfkvgkBn9j3c+r0WxE45ZImOridAmWi/6ScLEvgzIK+PvEXEP0XX6Pmk1n8cnh8g/9
C6avS0DFPkyrhtiISAIzK1BV6/mIs8S5LgmTyc4U9CykgA0lO/v4HCgkwTTu4dqQ6MgvPkhKjrXy
PhDXrx5aYRV+tQSQMmKgNEfqM1lfrcSOYz40DVhQkuGqbgVBqRmMlBaNYCryBF2sXOnxmrAfi74n
Qd8x7Fd7GBcxBb23vrUvJX8btC10O0+a5ubPY1X7msn93E5VkclQ9sQ9F9YmvNDcbRUVQDPhjJR4
wuP42amoa9qFT5oRBPUjSH/TBAeACjPoFn98eYkgJbsIJGOBblDWHlfArbYfNE4ZS0wfJSvCzbOP
cVgpE+ruxy1U5DZHBNDAFjWpWmMrWaD6NH621/7NU3gtL2AO9Fa0Yln04ru32B9er6Y8f0g4lPPX
CveU3EWCrLezhXPK5/nAC5HFHnm9cDIsLuDCR6pmDHB03QWFvaiIRwXLBuaLV3p5NwXdZcuNFWgw
3EdLwkJQO47jvVEQtSattomUz6UdjROQ2JLYm7YFBVQFKf0gr7ci1qrMbUR4ijMkjfdgmD/+DnhH
+rAMibkoKNYmat3Gdg2D7U9nxvTI3xV5frMPEDJD1OkjWfm1mZf1aP8eBeupGdphZxdLI02JwOOO
6aXJTHYjEDTSW7kLCLjzo//YbgKAEh4iuUKhyxW/ANSCaOFJnyJKoNXgOPo5kUusaUuHdhStC1kg
eojCKBno51rrcgJ0YsjoK7ehg7Hed38xZKtQPnttBnNa+abxbq5dsp1sWUH5lP3B30KOHEdE3Ama
MC6zI9KrJQ0j0h7U2GfDjzHIrokr7RjKezXwuHR/ROHgJTdSM+ACejbNCR46t6YZcquzBVbUAPgV
zo8FX9rzxbT5d8DkDN3bDFJaG87CEuYP21972B0TMfbf0e5PMk8MHnRUZqOve7ZifRBVVa2x/jGk
0WIdColgF19X0LcrwCds9HkxueGURnIA323aQli/if9jCPI455pyBEpeOYZ4JN0e3jieVfYxYfZX
if2YyfvlYF+Pq6bt8wTjVvcljlwZp9X2lw5Bz3x9OXPUj9WlmLQ5aMj/DvZymC/czmd9Zv+Uh0mP
AI1eYuzo6XGt5tsiULW4zcYc2AY6uCzl4VylAeIJhoO3p7xU34pJuYOQmNyULt6fSOFy76m5I7Ff
QigH0e/IbxOoCwXSGXEuYqyImb5ME7LhGkX4wbpfUZi4IBgeKOo7gn38W7vxp5jBwHYb6ItsTP/h
z05TUe82jUNquwJ5/LT4UuPbscaBwv9f16VbvKBn90nyZBDOeyonnEQ0kmVqPn3o5hLBAyocFbra
JNOZAn2NwhjgSoDBBzfHQIrzU3s9AiTgd+ql4bqWR/cJisCvI7opZm6RrcASXkbaaVJ+lkdzAIEb
kwHcZcdnbh+OIC0rh4RkGth3z0fnuL63XBiLVHYgbA1iYLCbPsYv+O5kIi5NlyTYr9/h8DlvARGX
bZ8r4CoosBo8hFhL+YFkz4CziJcZnjNXZ/0VGkwlym+3yMG/zEpXTqEq0Jlf44nRip5JlkMMVJy9
mXgM4FMmVhnStPGQat1nVyxIP4WVWWHw4PfLWqmZOD+cV5nxA0n/tXb9Cbj7YDtja8zgbVmi1Ncu
/RCDbgQ0bhOtNB/6wWDVqlw9jMxLTjyfdEUr/q6lVoraFmvCUOqPelEyXdvqOz6Dj1aTSqhCbYZK
l1YZTJZd36DeqrMXVwpYKVnApHzPKCLcm9VYnVM4tLJW4C5YmHukWDPKKkFZrmDg7VwATr5bu5xM
ZLVEru0TceH018LPoa23NlMgCNVDn1u/M+UFGERNVIysrTuN9kGPH6VVTKQOb2b3CHp/60+MGlvJ
odqmqyMaNstrR5GKM0DLRoZh54YPDiB0yIO8xejANxdkCIzr59JZp8I4wFZ7Q9HAN1FTGBS5lmtC
s7Z2oK8rWy7WYlNyuvFeFMPDkzpZ979d+VFwAo4/HA1Wy8C0V0hkCIJqLufUwwhI3AZVALbPOaIz
e650/jwsuyN65caKxaZAP3c+OB7IUDIEvDwLL1W8Eh+b4Y772cs3sbekursXDXO78b9hdpLSr/Nu
2abCG0D2UmTbBm/XsXqWLMga5dz2Q+35hQuyMd8gL5UBNYr5FfN55nSWuW7Q7emxS1WMFrk8fGND
qze8rhiCtLeoSMdMnDrhIzBPXLWeYsIOLzanlNIRWcfPsxHbEDpEXcatnKZU3cZcskZvpG7pK//P
xoQbLw8pwGi0SnbdvMtWS2qedxIyYcDeWFN5V7lDPuwDPlwXYmrCa76RCLdchIqdw2qsWhVFQJOc
f7ykN46UxBxVZ0qItx0ApHTdnVVlrq/lYTl/gqX8eeNCG/7Sftny5H1f50kQFGdmJ7O1PbeuoyqP
ZocvoJPnvv7jcptJ5kYj04zvqcHLMFgyXGUSZrCghuargRZu/vMFZSgUXjh5PMgWVs+Hv18A15Lk
d9/MJxeL/m2OxZmCPNKNw/eRKLYfIJy/Qub2UM1KS6FdYCSZLUxFaDBTi/g7O+saxOOCps2ii9df
zJfMjR4bZ1Y33/3vNf3BOfyLu95+FB9xnXIyokeqIwTmkxBUB3cElWvuKnpA1reIqf2wLHUfuZEO
I1/dfAxL8e2Uli7A2FnUO9juZXV2B0wJtr5LliPa1D8iLD6t8eZ3PS72jnpN4HX7FafT+a/WE2C+
2pzGHTeenjVSCR1YjeyA7cs2gjDyhknjGDUp3Lst+BQrVy+E9ROglYXNjLFjWuymwRnnJbTHI/UU
DYUaIKbHu9fEVOH8P6wyGQE7nZoWukCHhFSTJ+d8WV8+ry1TNz8MJr4MsDoxXXZJZaLCq73Y8v/1
voNU5YNnGhM/WchnXe0yJ5zK9Oz3u/d7ZCljA9jKBamhz0xXBYQD3tEhWe5P7Tp3j1k88c5XgsIC
5tGqQAv3/ORcnxTIX82ffQFwUDPx1CjxL/uXntMG3njuU5KWVKaGzSIkIh5P9+tNNGx12A3X4DNQ
btXV8GVfMT5wSVIaZUDcw8+Nn9+Lxi6uwIUx8UYtweYhEpFd936DX8ZVqIU2VKSlIiAOvuZye/HO
Y++vVhyKfm4oYCGfhhoJWrDGIzYR6RxjG8nklz9oqbcBjnMWcayJP9TCtG78kUI+RTvA8cYCfgSG
qzuuR+4mAFvVu91/XYN5enrswAExH1bveU+TwQQIdD3FEPXfJE2ycPmmHnyVvcjToEDmNhyDAuT9
R471Gqcfw+BBTFkMlZlIoJHQ06cjM/W9Kyy6J0vOYBFQYUkHRwL9zKfyA6kKJFkBB/S3xcj//Zi/
qp/X/rq3WdI3r1mYT0X8uIidv5b5KXXA4hwy41obnSmfglyuU07S/7dMe1t/1RY1Ab20XGW/mGFQ
mcNxJ8237lsJfqCUKEvOJN4lI4UDXlc/qUg0pWxPYpV5AW1Xu50wR61EnuJvxe/tPUji+iCpA0Su
0sRY3Gz6nceZzp3aM56UHuPb4njpzdOvuTL8LPVWsL0NAm2WZLOJBCltvC1AEQ36FkhDVa0YDBvN
O/US/f4ppAYhtnPozNU2G46VoyZc4vDd4uXw4oi16zzYFOCLbGNYLAxx8tDxltO7U9c48/k+Birw
5dLZauRz1Yc9hCWUHzkzNENUTrLaKZSZaWlbl8hKj7HJ5MEr2iXgAP/+L/P/T5y0Ht18TYNryGjL
bg8kgOEhcByqmGy7gId9sbqk6glSi+hwQ3TUIP+4h3tq6Cf7w+VQa9BaDimnPof6ijfaTu0WT1jM
2I8ujbj0qJpsEmhVxKbFZ2Jke5x9BMDTGFRkD85U+CH6pvicdErtESvLmIcS+wdD8hpP0FCAcbok
llaNqHKvq862lKadVyNRcJupQlA0b42lauBqFVr6V+FiPojbnCqHxmasf5ib9wp9/hrZSsIKMgFz
Y5RaK5q/YxdmiLGeym7XmCC24IRm1+OGxROUuVmAWOZ1RMzwhHgQEL2O1WrOnpNLUaS3RHii0Cww
pfwMtoXhWA0ejXGHU2/PtsISRYNkUzWMFrNhvmzB2M1phRN/Ly1pXRWLAcLANeKq73VZ0m6PlWjW
47sra/NLKbvzCU+WyeOnOf0oe+qIf/eS12cgN18vJsUfTsdoM1VuRtaSh+VMMS6RrBUIsLFf2n+F
8bHjgDRE6bV2qWt0ZGqpk4Us1tWk5D0BuH/3L6BxjgTi5JBKg6e+1oDKeTE3KOTtyIWskjofzFfy
pKDfe2F+hEDrsKfek2JAn0TVDxFpD4atKE4lTV5yzkSzDfBCdaCN1Fo75ufTHMP7+MKruv/Q+xXY
I83wbCHH7mYMnPXYe5g4w6KCk8nermQtUyDADTj4jsxRGEk2j29Quudr3HhDHhbQgECvKtskPgAM
/bgOtgJvWHP83QqQP8hw4SB0nCoQxxKoOpjEPWJA6WShtBHWK+ABc3UBFoTBxfF8WVYcreMQyqJb
g3XdCHsmfeopjncDiuWs2DhMkx4ZN55NReDi3lb0VuptU+XxKwQatE1pvxiA0VQiincqk8L32d8+
orbzHOoVUBSWAfJMFam9SfzArNqDWGBBaK8uWAIon/FfX31/EkDfYxgKIi3Fr5PNCwoGHpDbDFMw
AGaY7+7mD7d0UeKvjZRDCBUI0BLHm14qJuAyucvXCz3i504KgvORoopDc87umJfisPxSueDTYqM8
dC26E8TnPc91FVG5ehrULYZI0E8SSNMuq4CQQeOs8p3LtMYlvJjZRDOEY6QNmbgYXQ8mSY7loxPt
+YUI2hvKwV0ZtaJA85gLjqN/pNlN5aCo/LRJUUWmL7/mOxM8VAOqN34BTf6DrPRxBUcnQWU6qS52
qxP8Mkj2fHLzeGpW7B9aRa1hKEHcSmEjODxlKbqUR+/6msWYURo4YCT0cULXWUnVhyHeHXoPe5k+
1sSx09nh3Ie1LvKdOpp5PHdPHLVblnQSxPCS1M6KCCQnGVfmXvf388qCZzS1Wd02b3hkEy3U+hYR
x0YbDhuN9xfzpZpRsqwhTZKDTNBB3xt9iK/MB0fyhk4rqpi/6l2c0UrCVrzQLCaz+wGmyfyCZpPD
43x8erz+Z2PhikCzBT5cxc3/JCUwaM/GIzcCIRH3dphig44Z8OWK+y4+89zG7oXe9ttVOJT/9knu
1Rh3RyiO9p30Q4rCU5lH+TKK4SX7aB80CufwzxrWP4b8PpdpmoQu2VFcAtyowbisapaCqw931UT9
itUF+cqjga9g0Fx5R8rM8HCygu2xQuJLSgF14GvIucaAfyh4cYxi/SpHy+lrr9+iyMT26TXFkOiT
KcVbQstkztqyVNwf10rA5X+ydd6nb3hkP3Ud6xba7jE519EcBcw3tYUxaJaOT8KUqlP+5d3ltJZM
O5eWnhfc4jX0+pO74eMudFjICgZhfcVtKNdJAsuT9NBoOvH4MejrCWm8HbcKHBpspliKvR+EMSvi
YpkLIp9/YcuwMNXiBcLqPg/YzQGA6ET6pBN0bmmSXJiBBhpkXYrXkewtl3xg27KGTyDyuXyBrHhd
6eekvzCN5fCs4YkQEOlzmi2vDALWGdDnJW71yMwW9ZE4sCbKZr3s6D52/YR2gf6DkRqGmUYKJJr9
1o1Epgcu4vUqbNrLap21J3AgZHt/9Efn398mvsrdMLPc7M/yu9N4ShOAa3xTCXU2Fl+aq8LzWgLg
bkhaz8kKPuFNZmL9DSncvnm201FWjsI1a7GCIDMaCSloPxFbtAPnucxeULLPW7E0Wcjyk1SLLcyG
yDTVXgGb2+WX4Cg0vt4vqLLSNmWQXvmAbNe6/vBk6kpo9ayrnszdNfzGgr/GUFklnjshMMudaSV2
NbTB8fcDGVjWzpJemjh27LusDJZD4vBq4Ai1twgr0eX1ADo8XCLN6RS1mWKmrMxAYYHVdYzwny17
SwGgpb5yCXT+9q7SwFTfCcVIDg+POQ+HaXI3tirY2la82mXntmqxHnDY/20ccn3ZrElZ92t2aG3j
6V3y9rGqGEPwCmCl4S2RbRUl8BjYiIDRm3De0/mJ3pWcKQZVCl0yTW2g08+naOQKLIczQunWSkxR
lZ9FrPwJrBeaAyyDmmB/Fzjqp1qdw0i0n+aCMmmnETrld+6SjtUGbGgL/bhyL+r6sNcJskiwrZ8D
wsVgi7ikxhjxFSrgE1CbDe9wBKAdLFwTnICcjmR3D9vd6lCSqUO+ObdQICNWOe/kIvwYWx3Q0+QB
GV5aFAd2HxBSNGESHN+n2NOqVNEm8BtsNCBHQiPdt4GWGmQ/EyVhe9JujiOnMDskosQ8STkAKfud
XYtXTXa+eG7ffMAgpkrtA0DVp1dVxkHh2crKvTUTsWqvahCgrOhO96DWfPoPR/CSFXNZw/smFK4h
ByAPJMamXXM7qElbWWozz9fKSjuIa0nd/amkz9HzUkikIfCneZQsZKHLZk9xotbU6lwDwsn8fGRx
42lwIr+baAXenwUhuYCcpX+OvzzU0hnSlgo6jSvxvJcFz/TOQo0vELE/ddNtWsgkrY50fIEWGbId
Wpzj47hCGVKs+MYPlsMtXR3iGrFJlqG1m6LcFzb3xsefgpdfAunTFJCtJl2Iub/cqYOU1zHkcX3Y
R8eeFuXEykGb3s9CSnZGkNSF7OBsP2Z9hcbrSEOP0c6EKLjirpdQDLRRsbHtj+4iRvnhIOAEO0cF
Dyc838SC8TpaWNMN8EF9t7DhyzzjHQvPJ+oFYOqUrZIxiiy30YsdYb8KbanDArTC71fpWidQSz+k
pK+hLrfsh4/aUwcGMdJC2ppQP7qySSf1f5gKc1Nmw42rwVnzF6sl+1Fjgl5odGAlOob3Vdbw0Fbl
/SGzHyUBNceh0ifCsKLznSH++LLq3EO/NRJOQYDNb7bPN4NmMVQCnK4CNtklDUGfCnjKtNJjT6Cf
afpABsO/gVPLXVu3jJY6Vj/RMbTtJZ0924FDwv860ROlcO1ro1ozV6NY+USkaof00BlteKAjmJX7
zGfdBFM5TWzR6oXGcMEpKENrtkPYhX2a+A3urOH9Z2MvG4zhD1tLQrdEt9zp8fZ+VhABrlT/Oh4j
AMWJu1kW5pdSdt9gYOyIiksE0NBugRF7hSXjM2HpINYzfHUWwU5PhAd6xHalI50FCyr9cMZfJaky
2In+ak0NuGFrpQ0jnTxxCypPA5ii1GNUruxoW2dvRWHKVvDadZ49hd2H5v1mlbeXa4S0AiBk/fz9
sGZuLn/9ascdna6qL463Sa3346PeYW6hYdgFQsNJcoFT9INCJXt3w5Wn48hFTPWDEvkLPx7x6b5A
0CrP9PI1WK1Mpgev6Edv4S8XZLj8h+LIOd/j68Nry0xHr92caUk4GF6VVvzHTgeJI1XizYwHA7hT
NLKBAAvZmV9rBg9ExswUvDHlwKf2sox3uw/QGrRE8WCXNrJ9qcV/SQrztEZD/bF4XDj5gVzpchMh
DClqGw2Q3OtDPpWXmQAJ7S0/8YleFokckVERsEh8oFJwXWyRcWp6WlVuTS/BeKhH7Wv8XUKvp5i1
vUB+8cOO3UwWIsG1ZgnCYyQJuliDbqbK8C5cDknBoz/IfH/alUSsm7emtpRFpD6VT099rEjtNF5m
3AOBgQ+n3KizP5XCSzPow4A6cfDXokpBb/YKgW5QoMWgm+M2BrhMItGB/CXj13tq141CMaqZjn1o
qPpuFv5frEqYbnKqHF13GQPZeWrpTekON/xUUcwHFIVKhicgvk1GjA7sQWNIynY+TfrF1MGQ6dlr
cy8JNa5WrGD0bHe0hffNALoMDnIzpmRZ1RTgYaCCEWps6XdJQLbjiMyn9XlTLTO9Xeyh6G+LvcwO
vAKiBVm2WKxFRJRpNkqvLrj5esKd3f59yqyNAPnnJGVxc8SiF7q2OG/yevj6/dpsSXgAwrMzhh0c
d7JdvfhkLDm6JW6s79wFlsOAam8CW0QQjXq0nRa4YWXZOiDWxS8vUa++1/avWGePLxszhj9PUvor
sfGY0nip2S2o5NE7M6SM/CUKfeOd96ndhMt+Q95go33lZi8PokMEoKw6dBfUiTfW/HP83LPgT1YQ
vV+nsObz6QsJqIfbey+8BEPzKUHk3g3doHpRzoPHqki5HgJJmCxFd+lVWd4cw85MRVbr7aNfAfDX
iSE9Zpal7XwIIVrVBnDGeHRt2Tq6gAdPbCzpD+vlFpFtXpzp3HJLjpko4HCla9fZhQ2G+gQH7A7U
naM5Oa1O3Gfu7JnnndcTOgoJHXl4dJ/gPMOyJMTtnL14ehpVCfByanB3VfSeafU1FtNnsIYJUORc
AtIZVo8MYIQsa4092UHjnTyCbNPLxGsGCmi3Zibc4g9aXjKEC/rsZ9zLyITpEWbFGaE1Cvh5J5El
1qXR3l7n0SaswCKZcATZ+qX4XXYxhLRlZzMpV1zW3PJEQe8Unv7l4gXl2xNM14NKxLp5vE5IGaHA
PZC+hu1xEiOV2v9ELIplvY3o33Feqn5zfnPKZydjKnXlJNWohmeHf82hA3+LAM8NoLC3OEkAJuqF
0z/Jc/B5P26FBVGOF8qfCmJMwwhvl6SWMIdlyXD190l8VpOM87M4rhsPTChRDhHhPwkwKqJqHl/a
Dcg8ECF+4EXFB3RXDe3C8UfuY78xgLy3x9iZbOYRtOOyaLsRUScpdQoIe6CddTAWF/sZ2/M1Ehv3
+oaSEY3T08AKz6CO80XNL6gRtaNggfHf33tZpE/4wngL8aeaNNsTL1tFSBH8MKZotiVuBlKVukaK
Ow/WPneX0eI3tDmmfTwrYFLq9R8S/YT+jYIM71NEYmPCfkTEDLo5ohudbOVpQzR0N6/CKuBqpugd
m7CqWc8yOyKFuFNA6oRomvI3d5DzlBFIuV7fYyfSTBx87udQf5WkU5pGX+M88j+tkLOadlq5MArU
lFESDP/DHS6TtLNpaMjn9L/1ovzBEpz3iMw1bQEecEIXRNcbwi/vkLbDwlG7dxTaUTm7Ds8vwwQy
K/08/a2HQFUweBQbk20hoklbEQ6Ff3o5uGddzPkLL5ZggGXiWheasl3Ad9IGwnHeT+4Wu73n8dzC
vYPNIGXdmjrMTRL21NDMrieu0raLvu67VwVC1OITcMls1r3+Rmy1d67RoxgLVflHznCVOTLjldi7
sDC+IoCCLv+iKBKK/ZQfYzG3bjqCbVd0/op2gmELRJFSkG9fX1zNHH/fxTSjKlgDTjGkVy2nPPOs
fTRMoLhRe282Xp7o6mjHcejqUHpm4Gg3vWbvI3qX41PF2TVZk1aj4OyWncKuwKdcXAf4+gPBce/b
jaNKRboIus/43zVUfxwCqFhWvVz0ksngMb77JPylxRU0qB5nKP9U6nkiBWF4HuGXedxLHPZ/X9QV
OSW3MtWmzwez/QXlJtWPqdKjcuOZ1aqk94UsXckS0VNqTvuVI/r6W4KVNtU81tfskvQfWcydR4aH
9js2cnlrc0HS9vYKTcuPKk9hCfMYrdLnjKn6aBfrKvLDdoXIK/eqO3NqnhKade6PlVOR0ZoicMfP
zspyXAS5ZD31eb9lmUTIfwTHtgtE9GsQNBD1ijAqQ3XRZORqcuTkRttz9lawDeQw89uIu6CbCZvL
qFrpvamtDSrcLpMLBs6XWUN3rBIReUY8nXbNtwgUTRJkWn5W6tbnFoPqrnU34+QSp/xXZczfQ198
EWLwN9BxDlGGvnZtS6WYdFcTJTVNFotVGKy6kKXvjragnCZdNtP82YAT0UXzpi3h2Kb7m1OcXv0g
e881E9qzfzfViLKiTRhe+IZ6k1HFRFZVPOXH3oPlrlmYvLp2yTobh00to5idD2R+z1vME4pGszOm
aGYAt/ykK+YDG9uEqfgquEIGtLGV21ZsRpDblUr82nfQ/Pqb9xcA6iPnVPxMCv3g5WF7Oz61AQxX
4zo/wLJLYSf3Mo5Nf4sqLMVyyqnIyFWWIle0wyrUGuIlm7QYyioDuDAnMZwobJOJe3oEq+8SbGdA
Q3DYT/EHfCAhMmsceo/sr8Cy69FuGA5fa0UArMvSf8S2uwIA/xZETCq3VfncTm9s4IeGM7atBko/
o3tAkWmnga3EPOQF1+cjncNOj5o0eLkgWM5IkcIlNzTejddjcbZeQOWOd8ATt7aA3M6GwPLf6UOe
MjintGxvu5sNj//jqmWIzjFlWcQgGJPHxxH+E/e+aZksLEieob3JKvGzCmjO3MG6SP0JRRCQpj0w
qSba+CMjlJZdl1COXuc91i41/obf+bUmxGYfnX39sV882jWnp8yVEomeTve4W2JSIscMP6KcfQ1v
SQJf9dWyUyPqlDLZvj8EHZxLIZ0dGFNIIJm1EXfNJ69KyaRzi1nX/t3dsKC1isZfqghpxcOQbtS3
7vWPso9e1FshfBJ40tVDzRug/Qx9dHgL8/v1vE2mem+Dq/IulV1I/LwVqRURZHo5nYjQgCmASJpn
2SHFMMdRMRts4JBl8RFiSS6FLYYN6bugayWdEXfBwTGZokTKvDpJUAfksSWRG4xu/PydENZ4KdbC
dKnbfiZBa5XgkXFtuRCd+kqh2zmuF6ilCKXLBpy6Lem1JIv1eUgxvrnKhqT/9wTLIbxDcHtG1j+t
G1SHUj/rncUbJosTI1ihmL7VlzeGWy0W/oC/QcJqXCfVu7mvVpBICdAqJD/fTUMF9SfBBh+6U0gu
UmkFIzY2IOzU+w3zpplWQ2Ktv4s6An7VaPVhD1+49WKrLBm9GHpSPopuhiIDoIE5/n7wGHqHiNjs
oDdQ72P0RSBB4d95qhCQYyNfAbfuXsJwmCtaeDbgMpmfUCvg56jtUuWLkShFn5aU7pipyFSbTba4
eeU4NWeTuoVgCJnnS/UgaB860tOomwRNSjXIUh982jj+nadALD8GIANvVE7/Gp0IqNtESBGRGf4q
DUTdgMNdan63cgJRwZ3siJQAjC/CQ8oCeZacljZGObFVsZbQDtcG/RWWmubiGPM+N9drfMVWrxJg
nR9/kDse0q5kh4v23WpRsGgOdvhpYqdrdUB2OuW7Zue4AuFNgsyMQ4kNEfK8HfI+bSy1SOYCNfjB
mxzWGr1xrVBVumNl/pVuoneYEtGov02DnW9Knc+3D6xxO7lWWtoZQNPohgZ3OdLqOIU3A+5Dvvs8
j7/nEuetoPPUFWWyATjT9yjvUL1+iA1TCfj6GoBZv57/VxpT9TeFBe3vG6VmktCPpw3vHA8wf9Ct
pPhjxW/UgVsvn90xPbaMpKcm7z9LOsFsJ1TT9OIioXaTACcOt3LI97vmK8bmft8YF+p+Xx0hchnA
M3pq9fK/3whuZ9CzZlCEvL/nsrMYU9RYLo2pN2RqXw4vGbT0QadO8omnSxMow9pCZequH7J4XoAZ
ZUTJJlylbdqQnpwyRinSr521TPL7IyJX23s90KgFeD2IIbdEfsOPL/1m0gvbpXNrvSTCzyTfwmt3
GZIbFGXndlQjQKVFXQamx3UYTTljQ5Gpy1VDLiUtouxbMleDMe/OGNCDLMf9fgoPr0myC+PT7Uye
x0CAyfNAe+t1HboVYqPTOmgVJ9J0eODNYhsDabzL89RQTzSepY/5CyOlQbeenpNND+LRNoNRrnPD
usa2asKfwGsQS2vJ+nDAeDhE+Wp4QsCyEHxOZN0Xj+zvTw3P0l1Y1vCYmry+uw/Pk1vMwzfFoL3q
Oqpbl2s3VbA6fNolJsPufvQIPimgbx8g8FBWn/Of9QvXuKZlFpTBuRKfXMnGS94dCqf+P+GeYrHS
1+StGP0YnR4nnkRS/3CayMTzymMcAyYgPNamhmHah5utOepjemxBEd9Fahqt1ko8I05CG1D8LcEj
28DH/fI4CmF4aMi9StvW4LI3Nb87ynyfXOXVoj40dkyVy6wyumuUEn/fv4hfj0xNQAu3s3M6vD70
mTp+Hj3Y0z+1pZeGUz6NCfrQYKRQNQ29Z0guPA5F9SianO3x6Qiad8wb9LqVEztAU440wQr5y4UJ
p2+pSZJoli/rxjC69lP13NlWpwTCr88weZUC4PMRYNgAdtaihcHBmh7Gq1IcghX259ankjmoGDgU
Ck7h+DQezjHIPw2g54xuzRZcFzMQ+9y7EVTdlqVIC6IqWnYhyITkqJ91G5wzEwpPgHhZrGDJalfc
vDQTMo09Ne7eLVoUYLO6GyatJcxj0kCPgp/t3R/PhqQ+Xizr95mhABjEiX8JRP8QvyAIEPmAIm8N
eXFjh0rIVHM40a4XuPKyDBWyEgkn8kiep15J0grW4IyO7JyL3liRxtllGFgluOgbJnY7ni8DGzPh
SgwrnfDjP+a1TuujPeJhbyUhMk8UO3QEfz5SX0zXCm0TpI1j5WP0He0rI9jbVFE5cjNIMmKAZFU7
3Vns+K+PvGwW7Cl7tg72j+Fo5xVy0fia5fBFkIh+iRcaE11Z3yIOhAav/Bs5yVKjR8Al4q+l+JEe
16sI5Czyg/MTpG54L0xLYEQ99ppG4EOv+dHCm28TU6/E7A36NTXrW984dEFfLTce50ARDEJDcMyS
JczzDpJHLTR88lDUPX24jAqLWykbBkwP+2IUwWcl7JqKhrOD71tYs4EZaeRgoe9vV7jz5znIwTSx
elJL+nC52I6bkeHnGfuv4lMDDjx55DoUm34ogfRlUSS3tJwPfNbDrnTQrRmYavGWLhhIb8nHqC39
q0y9diY1RpBasMv6qAodY1KBM/nDoHg2KvpuEuWdDxR/d8+acTjyNBuVZWiCr9s853casSMNWnKL
kDmlwIDfRpnZMr7hkMqU8VUZ5qjdxl3FUbRLjnepr8gy1vZp25LsUC7yWK/KIjSD/Zd6AAh0BRMq
fF5hQ/K1oO3DFHYOkSqjq29e5PUo5OZr7nydyqh0vnPLjZ8USGSMS6vWAAiCaIUYxWwRA9wliJoa
qrmFTls++COB3hHs3r6+bxy21eJkDwAS5olNhXEKEAnMQNFtRBo0xkANJhsUnux+PN72X72z3qcI
Rhup0DBwhhzwtf0rcszZ/1B62NZeC/yMgyFLI4rI3Clydj+U2kQsF7tZExT8BKK0iXLVakmyRklq
oH3cDLhrmDOORsG1WqR3TPrsJKDKJalUiPMF18JpJIjoVZSAcbs1FFhqI3HVDeR5Qwc55TLvB0F+
rClJLu1NTXaJcONLh5VJX+jhOoHpCfoOkvoyLUn5s2lUR0BovrtvezLcEeGfFV6GmeTsrUX2YIac
kiNuu4G/WAlhvKYmyq9UGlaXDCX1sNiK3zvHchxpe5Ba70Js0zcoBLvD7LAd+HGeUxbPH+pJeY7E
motGQNvl9JJh+YaDxrFXIyd32+GAlOFFHsKwRNGHv+bGm+VHygdZ8hGws2gXutQok0s/IkWWbbcf
3Rcc1g/tuSVkt4kP/yLdoxFYOrfOazK0PFYFVF2vxfl0lsXv5NHyGoNietLjhkgi9Iw9jHfBLkM/
jUVDZXi2Kd6SRdShj81c46A2jjnTFnqdc7Zn/eBVq2ShvEUm1Dsl3IfocH/ycrJZ8/7z4O8iDjtV
/QK/jMQ7BxfvCZ00TUFabIF6R5RYLomXl4jPbBcyHLAFNtOEMK0/ohwdgRBnM4Jz5FkysC3qLk/d
lszzU0h23OswlyaekV33aFWD+S4n6skh2U/H2HwIhqs521vHyrLwre+Z6HkfbEgdi9/mBH4CnKq0
aMuusVkLpRy82QhfxdGpLVqVhhe5MHpD6NZy765ilc9JRpy0iZ9UzMmmzFAWy+067/gptlN5VR8x
oaEQTm4PpUKppe5Yl1w1p2cz+I2jbyGUVza11g0bLny8ucZCaVIUBtPWWTWG0Z00rCvaVhFoyVTD
wmSKxdjhGWeuLdzB37Ge1CPSYR9FOSN3sEBeGYj423CY8kC2DnIw02J6EvOG/6r0euM1gZv27rdk
HUcYcsHkFgH9UYt2SWtAiAQq0bkYUr0uK4XTP/rYUhMTAjZz5K4oigZJL2SWzRRfgD4+mvIEV/ew
FjJwFM3+Z9g2Vjd8IDmpdMMcNWU/Uewcf0b2HDyLoNzFw9mTCQc+jA7RpzGuCTTpY4u39/ygBWFJ
xknCD1E32U/v/fpACaCBS2qygDl58kl1DoQkrhuDj7EsOKqcGImGYdpMEw8kTfsq2PaJrB2l9v3E
nfgy/reMwrUudM24fumfZv/T+DCOeA/+bjOFiXUapSTJn9b6eRk6E2Ahjtqk2Dp+9Y0LJDK74ht8
gnbr2YtRNBfFXGXaJk/UM/4rlIlD6v6edi2qln2ukjIskHQT8bTZmzqMifGe5+1Ev3F8suFwUxJZ
qwe7462k9wiNYTpbN023/AfE4rnskUuAu+AivA3OPy6Ey20MQr/NqHUf9euMXNYtWePZy0QWHRXM
py4c3sXBEtXVfKFhmRFY0z8P/KyePGYVav+/RciCJuWLbB8FE5mLN4zh/HgC4kiR6IRU/KrUdSSh
K9S+MwovKHzXnoQ4d+a8f6P21S3XRty714+/Hh8Af3//kDIruSvP8mSFQTSKI1OsAqmPB3yeN1OU
G0SpnyeJURmGEQqWk3sfDGwooCKz9gLXyxsnU1lGunKwF+9zowyA/ER33eip3g6mFeGlOoeuAXNM
SBDWKfvmvoe1obZfqCAMWH9EGz1eX9P4uQCaZf8NOR7zKL6LINUzYjnDR95He8quymz27npJ/Otm
e73YnSIwrJs3DpgJqQPSEEx2LpkgIuzNwuK89XsSpIHUiumuxVIIauCKAyaiM0vg+mlSF97ljmRw
i/iQNCA1NwMLY36pYIZKt1MZlDaxtC8MJBigvC9UM/S6pIVozoHmap8YTV0TGZ5pxq5gyk6DkFji
znMBljGj8qN1rBGFMiGkMmN/tUmOI3IhXqz38U5Sc0RlizoURb3LPwjr2sgYKV/uUYg+zQGSb1bR
pHowzcHlITsA3/54RgI2A/KzioBHR7sBlDmLkpWnty9bsrYmLWdmoT/zWtr7PREAcgPDfMf9Vl67
MOU6FhKxOWwRTcmvlMiHHuXYmqVlfsaMsMFcj6JLzkZnsHD2P9DKYOHMJrKEribucsZSETYpDo4Z
iwj8MAwRcL/75ncAnwr5tQ6IkXO8zwT/FUYIsenYEk5ZAUye/AKOBcnyqIR2mJF7ECmSTSEPtxMq
+h8LfQtz+tsWzx4NjTFPjgGhU8Ip6Y7sWI0X0gE7QiM9rEcux6IBoWPmeOWh8NYbvNm0meMiYzr3
GkHkWIccnOpaFOTocBA4tKpzJFN3nj/SjUbG6jzz9MXlgqa7lDTCBPL9ttukdtcsVE+NAqScMadm
VVrFJz0T80LMlkbQzICW9iqn9wsMRs7KJ3igTi7WyhXyFRLku9koo8I4VbVgnwlitd56hFyzdUR7
7IX2uZria9HJXU1lhzcLLPFEXz5AB7WENAHY7KH/yB4dr9aUTZmYBd+Zzs7FlYdLjL1/wiGDbkvx
pDXP9pUaqu7V49kBP4xyJOAZp1UY9j0Y3AlE19j4+q7o5ZElsMjzVpYNCFOJRYUntHMdyQxHudao
yGKjFBz0pSxbxpzguPRoHk6dwwPMFTxP8Gpxm/jG0wmWch3t7bpBc4Ta98Xgn3qnngVpC0zIMjla
trFCU54Cc89Hz/RosV1EUy5C8y1eJ6gj+DmWDBu6wM5hZibE7icJBIQhJyf17rr61Q4Zxv2RLCg0
7jNZoVMj3jX90uKk7gVCBr0PncwVlIt2Gnt00xW0yOYIRepZ2JamkP9lnxUXPxwClS80ZO9k3Byx
6eC6UVuUVgZBmZxfifcNXD8itRXFgISO5lLwNEY0m0i8L4NCIL4SAQnmnO75n+EgzaxetK2/3hb5
N0axEI+Knp4MTYz8tY1pdmIh7vP0thwTr0IR4U5vf82ATKPIRPJClzSGIMWn/eW0br25Ive8oHxv
P/gURI5Uq2PlbBPjZwH7Z213cNrMHtbSe4gegf141xPxoV4Y44oKmCDCy+sgAiTe5WHqt6NFUS/M
MgeJZYC8cgWDAGXFrckKqj2ooXmrME9ezsdFaRg5xP8MGfZJ4To/oseaTzBYD/WBD3VZE/drKB7+
fCfW3VCvvrcwrREyO+nVwbqUQ9nblxNj/RiVMDonT0uFBSuZ6ZMqVOdWq73vYyoGTTO+ovNQs0W9
eL+6nNilWG9PnlMwBE1B2yE8rYbwI/WvfWBf1LHSG/cAv8wAmrFEAQ+Oec7vDtWOLxk0KUn2DWNz
htW1yhw6Uj/71+RAgMTYcoBI+K68Dn4GVNzB/9IrajmwYVSWwaYkkfDrOtoQ+bTxwnqccHf11RAQ
IGXcm+V3VtKmcHKLsg+vLbCEU5HNO07jNcAcBLwIf3+XPutn/rpYVwGRT1e5WFtjfzP0F5tmTNJ+
XXlT53bYTLpwcqFBzcoE+CxEpVtzd9IcN4BXWPIuGBkTpQt6IN0skju0iGG4YrM15AgX316fgi5A
C80W+s9awGRZ6SYzc4e6B4ndITF+vHjULsCBWjawLG/56Po4CIUMFwnULBRsl0tKYIs+dNGxqtP8
uTmX29uk8sq9LfUeP9uVYwPrDHJiui4lfeAV3m6PYenWNzduFletHpMKpMvOUAFwAv0WFNcVb/Zr
+mTfO9Hcd0wqc4qSub0YkO+h+Gac4lnD9iuogJqVJb8vDye3AfxUzL+cvmpSYqyiZp6K7Pr4q61n
FEyKxQeuN/K5QbLQwQ7D++82Q5HNBdk9eOhSLSirdYj4XZ8+bF6Ifh6ciclie2ghrKFwyIelHdz2
R2sCq0Srf5ANMeJDM0gsHrSexX8iaLK1tLYYbnlKAz8BXYSF2fqVgo7aKEj4Bn+MDhmjHr+QlCEc
YPOq0SYwAWnz1q+wHp139GnrW1wyxPt5hPuzTMwZ7W3xIAdGrz6t+H9q7bq/vLyXzzaJcxX4N1tT
EkPXMEWupYPR7zhpSU9FWrnqS8F0idB8qRohRbvzML/TzsooROE0x+6i2T1H0DqD6z+73q8VA10s
v25C+t28lYXsNMr7EVE59qhJzpcG431WJ+3GE5Fi8Aqc/vHyNrLmPkNj+NbGeP5ZwK3dhJu70BJ5
aamqEClILd8VQz3q9qGiqWTsnBqwzy0KZhoi0koLYJYxbd5kgMfr5Oq4q9Da5Lv8RavG9Rmb6smY
3l5LVX+SQtiq+haAlZ1eu3NDOGRCgg9vqtDJDgzuk/030bnE7IRYvCh88X9ANQLa9IHkxeWr26BH
/lr4lotU8HhQUkaj3bvOjAkd45GA+bfc0D5nYYcBGpf16Ya6dMaVOvH/v4snmPUp3bM2chc0Hveu
J8v7570yDqzs+ZveoQwIAKIHlfmTwA4YXYl3gCFc51D1gfztuaOUlxuUmjEAu6V5z10oNUga2qV3
DxUW5xGKjwZlfTMs0gNz14rNb/Zfr2mwsyXWm8WZMEbD7pZv+EaawpwLuVCCpvCG8pJ6XF7kriLa
j1F2WL6VaUOjCG2H7ytuUc9vOjECh4IoO3oTZ49AN/LmFo36NDima18qCw3X9p4DUY4p4iEaSz/J
kedLTfszQkWooWZ6z5P7mqMV2u1cTU+hTF5T4rLALp10kQcAjnu1ASXsRJtPgT1Mugd2RbJ9IZHK
K5dq2G1BAi10TQpvtV8Fk+gs9ifxGmLLHYPd6IbKSIeo9YfkVydcTywpmCxljFX5I/ggAJLapRV5
ecjzTUD1VZCDaXUUOc4gGDhnaq4Mz/QsGhL1EW8pHTmTN87gVLWkYl7fAroTJLoqRq8I4aYRvyGU
+S+BbolKJFm/EtT1nrna2cWn/8SFvUU4zRG/bGbL9c5cf4CTrrKgfjlfZQMCmA1tm1iEJ7YYmRQe
2kGbR0uJLYilvXJTmLyg2MGO/8nRi1w3n06md5zHYyBYKZhQOGsqMPhmfDEPtp84BAFbxxLCHzN7
Pp7GVtezs0fbelfumkdyH3nCtfweujvE8wYMcoI+Ss3AiwZD+hfMKhoygKtSPd/IjzdiMH6KIk9F
LrbNOsJsfIdGZmWSdQJjGoO8ZAKPssAbTacX/Dc2ayXsqkSSgQVK4k22jHO27yFr1EBIW3pnr36+
XOKkbw/BwWsqnkmnxKLjUzbmL0OkrVVFjfmG8+m8V24mdmD60vY9gIRh+dzOp8l4+iWRUaePj3lA
iJO4Gukpo7w1MfsdLq1oc15huAUVtensCrOpoPHph5HM+XiI94tZZsG+vwEm4qGgf/nFz70J35j9
Jz0I7iM/mshCSYEdQ/3UOxnnWZPZeXVAyehS+rIaNo8aeCjwY4gDPtbA9WMCmnB2MMWAUvIQs8mA
b1vNBWiDuT1uGNyWzFcA82YpquxRn3I+72ONqecl6xz1AyFR1wDbUu75rD7vugoVpRfDQ7mYE3Q+
rRuuTape8DXVw78bbCZDAJth3YYqBmtTsjJtH5VToEp9KOLNRfzzf+lH5upV9aLW9oWJYEaGMSY/
npDef51wWwAZ3tJMvOjLc559fLLJZyO9Sbo0DDCWfDSFf/mcUu/FTQcT0YB2BasWM1lmrSA8QpRX
bFb53L8fbCFLrgLQ+gyAq2hccLqnlX0QSbmleZXM0zTOGH2wgq82C6tEtgxbzmSuEA1k5DKpVZuT
IaET2RrCIUWZPu71jPa3OBEv8xGDIB+Wr2N9sPzAoEeFmGppDpW0LOazmvKQAM4nUtF9hUQy3j05
m0wh/GvybDz69GzxmMY94tgEe3npz5pzvhmtPMjM59z9S/MvZjejN+iXqlL8O6CdnGGYkosHDca6
l5QjWFR0gexgbOfVAo6UYLlBlxMS66IVPL/agPmheFBrOCj9dT3YlSQTi790O/bnIa9+EnR2gxjX
yWTR7QRGf8g7Iktk5hPRVgRB2jnN7xr+vl1L9xce/d0ip2n9q6PG0Bd8+0RlRFYj+GbxpdPaSaWE
TfwsNUOQBMzmrJKOnKrVURsblMCG6bRyyVBNwd7Qn1MfS3TyVB0FtoGgaIIEh3RNPMBzCbTCmcC7
c3JhvgxYtBpzUHFpD2HCjamGtpXu2C8CgzFqbPqa8d1n4UvZ+CVsEuZrzb0WC/ewOCL3QPhv7znp
B7UTeHtUWeGU3nb7d+Bw3IWF+/FXpsFmoqtiqN4lXko6h15W+rOSNAtpdOhF9aRRO8eufqSgJE29
hQUAT79+olmJ1n+jfhqIvjHomOA4C0P/3PiqL7yyrfEF4LGF15hryIpP66apzwhkd2L3UDjHTPrI
Gs1BuSRfDmN+3gQWv28wF8m+jezHIcwhhvaGfbP3+A2WsEqWXgrStHSD9joKZAjaroDaGYaUrlw4
nBObWbVz8jaXEiID+Wrc6WhWYXZBwiUATOT9pRbY+OhFwNHktNTrOQ7EzCW6pnsnMkYxf1Nh8SUB
zgibIQe2R443R6mIpsENZizHrw2fX0G28dAzp9FYItacEWDsS9kFarhx+68Jp2Yk6yqhnqPT8NFA
U/u3s45IbUcnxxyavYGtT5CGvz3f61strOe8vp6S+WW3WJ1FDtmqAnMgR5fD3xxM4PhTuhksheYV
qKE5y8ptVw5f5L6ae0p1wHHbr5JssSRZft0TOfM9EH5T13nbD2Gj6vyOb0rwWcAg0P48CTw4xkKw
iGvlznRU6JAFiMgc6VKF6xN7YULa1DhzkvSJjgQXtCW9SAEFfApGIbuToql2uWd1/i8h7/eOELcU
VRrHzgiDU4cEUxV/PrTKObyOnaVgkXOi+wvA0c5eUlICGKHtjTN0sqbbZHHGZsD7mH+YdLYIcIti
//7P8I6YaCkaxOM8cDz7jhR+5cJ5x/YitWHkZl74ybewxTEVhOP++7cjeaAS+095RimyCS5zrAwJ
nddJ0371HG4wd9yJJf+Lwn7yOM5QlUTcoxCLJ3olILL3Y4iIqAcguKdYH0swvXUg8RcAmbipDDLi
YR7pFva4ehA6ehSd6gzlyOnWyHVnm67AyXv78Bze3jMoHpWQqB9Cz3Jnp9IlpUZZv1wtc5JRyhCB
cmSH8s7mAnOAgAQvATagIAsukH+BCYhNpPnESt8vXcidFQCF0I0SQ/T/E/IUMrn63QU/5iCP+WrI
xp2TvcqcTkSRV8mGF8uRntuOr8tBLTdZsma6GaT8j1YhVnAGE3XE8SmzmvMzKGUfEGfQPgxLEGvn
gSb3EE9N9uqzyO0MJ6TOfjk7xhMQiZuCPppHa/URQNYSzHInX28fH/r/DsG6Kz1A5YULn98nNMi/
fqyqxYMJLk8Fjr+6cnuI0UkulnJOc9dKiGViyMl3HFhuEal5G4jZfZCeEoXIwLRatlge3K5wWxVz
HjCl4kITe5q+sWkK3YXvxlC4LZ0TCschUMTtkxtnebqLrlMZ+aFidVuUfzheiq2NcYp7OR7hf6I3
FMe4/5NKATXkOW3/rxP+Ufg4ccxrazZ691Owss3vuLMg9MT68hF1LzQx5HA37BF28iFhEnjdhwj+
gc5MzPvlz7BCBiP09MyicJtx3yww3JgOZFtZ9ex7/4tucFs3dLOflcZHHiUkAkr3Ifo7vNu8fy7/
ailNOEBQDgD1djGmPCAfM6/HRarK4fcuAiSpCxyHcl7Ot67WdsB7kMPSOjgbHlnlWQNxE/YJ6vZB
WlVsbKvAw5mcLImJqf7HXOnrf19VTmOUk+K+gFK6bThruN4CgCp+M9Tb9VgjoCewGkOqx8sbv/ab
cTH6bSKlHbmUeeDVPYuje8fm7utTXc6cTKNGIR6Yp/Sth4bBgGGm/ozVX4VMeB/mVJhirCXWFDfB
Zoh8IJiABbxsJF7QSS8R+J7/d9L6j7i5xXL7m5WnsgfwS0mWVoNXcquuT3aigGURkfaWNB9aSq+3
tRVXGu5Qqrb2D+ujU48LFjhLVe/Zzb9aoTGOi7txR1YK0nQvtwBwic37Q6FmG+Nd54/Keq9a5TcU
RS7himQ9VgJUxCvYzv1jNXUBhx5MzEqjQFmRWGS7TX0XlHphjDzNjECh4fjH5X5dPL3kukM/wT5B
IuuYwPUkuA+0htYh4cUrQa91GniA2LsayRBO/s8Os5k7jcV6YabQAEl3wzUnpr/ulovSDu07A4zb
8YN2jGWAyYx7KRK53DEaidF6HIk+HvDJ13tZbo138QwPI1x8TwGB60Q0Gd1oxtTo+F5ncJ3sgCoR
va5QjWhFV93rU9DnPy4hdhOjMxdRhHcetaBZynWGRqg8ylKYkQ2j+c8GFNWrlzbnMgYawOq5ME08
xffr+I/bRdrqZNeufkjUdRKRq6cRqjudEUH1h1TweyF+WzQkACc4STBvxmETnC0vr9LNEIs+tdUz
+ChhNtq/85FSQdi+xKlhCqQg0oYPSKDmz3H2eIYXaLkDBspsGFvTfK1BnWN3RZ1H1/hLF/EZ1LlR
jxsEr2FrksQw1+e2V1Ox4+IWdjmB2ltwka+OglyNB5//rgdoQmRbuKKu5Cm2pC9aFC5vQIxCAZvj
8lqYHDxGwiW3Dz7RI5wBLOtt4T89WG1rvYcby0GkqElw9k7i1WfMQ3RDZFxzA7A7Kj46yEGxGY2Z
xwWhuZJJT4cNc9fQ08LDqsx9vwwP2o/lMdDzbyI8e6YBLk0RIrsKEpmTUe9yaWGxbevYJ0tfC+TD
bcysBFI+hFLEivg4uTNSCEfMD0IRDkivYPkyn2yqbXkegapnmr6eXWg1jxQRXeTjJ7sM2+WoKuIE
iIkUyKSBzmvUd7BuQCYzyCbaQ5aO7ujjIiTA1TscAEjOLb3RIYrrt35ZJxZJ9Gi9wVKny8YgrkUp
MMM+fOjuMibzmBXwWLCcqQmlDLpiJnPEtg6qn/ql8MTmNcc57u7z2+lzTrCTRLW+hqEj2P0TZ3eV
VcaRl7nZA7e9SlyzJ8RCwJt2+66CZMJZsKr0P5Ohta6gj3CIk4bydvpdaA+oymKbQ7YaNEn6hxMR
jrzgS5+pxbvp2shOoilcLqjazLqNh/cp5oJEBi44xPGB395eGrEvGMh8xY0e4XKxH1WmVoxTVKst
Fah3L6QofzcjdhlwiMLK41eEUbbxvptIhzscmRcHAeJZ2Ki3U2aYaucE2ni1AvMCy/h1fwVsjnQ5
POomoxHCfkuOj7oYNS8uQX1oAxgIzvtluhIyB4FVJxRkN9z/1AatAPE1DtEqZvkxsQ20aEBX6Faj
luls/pqbAjHTAt1m1KfGM3hSTUsCaX7WuPcloFZ9V/uLcsEXZdX0LuW2t6v2XeifIq+6btWOXLZM
ZpoGohOYpuvigcb51BooiatjiEi5SVuf+TwGP6XqFLJQDIN5rDWs18RVtvVwDxQ/K9C/OU8r4YdQ
jda7Uk4yDfDrSP1jZxnRyZBh9i9B9RKJiVlV9NEzC9opXMuOWQEPKev4HIQD7N08drD0v+WoIyVh
++KtsBCBpGmlKdFzswBORFhfVQCxMuWSJluXIOg9ww5D8b1V03wzpvG55+mpcxvwBsLEpmOdN9QV
Wp+JQPGvE7Cb8xMvUmj1R8lK3LWopniAElm/lteNX/5k0isfsxqp3cpmHG0qAUDJyMxwZcVpxWo0
HSSt5PAc5ak+XZQsLToby0bqWXcYqpP2J55v4M0Yx6oi5XF9DQvOsdaTVhpkRNqwtUypuw7BwyEz
5QjJGf3c+TNLwnIfRD3lvRkIZuzCbIBnfv0j3HfOEH2BJpJZMScvUkbtGXLfb/ygZlDU1AzRIfcG
s334qu/FB5Rf4FjKz4P+jsG6n0xZrvRnMmH99CyRgQ/l0W3o5EOVkZDnJK1NfZwT4OOKvwDowie0
4AYDWIdcqA4IEsMR5mSNL3RTp7jdtewP/Uk5X+BGC23f0deSzvUaBsDAjCAJ+BQ5Wa2ouQUzSjyd
lky4kbQ0JEpPq2FMVc59WcrbyUkQ5naZ0iuw00Tm1k8Fbj77OONWNDta8dx3TawYwoSqbcopq8BS
LB8GGTO8Z8LCKIxrbvPu8tJMpE4w5EysTFGvjoE384B/O7FQosNKZ4OtoUbM8DQZR9EFXaIpQ3M8
nnJ/d/9RVeehuNsvuO8QRKlLLBUE83GnoIo6F0PpzXtMRWn1bEQLUp1o/upmp7HUTl6oZkT3+w2Z
0Q4GYhE+DpMOZMlsK65gTB3EluvQ75J+D72cujuZeavb+BxX2mH9UEJ5GW2BkqvCfl0kUju/Y1AF
VnE7bdXdncrs7CTNkCYBHNB1SrJf06lTyJyUU7BHHlqgDnr56Y03qn8F/P5AfwSPN1x3bM/GJchX
iZKja1gRu+4VzRMONMqQknwed5M3H2H0/CYcLXK47gM2/GlaHlJNTllqWCYTLX80vXnnIcplRIId
SV4IYmPi29jRXl+cQuOCFBG5XfHi+ACYImEQQZS7lk3a+tS4RP4IsFjmbvyNrWJFoGdAiQ/sK6kr
FyiSaT6DYOOOwI/1Z1Wj0xobcS/dv1iKP/pow9XIObg889rq90pVa1PJRyHYqw2Z9v5StCje3Wqj
atfZXYMIL1ZW5Y7EKUdR1Wv13qDCtRLgq+Ol7lnJjTCco8hCzZDqOu7QSPK5kedxiIbRZhzv+Fn2
ChXcV556Vo+kRY1QRdhb6VVl8P4YVkhLFx7GrJEAABYtI49qZmgjEIE9hXVF71iGQmjrKe0pK2/1
gCHsqYmhaAXWfUuZoTao9Juonq7ycXzmvG8p3IKhOgpDUMEiWUvr0o90Jof4lHkT66JoZ1OorArP
WMhLThGsDg5l17fXG2tHn/UQlNHbqcW4+0emA2otSl0nbKL+gLjVZoFBjvWcRT+LngbTJINoryoh
MYenEFssOKf0pfL3JSYVB8wDRBnTKfYZY/RIY5eZlPaf2/zTqIbPnSRUMpag3sQxE6oqrJSA72ck
b1FudL88CAYie7rPc5GrTNWekLJsiHUJnln/EveZY5zQAACeLVayZxmTHraYDCc3dCmdD6pZXvFc
OQILoePU6F++BAOoLq9ZvJoqx0wYsXzvj6AJL0BYfOuRgoMoHNdlT5LNhnGm4t1aQEuf+0nI9ovP
gOwOBX74ZHaNobtxz3b2Zt9TYNkvWFDAOOuJvVgPM/dWy3pBw2gzXr1/x4eXKtZhRclwsT4enGwC
GOCv8bz7uBpshmfoTLEblxKXIJScqXlL+FfIzhd3YUUCDPK4CfcoEeB1YQ1QuS2DImWNaviSvcQf
Crl3wkA+M1lWVPZtmdF1HwCHyXLas0uN+vco/VGOqGWQ6uDNntasGuUgPTtK0c8Civ30IE02Iq0h
FcAgOCCiRPYUmrU5PHq2Rs2SRsWgyB3W2D/o7SEyTAHkMnwO51BWAFKCBwW8nrbdNqo6C6Zk2pMc
jdAQBPTquFVf/K1p3n+x30lPzWHNcq33thyWibO1YHg/CuyfJ+lsiOgL5g+WeoN9H7rMoo26Qwri
k/gE9y8vSneq1dzf/masn/k3GukENJ5pnCObwJ1FtMRvJNnIeGEsVcJ/X6IHqlmitSoA6gXkIGnP
XFvsP7klwLQPF+BLXVyqmC23USft9HImQ8tj6YHapLV4y83NxE8WI3/A4rdM/8VkytZxGyGnicrq
zIbmSLguf5O1Bd6AcWhxdez29PWuLey3QvYWV70SPKqyg6E7x5o7aQhuhVfc/d0b8YHC8JwNvlxa
V+THdaDwV+09Y1Ud2j/h0namcWHWNsOSnaMjEQsBysThGqIBUJZNTkUA5696wop1CVUNnyAsB8I4
7QQOC2N+lYaJU8gzlxz5XXjCRGCrXrnf/f2s1YVudzxemgzLKpZyaCrxKh3/DR80s7WGLGx8psux
LaC3TO4lxmXoLN3ZY+h03yRomYY17Jwcbo71415Tjd+Sph2xbwjqWQZPofdI5nWGddOIQ2eLFxbR
f0FNgyBGyvydqkDydDU8K14R1qNBODPc77rbCBHhGfSUVFjsVEZI3J15Ghi4r3RgyGMhfJJ2/zNH
BC5xirNtp0+Tp7ZT/ISvjugxKrs4Nb6t+B+vcd7HklbYvzJOpupLuWX7xT/wqWnDrE8NC7y68ITf
BcwauilAupMHVVPLGEv9xexvrbBPQsIN1eWmdbBST8FZkSDFXMSAFBOWu0O1WoqCp206gB8uedB3
8vqDcUx52BS1f+jCe9x6hCTeKjmKgrx3Ay8a33sKKKK/P3nbxRF2CPRzX+9NvDARRofgwDk36Wvs
ygM7NSdRvc28c3ujvMYPCezgEmgDAd1GM8goZarilNqLaWNvJGT/HNjQBUMdEO19KiNnBzUqD3LB
8OZETcNCrhbNf84Ft7t8HShggfDocuNnpv5nHakpUc7RZZMtVSFX5+jEvKk0ZhuEieaoigBzjtkv
jrvALiW5mGHMeaMSn6ilf9WDLExKoQPSWmMNMXaB2mssQ/3KX0pEh/nomJRGrnrIYpmi0ECEdE+3
7YuhBAM3bJ07+27KIiKxHlfifcTujk6aZciHYiaNTwNvy9D8m2AxQ7UZWMMqIGzNxo2rJjXgcbcb
zHp5S59GiNDqFJMTIue4Ldw4/DHREw62dhwINzCf7yxb53cBfsKIjhFr18VGDQ3LWLZZFz+2h5w9
Im8SOHcdKmT1rBy6/InJcxXVW6TG1qxvm2qimpsff5F24X6SBAbPYEL9ZHslo/fqQ72dzRgEe1lW
ILIvTVuhjr+byQtKUjHATg5/AqBIqi5Vmad/u1/9GocFsAaFpP6u6QUrpvBHttGdzjElwJItpmMu
EIjuXwlLxziLveZo2YFvZJm0af8n/OGHo5XWfzTn8dG83PAu6LgwKgi4r/XrJpKDBa4Gj6pHb4bO
G7CxsqNvquv/nE87tfkGZIz4UQJ6V5C2m9sSdUtvfWU52vHq5T/lc2B9w+FYfwC+B2y58NoPXGor
SDYOFkcdYJqr5u4PZyMRlq8Nj5v+Ybd5eoMzMptIei8eex4IhyXNinfJ9xiac34FE0uI/2WveEfT
8dls2xVeYaOld956kSMUT3dt6WwYm1YDWmYjW+w+ZsIvGWWucpFxZYf6fXM0zMYZ2g55AuaTvUSG
U7burpzng1vNdcImnEz96EtiJl3g4LRN5QmuFNkj0lWt2c66Z+7DcxEL1N0i8RvjTuDIw7aimjgW
jn77MHbQmDF/fUN2FZGBrEjPANtgEiWEgCBlMWfPnMIkqozd7O2HI0dHyjlFjauazSMnI6Xiw/YD
+tOR8P9eK5D6JYjPAT2dpIpFwDNaSsOH45QpsU0RZSJzTUWI3u8SHUuCDO4uqDJYmpu+6MTFGslV
naZu0i0C9NwhdfD9PuvMFoIoXfvckB3OPvdZVudefcQXDptUqKa2sfp0tWyoRDFT1sU4p2R1TsaK
CDhYa6sPbGzqcFC4lquJAMRqSMZovuhsdrkvqQQxcTH4hBYAZugHOtxm/9dAYA9pSxhsQVvX1GU+
1iYnbOk8f6SHF7FtznS0riLVuZYIKRLrwln8ojUm+tJgWjq+QqgIA5dax4pWocTSuHe4OoRJ79Ns
jv3HqTh/iOVGd22oeocOAq45Hi7rIGLus2vGsaR4udgg1/pjiJ8O/FzmXO1d5/Zdqf7BylB4ZOTm
Tc8zL5R9dUS44tlBAWYnrGq87XMB6GQ9C7tHn8XSbe5ksVrJg0a/fPyHezO4SFtamEsqqXDZO9qY
aXR8kcGBEkIZQAm985iw/F6xpwNlHMsVYBenyIAFoPvJCUghXXLEVhWDNonYh/LsMuE0/kkJ4AE1
rL3vU1emQ9oTFBEk4rY0gQ6B3nqxVtJwwmZmLOi1q5o3qC60edF2WXGr1cNzZ2Zy607+OvNoyRg8
rCWfQrwHjOxgK1M8B42LhUwDwnuPN/GZeATGW2YNjlCZKOBH8UdTKL0ZVVhoL5CcZzXENBAWxFLJ
1bYQmgtmLhQv+8I7fbkGx5eosrTGOh0VE7QWP0QCs0mRD3PiDL1gWr7x9XCNLz8axoIVKmUua6Js
dAc2vrQtec/F2wrWRLYJha6/rE0ej26UZRX5+RJQpWgSx/RA/b00ZFHJC0s+PeUt26Mz28bXyvKb
0ktTSVPj5AlUbkTYAlHoufW/k48x7SjAEq4+7MKt++tbbNC89uNNJFx5dg/cR2kL8A1auw3xogAL
ykzKez4r0G0zPnnTAsIYwRXb/XprjAMIPHcBXtyXpUa0LRXO58DkKW8s7qf+d3MGeafYucoMU1Vo
rFvzqCVX+1coC/zQp0YAW3jcPVY6L/w+teOcWowDrpkhu0BWO9VlaFqDeys5VsHGncYWWm0L8wHg
oFVlR6LHhvFsDax+SCzFLxGOTQRDeWZzzNnZO5BfKpB3pdTzojVF99m//m5GEaKJQdZmjNsSIhCb
t5//MMbNbUFunhCKUHOnHpjClfm9FH7l03Uu7KwW2giBnNPOKagD7YHEanGBQYnptxr5jCr3xmOV
kg38c7sVK1I75IustNM24fhguqDFtlmLVv3ImnD9JYS5CtpOw4s6mjjxiVbcimO/rDS2AsGx+3qt
uOWMdnTSuJTT5XykvtDxpt2BJhO9mLgnLiOA/bBB8XD6x/zBLK+m4sYFoSXaI8FkxbvgYz6Pla2o
ogEDutoi6CE1SOHClYGlJnof8kcsQk/pieYiNBeSxrY/H/E8n4pRIbeb/Pbe/Yz8udQZIL+4vukJ
HWqddjsSYwCdkw3OyE5vYMGZwsNua0X0B7WGVxUpt8eDPotqyelRPbqnAEoCSZMDzFb3WJPqvzE+
Bz3d8xJnupfYW+l8a1CQtVqJhIuD5S/SDFZoI2JyzD34Pf5yjAY09BccQ4FZFse0XqNLdqbrp0EM
bueAyHsS3I96sGkcS4nPSSq+Doc6QNj2N9zp/jrPpXHCdqFRmBaoKgQqSD4DjTDCqF5+rfqwzs0R
A5u3x10Frxr4bX4/iQwdAS0LeuePdjDqSHABBEkV2BJ6PHvFLhPIJYfZBJLI1jVn/zqUYHT3NbGN
yMdOBtakuXliD8/w3bp8Ir86vuL6BmJXpWcRmu1hq7NZgtIYHlnNKOcFKJHiIFGF9L+GzohalTXz
vSrTu9WMRbwjPc/R0CeiqmmRNB8mIsfsPdRbpcjx5mQznPKJKt/iv51Hmx+8WIEbSkuxwclRsxeX
h54MyJmES5u+at+hDs6L1r0O0GN33j7FjlZqQhbb/T2bbMH0Dj+8lXKTaGPlTKIb3RRPtdUd4pdU
L316Y9/P+SSzYsAHDPsQv6bkrxRek4Csd527Jkfp/ftAJbhz1eUk7AK9TKaAaq/GEUv+yLFfq9XD
4gRrmj7TUpiSwgtQ/FuGX6lDs+gTvfAVVN2RtaN68mDtPxPYRtJ3da1yAymJ6S2lSRgzHVK5G1qp
TRch+Da8gqTyIZ8t/hTF1673XwCpcSywS3NJTSmslKnRF5p2jsZ1pRXF5HjsVRZ9g7qqZqHuifHr
HfZbbo4XIhHyLjV7YDjKipweUd6jDpHOv9DVXDGjUthzjhhb6nPQ6wriCxX/ZvEra8kYtpHRkgTL
cTO0PCQaNgC3tHighQTlFqRULev4F+HktmWP/Jmv4d4PjOZH3jrE31jDoxrOjVese5omHL6XBxtx
0dTtRjpCLninao87wm64GkJk+0Nl6LJ7JElTNeYoDM4sXbunZ/zyBTd5tOkytQBb3pVuHgM3iXf7
+knbTAkUWNZHcs8xU5bX/FESoQI0CW3Ai01u1IQKASnMNxca5GEey+G43SqGyiD9+n2a5vtdbVfg
JxkspGy+6Ou6Hk+rEZZdnwW/mT3+sHuZ7P3wuO/rBlYYZJxW7C0ASy7lyNxQgTO7XyDaoM6DPCuF
DC5pvEDfXgVelZXHOy+WDImuV/l1d/yVLo96TsQ/Jtl1KDaaaCQmiVBuZbhKCBrwjk4YTX5vyR+f
kIVhc9k3KgSwfYt8hHiO1IpNH9objte3aB2CWESau5N+9on3W/nWSMvZPJvFY1uHQRm8hE0jnfNz
rYteZ1KOQLA+ZySop7/tLhHTZx83BOf6F/uIJRSEoA/eborvY/X8+nsSeVVPjeKAbuVaNk5dlIm/
eeS8rQYsniXCsIuYAA6Ijd9gCzgPE9xhHdqlamLrHCiYJyCg7i1FbmAAK+Ao7sNQmei7C3Pk78+t
Y5ShYf+MkZIO+NKnjn6LCgLTiAs9TiRP9SEcDhVVefrYAk/Am57Q26FjdgIoOHvLd4u9qp9qfJko
NmVskzl4g9MpTZ2bUCUwUTW7c0e6uf1vJ1xu8Tr8Rn32TF/XGXFW5PrYMCCOdeGnaVPSuMrAVN41
rgcG0x/61tan8alrPh5E5K0l/3gcMdEogSu9Z/wvB2xe0FqMZvnpzuVdSBdVF3hnisNhiZ/Gi3ag
O0zP1RY8fZb3Gvndpsu4Y8d6ecBB5PHUm+gk4QiFsjVIXJJqU4iZd3WS3pXa0XgSmFbnzBM2tiDF
DiM7Qa7dAUHX9wQx06OMlHE49SjQJQeR4MnmukNakh75dRcRkJ6S83rydBQZ6sz7QJualzsiNJ5/
hf/QanY2deUIGWB/eZFeEG48gIpg3MxRXYha+pwa/1g3HLrB/6C2E3uDD7DILMoPV8anlXtFmDdk
Rx5aE08TDBv17Pl0vbX3ekScKp3FULAwgqbaNRB+Df5jWkMx8OLC/xLreN7mLfWeduZxmf3JW8Mi
b69okgop5oNGVTqSHm3cpJetSyBSToyQJ8SIwez6ToGm6eq+xpjSwNyrP2XGqJDgEQ+iF58WtGHA
eB027F0u8TRwMkBGIcd79jegeYB9mZwgzi5oWR7G8MbOvAcuqLiQvZNR3V7KiRRGkXW8AB4X3Y5I
J25U8YiWeNDqXPp7zWOf7IwIITvBVIQlCihQ21Lbwq5tG0fLeFN6MIqTLWqV6MuzM2GSYmqQxczA
Qv1fLHF8nrSWsRRKta1slxhRanRy8cZm3JI577oq7m6x1b9sGSZhpkag2FbrxAz7GIZ2ZGfCAu9V
tMtzMyU3rZVG99PaqsFh55i0vtjKzpgtFy/YQoGYKMv23PLP/oxgcTiSkU3ksQD2of+GYX6KyXNX
noa+rBvu+5lEkPw8zCMMXTvKmOdvjI6PPft4gzT5XOytomni6ce02VE1m0n3gNkVOavT18B//dCY
YR7ESxNDdgid2v6qbRGIgseIdeuNg88FVQnXr2zgR1XRCLsrLFKbN0v3GU6VpH0pl0QVb4AsKlmC
Mf0t9vtkEPzfpGLccV9zm9jkGKBPAS0vPtTwVM16NRhjmCyGBP6EF1RvEXGeJxsC8egZUTtpq1Yo
ClcRud0L0HX2rfFQpw6+IjhbknMUnatCfUO5lCLxaRF4t9in5Iw8JvqYy0EqDuq+GDfxHqEAoRle
XOKVDorzSfxwr0ZI0+U1JZCj5pCarhX6lAHotLZBOiMj1R3GPay5FpY4WrSP9jEdw+qU0utHYv7J
MkPpV0auFyGRH5ZOz5vxZIBff+7z2+UOgSKZsy3GoMYV1FgcIx+9ZPy/Ne/K4fFob+tVllXZTYNt
fT3Rkxv3kM+Fq5+EaDBdX4lTH64I1Ea48FdIkornRkUCA6vEx2JV/IVQXaBbzwzlUddA3cWbQu0N
lL/zezKUVtHsg+UoVTW7ubUNpr+CZiXGvtDmdm00+/2qxLKrLtuoxFPEDsx+Dzz1LAhdOkXtHCqP
9Eam8Qf2clQ+UQ+hyTnLldq9P9KZW//tq5YzU+RhgZ7TU2p6fBJSl7KHlXn/OYRfBFRJGu4AXh7I
eLsmZve7VX8HBd3FZwlJ/sbQ5BYu3iFbq7Sn+exkQ0a2qkcvS2Q3Cqe/K536Il2F2OsIu0NKDvDg
E+BrlBLEU7YHg2FO0Drikdwr/9WJKbcjBu9PHABV5zjGyuzyQ1nRb1n3zv+duUVVYFQPZ05oTiPz
lUF1vRtAqAHN254YJvPB/14ryv2xvsLpkwcYIWkFzR80rE3lu8D+67VAZKjErIadRVBwvwlHiRe2
Ojq0FUG6udtD1JX5BgTksmyk/9AJRYFF/zXsGdlMzQRTg8CLwud4j+OjszZSbxE7Ti/Ig9ABHPPf
k/mq8WVjdDf9h2dXTTrq5tgfSajyX6kLbrba906B29ofFvaD4U3FiO0+0NNHps5iU3S5YTuUTBEr
mReR26EDrgT+oEfHQXVZJRZ4YBkFtbfYluE2yKCcD7Wbd2IH33yde+7xhGFhPvI2XsfJ+v0+5EV6
HvRF/ssxjtRuLQeCYftEcmymmpCzj2uC8akB3JEHVfCBMQWGWLOF1HJ00eZIVIaylyFDTlhaDPlj
Bbv6M9jEaw8FQBBbShO7Lcniaova2itDYvIblWDxNB0BSnNJgkb8BFv2ELaB0xOKj99k+vU8rqG9
rxcvFlS9OIF4quGmKJZq4hxkHOc7U1eWSZIZSz5ZQ+khU+D4B2Pm+r1vyDC/UF/ATTfwzckUACwg
iZR31CPqTaUFsdxqiKMFT4ILNJ+vgMCusRM9TPCDZOUb5DhuWWaAXNrhd5sy6UHWKXBE84THBdOm
pURRaBeroWoBpJJdYUrGIHsfO2mQsg9PgppV5gKHlMtxbMLzrudp4wYaE0WdsO4HtbdkqeDk2Rj1
1kaEEHQ2ICIEGLXja0QDqqRwT7O9r1cbw/4FrXxcnhj2ga/oKg1VhheMhf+J3IPc9Nt7xqn4dbGr
4hgJq2CLTbL/KxX8HgLxDvvYePudfEw9I8HeGdJk/meFZUxUJkdj35O/w5DqDsNPnxeQRP7l3Ie0
UP/8hxyAP/45YFSJUSP9pz3INdmAf7jV+qkP8dRrOSXYdpP+GcIIO2KrpVpq74sGH0e0Mg4/qFYI
YhSV5G3wu6yxHV8ptqMP13Lsokd7LI55OZ+squgxGWR91KnJdXrXGBDDapCV35GssdIFlIF+f25O
mDr9Uol4PZ12SHZt4AKgxcl1fjZMN8tM9mn/HCSO88y/vmf/NYY7AhSAfRuyuWwf4Ni622TVg3WV
VkMaEY4+0K7En4tCv01hSp53qqlt/1CZUm86Z9PaXoy1ubuB4uNoabcUZYdr7VjTPleulyaDdTho
rM9+ri1RpIkPntfYTbizGtAu/Rms538j6ga5lvvtsSyz1o/iGoGh7ZNTHDw7irUMSYjiRt/Ak1ba
e/7TtCHc32DCTBRQij4iBkATpiBCb6HGMPQPqCaDCTzHNu0eHix0jVHsI39CBaCe2nGgZ0vmhGNi
0r/LLqG5TsgGcvjtyU5qQZ5gb0qe209om/tk8Oc6C1mNLQVnCvCUxPfZFVxumbdGa1V5GnGI+bHG
f3JswYSop3vJb9obQy2xmx6P2fF6Dtj+0WX9jQwN4FyG4JC7Ru0WVLwj0XJ74tF+Py2hJQhx5Wxj
8Ocglxq112sP5akW7jvq7X1DgMzrzJwd22whIkFkGuCdJ0/F5AJIJJho5ffY+SBC0FtjC+qyxlyn
MQfxkyjAlYgkjsrkc47atxPflSc6w18pvlFZWF9nSYdBGh2pHmGggOv05qitJzWDDiDSO9Cz0WxJ
GB0Ttb063+IXA8aw4fRTJ0p7l25JQyIvwS+eF44L6tf2bUG/KuXTQCuv+MGZuZOGna8zTKMn2ju1
E/eLuLmBcGhg/QzdacQNieX/CDwuCY7ONtdnavBLaiCjP1MADd1RizijXjS5lS2WPQZp13p6nndR
seRje6e1/Cu1SmRDG9TPQ4WIiDjR05nO/gv6j/7gANSJi7tWBv8ZdMsleoWJSnhxDAHiq1+zV4gE
wmI81sgItCa7Cnrlw/708kutiIC2kIv6Sf7IBBLvyJGvUvqSFxDlJY+L6QVfDEu9nXqH39N54LbF
+Bo3B8lQCKbTM0tjLN0L/v9brNgGMJoNAwPXl1Sefrz76cZkRmfys2jc1oeaY/HwFmEJitfrKLoN
GKDBsU+8n4u05r+j+FYFgGEHx87hOMRXbd7k2qrXQm0760DYcFKMlecFrNhCYy+59cZmFBpl2+EF
8olUl2T6uuFG0v7qrqlmOXzKvsZbtiqewDeuiq0sBp799SmXuL5IEpJHkJbRZ/bDe/sQTcadCdqP
bw6DzGXdn55IreToH9r8YQ1kdr3CFG21bYTQQ32SAB00LnlVq37vWTUArXRHoBCStxdSbPQWE7aQ
VNaFsO3642BjO8mtuzU0ipDQZ0rrHtdfECrMEFFs9zCwNL4fqIlvZRMCL99F0dP2Mreaz/fdd0AO
hOK9CKtm8ff/Fdg0akFQsecVuKSg237VlSP0IIerKJHHx0ANwMxUNzrUYHmUfB0gM4afJUpJuu70
FCHsaN870Dkrkp7c5cfsj7kD/NK+zqwZ9SEuz/qELbEasB1QIny1R+V2If6STlD8Bj1SpuFjK20y
CRnLolTdDRlSvw8WhTUfCDl575YD9ez/U/aePezHM+DqWGFaSb1pCq9u9YkI2+0kdm341HyBGD9L
kSE6HHuXbCBaVB7XZg9+V5LX0HYD/fQHLptpH0QWYWvaQf3Yx3lK59E5p8e8K8Dlle/HWlCP9djp
fxKivcVVpeVZOhpky6K+Py57kJ7qVn+l+R2B0/kc16cUCHb5FAylQB8EMKaoIYta+mFkNYJNy1Uy
Y7vgo7MhfWEj51DK787B3CNGDU2mh8nqv9cX6OX5qaV6O5ZMcu4hULPcC6ZeT6UZJxXbBttE2QhE
0129vNIpAPVrhSbb5YhjSM3WsS/u85VW7OyWOyyoyb6Uz9WXzAfTaxd4l8Af3YaKQGUlUZ0yk4YF
RQshrspq7Xuhzd8q3fv2C4qIoVOi0wPARvD4qugN4dA4JURpr8HaNcfI1Eyctk6RxAYi5DHbzEBH
ZM8qGyIuZHaZsbrYDySuzMD0RndPqXI2pfcsaUZXL0djIyKFhpw6jztnw7cT9/Shb3aAHiYmI0qw
zp4p3DKc16HCxjFmf/a0uCZbJ5KKSXO+ThYVRdO0sedRN3hMCYEiYAVfQSLGw3xB6uRa6d8BaSiR
pMGibwdAnErVmeauv1BEC0lxoGXmZE/8o56R1RqNA4f+43NwzzKRuerr2dNiOauj9g1PBSq1AU4k
mVprtg7wVF4jCDZjf4lEEkbC1/eYQohHquyjNl7pDUSJa0+jNHbcYcEtghjz46y7TBmt6Gqn8FlF
UD6T84zp4IRR90kokIuXecrbbhaZ8SsUPe5OMcMeFmGO12G3b//NGmIYH3gcQ/ywKsvNfNXOC2z9
SYV1vtJrPZgazpQgflgP+SRWcQDi4sSw4x3EbMAKOR11MSS7wGdSwp6MeK7xqwYieP/S76wdALcw
tOg85KoIpiJT78QEkTFFXXHYnytgWbiWrWb+Y0u48q2/khFhFp7slESfmBfssMLqPx5Eb6QgoFY6
fPX61IHsFw0M1U1UpMqSB0Lx2zF5WDCut1Y3QfbChA9M/cyp+gQPZIO23yT9I16embqsNgyIutYc
x7IrKgspS1JZFOrkG8fJgDvzNQ8TnMkoXnRStL3/SB8sP3JbgiwYVuo/wPAr1X2IGEJYME6JnGxn
REq8l6mkeG0Wyew+Napd7oxWHN1QPSQGZ+YHTo7sZCAoP4Vvzy78fo8TQW1DRbXymM7vfM+rKg4c
EL01DcLopuzWgUfH28Dqf3aERrRYrNDz/T5MbZY14T/LljRHKEMWoP7Cs1YrCww74U2Ibn0fj1Ts
H+Xsauxw4r7uiv83FNc3FQtm6vYOc7f+zvpTAU24YNaFwQndNcxphXhwXVCxmAOu6DG8lOIRmSix
bDoNnbzEvJIEd6sQhHspnTsGOHr9qAtgHRy6SbHQK3dknx3k8CKTA8TFoxVWKs78UJb9kpwXimo0
hzHhBhMvAXK1tbszBNM5i1sGnIWLjisEGKXZ+gbmuX+jyqdqzsWuapyVFT4b4wzX+eo4a65uvQib
EYWC6YcAeRrZlQHFWm+Ovf8kx2sKmgCZb7YnMF1FX5iqD+GycQMo2fY/74loONPmV1Eoi1G1UjID
GjTTJYiCICLuovJHR+HfPCjqRhYMfwGcFmhRyY0NIdNRdHIG6j8aJlp15i43R3ZQQnkH4d76kf4g
rVn7aQ5mLHm8JaJlzep7Fcr5y4ml05kIzWJbffmXXQEkG2IFtYxH1cN5ps28IfyQEj5Q6qASy1Qe
MuatBAq0HjGErAJzjeF598LGfbjaOlsb5fdkvvGNB71QzHX2WUO5NykqECaPofk792rkQU2b/GLe
BERKM7H4/0Ja6E+mx34jGsVqLEVSG6BX4pqaTMlelbcYRmPrmTPt46hwqxoTNHm5h6ezfAbS7TdJ
nil/h7rLHxqqIAcBMCwnpNPKMkkDzVjBGHLZpp+vcuaj7pLm+llFzKyqYtuAq/QgnkjPyVRJVCp3
/Voix22ev44SdcRTAMOebFBObyoUwpAtwexIf+tYd34f+8uwx64GbZZaJAVwfX7oF5YlBjAPMlbg
EbCsYdXlcsVsvIHWKpxBBfz1x7a9Cnu8+bVUtBCfiUn12SKv7sUZSv5AyVi9hmDmzAXjMI3T89LS
r7NiDwoJSGg3wmfDt/322ZqDyemuvqAX/hkhTk6kB2jOX+0Qcrag00kww27gZmvoAZ7MAYSlB+1U
DVHyfhSO4jtumBgkhfxTIJvrQtJ8axfzBa9nItnB5QAwF/BVJbALLkYJN5QaQvj016dpWHujYHMA
au/pYYQlh9FFgLz/Jr47gcJnHbUgb/Ar7JyEsUNYuP9hWNfnNxy8QRWlwYsqWU3U9l5hBlSPcPdR
k/0XX0xdvf7YK9aFnkLfPU40Z9t74ekWM846atVX0zcOiaO93adGHxhPTBk/pN64pPtQZBCmtDGV
4tl8fEBChJ7JVG7+nrlGbBSs86SkMtB6bx0gxedqRLu3YZFRO0ON99zAdX45Hs0wMtbbpZR+WOiY
lgY0ZaAG4MRTYuSoVnhaExqz0Pb7XRTWydsPe76jgYvuo2ZEaOkww6JgSgY+XwPo6fyh0Undg0RX
g9Ps5Jd7jTpURM1HzXlIi5MPGXrPUq/OaAYFurRWAzqGBbhdXVDHiOrLcam5MmPkGPhA7cD7pkJD
KlOcJmanv+qfOse0EBPIx950yanAy9kCfbr7vOC5A3wHS1YCoR9INnpkbcJ3ofHKCbTuJ9UORkG3
Ea1ewD/JrNUb/K/4eXoKjYV68IaPzz5Lnx8RZIx1VNSep8nSAxanu6V9Q+M/VVOC3dN7HiRsq0vr
mrDncR5NMtWczIe4a+N1KO9+GDWJeeks8ZV+IIQfEETsXn+cOmb5UXZQ0FiMT0lWdhiWbYvL52kI
we7dn7CwcZtVvBsAXl685rZBTe0rSQE09gPY3HzGZjliTcX/PTmdzqFYkNLT2wxVtvQ5HOx7qLeL
TVn3EsAhs793LcCyaXsKIqhtBbHizsezXMNt/kTQ3FlwGKejjlr/oDazONL0hRqm8apX0CHIeLZJ
qG9WXqQww53NOAFf3C0M7MNsPYEBBYZCy+0YYO+kT03jqVWoCeA+8qJ9499n3ROTzlrLQkx96X8F
dmc0MkAJ53bl5MydSVZZ8Llgn/E8gSFbqM/lL/2U7ICEBebtODnNC5bR+7v+2soxuYwulCP/e2ID
sdQGziiNMLQcc7iC5MG5rXpirZqUQcGX+0TnDJ96VmNnesswQ+X4FQVF5RIILspOpU8kMrpljPHj
Ssj+ym1wDei+AIQzyWzaGZX52P3hSwUtcXIXNVapPN37bMWWrewp3iHsX6Vfz8/rWTYM4S7998Fb
dE38nlVuDKKf2sQJ++pjNnhk+81wTM7vnJw2xcbA9q/HAukbYEpRpItt9OuywIa8aB/Mf5sEaPJ2
G1ipBOLaOANR3QCJbjEApi6BLAWMFyUTcXHk+pQqMKpxsznWq/5411lLzQuHTxujia+BldJTBssO
NnSy0FksywY8xCy+Y67aQGM9ZjAW07Hcht4i5VkjMQnarfyBe22ubzDzu9WFcEXPPsff4oM2CDwO
auLIHZaky+Dqf5AvhvR7cJ2ahAL8vEarcULQMAEQKsLnX6qNj/Zot03oKrAS8S11iXbFQ96wPwzb
tLnoBDnpvhwqIazA0r6CLvnke0QUjN40S7otfefG/iAgaFAObGvBA+RS1EGm43ByKP3C/VYk08Ua
2zzsjtwQNkrYk3Ozn9Hxc2ftC3m+EdoUyXmK4IYNTstv1/q0/Y6Gnu5KGi7whWf1Z+bSdVpvQwtO
1popDZvb43zYnSzg60wfa4z6Gd+lfg31/Uew3o/LHrcAGzIPJeGF7XSTjk4tl5qcW4QufERfOhH7
fi+0bFT/P4cOCaWh1RzYRZKlJ6Ldj+3AnaSgtKNonyHQJUaJg2hUN+X+/ePx8LCn9UFfBnxv6mqD
qVTK5Pfm0PBvJjWvRxX61TV+cqG+Vbc0V//GB7U1wQxaHZuXXJKnEVzQyJ0uM/VFJhc1UFzRu83y
yJRTaO6h4PMRXt91NBE/k8uxWFYNQYD2DCZCR+K0XEUnbJlT1vqLRjkSz7k/6a7Z8zHYJ0beu2sf
w2oh9NNNAMEonYZcQ2jENY1ITBhpVlRNIpkUzMe/q4um7wqJxWPwKhKEebOZ2P88dCkLHTTvVVno
3vc4KduxV0IRnAlpcNYxiqSwq5zXSsDMZKf77gMhYoYUbM/x2sLeF1yo/Crp7SDi1/PGR7miQn36
9chcoHWCTHzTxdXp3dQI/+2r5uZKduyAVkLtG9IBY673VXGkqX/QXnaXVg/yRs8560dSlB82Ytd4
0HyvemPIZGRtu93ywV7ZpcLJxnwWkcWd55jSV8km09EzpOQecuklhpri0G12IfAoILktWNPnK0CV
BPJzrzqi8gcbQqRGykifnBmeYCCXfv7YktkH+jW0iWiwnEbNA09CSnAm4JWG1BXmGunrJRDV3yu8
NAwkNiWIyWjHw2sHdyxV0SGKn3yz+ZCnWj8kTR4gNvTmdR2JSx8dQcN1348dSCzX9fcTq9Miq93/
kXrZCxtZ9zVmyXHlYOt74yHOAg+gGZOHWiZEORVkSqn3mKZJ7bAa5gJUSuI7slWcEKWaxfLrkwQP
PoKM+yJmTpF9fnUTA7kAbYrT2Rc1WMMB9htYYGavrINWC04B9QurcODPT+eOGnMWQgoehjd3fteY
r6/76iypIPwSHLaw2Qpz1kMTPkeFvfWpMCFmHOfqqR8hPyARggBc6naY4OEc0OTMt/myFmyhZb6C
xnW8C8GVP1wOCj0f9sR54pQmzJMKyzy3awTbGFvXhg7WRg04q6jqsq/8tKAWBlyzoBS2uWLHpDJm
aqw96ZR8ZnzpoEmIGZ51I0JI2wIyPc7/VSh7aREH7gNhvnStpNhi+tY/5Tg7Dfo1RXlWgpKd5zrf
TNw5YiOJqijD4aW6IvT4dL+b0SsDeF2dyZc70ZKZTGBMhhYlSUwqwKekXIU9HBPXa5nnndUbkyxw
QWbrg8Kmts8LeYYaoDxGSCYC4lwRbn8nv2cVhTDZ93MhEVO1nfofhW8HVANYFKg7SM8hCtVku9XB
DMaEskEvFhckA6F4RYGjr+yT2LIKNznnkxmaoJml+7MVVTH+8WsjVpZWGyJDUwOKrHrIF5GaDjZo
SGov4UyETBd94P/emnAnkDRabOH4A2hj/oP09YGDwkaSei13lPrfRtWyp7r4wG+13m8Gt+s/9kmk
skTW7kEMRahmMf4x3ivE969JlhF1r21gDGL5ngUP6B0a20Lf15FglML+fyPx4TwmaSK/yNr/0gsO
0idj8gwJO+Xmyc3hPC2LCcOYNMHl5BQduPtKjj/ApBAYbZswpkLQt1VCXuG0LN0FI55G3uAHB/U3
TKAw6p1zugmlQnzPtJ6ly5+sReACKJwRmU0MfJG7q4LtXoRIKxMPSizAui5v2Ik5soIjFpm13dRP
HMfnAoEXV1Yvw0BLmFnpSgFZvQYtp7nMHsqHUPSTX4zRLc8jh5/pa2sZwLEeNWMJ/FBlWGDY2v0d
ZioJIsXWjY8ftQGycI1n4l7i5zNe8+omTmSlixEgWD7BFWQ0LCxFPfcTN4wp7XHOpdSe/BoqT5JC
6yRrJMnCb43QhPfcA6bu/zhlSClWm1TB9Hm1GIgB9dhlet48t2S+yRvrRrQjCs5wXbHPqTEQbHmr
yN+s/g/T/a3jHUDCP0RLfLUdZQ81vyUqTQJg+ZAOT5eKWsetudItJVMrbwgU8qGcEsMu4LI5UOb7
pH1AKmZZ4vQyCW1O2xFbsoT64kZwFa7Nyqq34B+OKr4juUqr4+pvUF7/y1kac4h/oEuK5MNcpM08
icaRwKHpfEYfW9v2rily3wa7ZI42aU3fb6f5xw3qbx9+3yQZ2Q5rIzCijQzz/fq4hGOiVLmNXyG5
bQEmgYtIXCMbP7h66puAdviQpfRXQnaP6/CaVasASnl8gWKvWisQcyY98IHpbtYOL7gVKOidEXjz
PxbXfEuPHt4Q8f8BzuzL/SPfxEu6f+7cf6ArCgeVhcJI2qt8i4Bb3pmzFehsBrjSyvUlsHDhCeUR
Nr9uk69LmhhBAMVzQ2xIimpawvgFQXtyjvI6WlnJJq/2wVdzK4jHObcb6ZllANR4a8MB7Zgq6fw2
wBEPX5vsE7ahUGaV6Ktx0ouNvJ/kRPqwIwMPmze8mMKgmypvrGjl7prBRTdIu/b+gBNW6nWUsh05
2dSo0+BKCU1PAEXGjHuRzYDxv/EqCoazXGvZN36wmc99a0DTJySNZot8m6c9fQLJ8GkCOlWHUva4
t+v1MB4Ijsrwg8KfSgIR78t4Zo5bDaVcHzftml/5bBLIBowie/QpeCR4I/+pcRspDHcn82KH43Y9
jSzsGZk/eLZK9HI10uGH0tYiw3XohxEqYEpMy5V/VNO/OSstfPibnYhVdl9qaeB+dVte1jsqlHP7
YGiiRNSe23vFl5B8gOiP2eNMkg6MHSHzeRJzaOXOzJVsQCnrSg+ltD6Oc+WEdAkyyooYEJdE6Hl+
Qu3cmn+5s8V4MTfic/VW6h6b+mDG82q+GUOV9YlKoNhXPK/w78pOjXVBwwp2OChOMf3GDnkHX2JV
lcKIUFpK+IrML9UoJ5qmZu0USitjsB5qXqxM6w8rFYJ/D2DMGnEsvEptV/b3x6YpOEXaHDijoKac
Qpcto88rDzBMOGzNxZsq1wPs55AugqePyRdcFqcQ4mD9/gyFlYT62r3m4dcLInl+no9VMrZiRMUO
/19xbHMJXloJPOc3ceZeBlj2rlv4xxHFSHHY/OLDGdMEE0m5cB3QkGB3z6SPFItHb6avAGZNpBjz
uF7HiIaME7FPpUU8eaQYVEmPsdbJOV45M5VnDcuRKQX5fz7sAi9sgV5BzRf5B4chDGN/24Iq5cGQ
A5yGK97gQv2sQaWbqjOchUw+9IRakfPGvQkNXg04VRRjz3z23BelDD4xdwTmLKdg3m/MWK+99ujT
nFmEH3Gq1sLbfOA7J2eFNa0UkZSoUnuQSAg/ualP8UBQQ5uIpOjB15JIdlBVewQ4uur4FKu15Ylq
AxDz/l0aSizLkm4ZHTXlDtWrLBIn5BT6Atk6XzYjJdLwWetio3/w6p9rN87k1Z0H84l3qJwdTkRC
f3vifRkdCN8oWu5cPTkHepvXasLBDbnopQIWE4Heas3n/DwKVKZP1c8OYT5E+5ewBg9ONVgbwmEq
QMxq3E9EAXr+BPkPSXE/jr2oajkR96jKoir6008+7hJENeRHN2inP85eyLGHbmHxhfk5Ke9n4aFT
CuVqz5hFbVCbMul8UgeeUAR4dspB21cj42RHJkIlEmCkn8stKSwuTQHPJ9/q5Nj+stFILHywsuiR
3qC/pX0XoxupOTYUQ1Hh2nizIWCAV+8Fl0nOrR6N04fzAiZpsmLR0dV97gXybY3XKh7TZtCcqVdh
ZnCFAWmwTNybWy9m0wurv59Lp3JarEWCFozIkeMol2eoPWRRn5wSSamrFm3E8ytNcqITM4c03zYU
SGffW5lgOpOPnNE5TnRgjYAtlbmhxJoL0DbI55v26ubBFvFjWz49kOXusb4WnxNJI/t79sIHwBzX
G1bZaIN7uJZj7bXXQHzejIcliLEfBhZVD51djRCDbvOM14eazSF3Sf9YR50fA5jhhIIkXnB3OXIf
gMz5n7ZLR9GW540kW8SxihY+FGvwpL9wB8iEgC6lgAFRKvAAUya//gBra6nokwN7PNXAfxN2+WYz
5bCANWWp5lrp5Y+3OnsTbzFKJL8ePTtlC3dvqg7Od3w8zjUdxZNSIM1jPB+NZ8BPpeX804wqG2ZY
PmjIauTj9+bM/0ePgYJOlB7COaz8JyeMIcjwvkeVFY9ibjcMUterYtcv5PeF2+fQiomrOQNfU7Kq
biPoyXCMaOh32j6DsV36pys2gcDiLJWxVOfvEWDo3emsJPP4HVXaV3OedfJEqMvGf/8WGId2vRz3
DknHfX/kqS6DIbj9XG890wmksj6g0GC4MxavgOxoY4c0ZLnZu7QkMpoG8qLp8+IZld0byY1puDhI
Z+gYVp8WbVGGTCXGXbJcnLzm+PvyLvSogUxfFjGZzTyamYnWWYgW153gQ9ktVK+FK2YMykCljDH6
u/Qe9s5YgkjMSv4FTeh/kD5R1XWkAOzLW+v86itRqdoXf3AG1Tilsau97wK32DB912YmWI8jlqv1
V7xEUYpPMAJesx7Zpnmj9n3mUZAqwOFlFvvi/BrgWQjR0lSq3OYZuGQRMtoXXwbkruaqwug6R9kS
Ge6cD4yBq6tYUYtGP3UoM/BMPXD28GkE599vGYqRyo1IIjqCRfvda4e68aSTraZtsIx6bq4oTr3l
HRzG9XQXhh8dKS1DnhG8If2mDNWt/HC6S6TlZkKoBiaiOPINR67/vyaa9fZnJGdcTW6fVPDdkb1x
ZAhk55Nal1BRwErIiE/XG+EYxuV/jFEUo2CAc4LIlx25ROfItdaNTxyrFCBrPf/xRD2oeiliW+cT
EW7pKMwpfRWmaO8908sYbkfCxIh7NhAH9vMl/0B9GmFu0NiTOKhR1IHSQvWgSHFtmovd96eHkD0d
6fN0SmEbFlyeaLQCUUju1QMnefWUspYn17Iw72s8dWthLA+XPGq/l5+ylpMYjtG+zoFls2JIpBmQ
U9tAHpYTV1sAQLdlowShBneJ6jvOXbLUoj6WboUYXgn+EEnpSz2/m2ugjpOmZsRmGEPQHuaM+RA8
Rma8ITq5aE9KG0x1uwNqLljApVecSnvrpKPV4mSqFmma8MAk6uz/wkgd7b6FQmwPW0GD2ta8J/m5
ApVnwZM2BCoa4cx5gjK4aH5UiB8O0lARZpsg/6iUZ1ylRgiB2+SYPLc3DdZYRsUgAqJ3skyue+fW
9DkMywZbTzixHSb38yYgzfSZGkNb1Gjw1VeEOTmg2shSDrzhvA0j2q2A5bK9Syr9QJOENhubJqky
TaZkPQzX6BeCJU7MyVmNQ/Y/hh0EwSDu8dyRFGdpdXVNAmDi4vbrtkhtI1MHEOJRbfoV7FKhobCR
a3socdTgkGfhEaSIbdNI1grsOiYNvghCeo1/2DokYrp2hGvQSctNCNeUp71rJZhUYikXzunyh1Op
/h5t5xLxqexSxCz79ELu/OhPwZrehotk9MZCV7mgZZOGCWZfr5/laQJQmsSgC03ZcjSFGC3PkWD6
Kzm8ViZqXVW9bM/15jXfIJgdmsoH0sXbRsoaGxftISGfBBQxdCSObKdJV3GOvpeE/vG+1fZSJYFe
3wnK8XRvZGatA7E2+IfzFk1aSdYREfpYL2PjV5H/fcSZ8hrDRQZ78laIWfYTWgNCSKVNhv6qNWBG
j0ZPs3ewDnWUqqFVUZfjD75pXtQilKOOYFu8N/HgQADH0Z+EU5LkkjP53/NXqfaQZSF4xrifD7Wt
EAaSZq+2lcd2eDjmYbUI8+mEy18kcNaldbThjEv/OvaaY6EGN6oYQqdmM6QmAvEU+e1cQoBS2+2G
mKAxtifpAWURZULsWWcsxNJudq2D4R6TQ+5TDf1ML02IZHehPpR54ohQ95nRLTYdNr3SeKydQwR4
Bv0IMpiBKTvSIKozgIxIO4MVfe/QEwfvuXS0HPmhJtZgAqyOEgvlG8KdfKbQSbnwSFNOvOduwLvU
UcAKef+ZiBrD4pjzkDIaca9wQV4CeD6o2sKcVLq3e5JqAxtz70h6esCOx9u0HR0k9dW/97lzpTVO
aRJwh3RKK0/XBz0SKLvdd7yEiMsFADCdz8zm0/jWXT8um9rRLClOkeZWlLuDMAOJZHopTNHz5SI7
61ZOdkymWxZegI36JFqvqKKkayZWaoOWQfJiZafnOt0Rhxzc4VEPDcfUEpsHtGJIjOqFvf97/Iu9
Ie919AB6WS+XVZ/Im7DjbKecGg/Cwo54RKsDwNVjxa3OPZXCLJFtrk3l/puTT1sjbXcwuI/+a4Vp
WvrdesKfw0zTYY+GcuMqKVLpstsjWhncrZjBxW/YFDYWOKYUBKNlWPHgHWEbPGfiKC3n8WLJyvi8
8yUtoXpuOgPh9ZVIcUGujUPADUCtXLx9pJSR09uxUE8sIuUYSWEOei8HJ5yMEOZq1FSwHAzDQUN/
sdj6AEszR6riYgp2ml0Vvyd5gsdvP5n2CBSGKtDZYL17rzWhX8LSEIO4qjlolrPrV34TNUZn54rX
RPCavIQ+6AGCyawe0m7f8bhq4j0/kUixS2bORgMJMWd2J+QjjirNgfRUuJEkXU7AYEp1jTBa6xFv
ArHg567jqcAdA9HaVn6vp+/2+ctOn+Hu2/I9OJzWRqLiWFLpLfkgTN4G7EtZrpbKSM8TGzifWD/Z
/id0Bl/MK7Zni62O+SVIOM1qhwi5zgY1X0if5vWcKh2Xu/oVQ53PgFo9PpsRGYQt8iZyCYW6IApF
AnmAKJQg9VkbgJ+VstM00d9tJomHcMp2JwAin8qztbl0pNwB7p5hpz7QOgPRRTKOKpmIQrTJy+s0
PjPAF8Y+hneOuS1CHQm894g7eFfIYKbsmg8Cz+dIxYmpPy4e44wOND8VjGgUvkkECY931Po7/bqE
dEXiRnK7lll1znkL84xgTvnp3WcoH0+YY0487I7NFQtUqQCdtpq3to5Tbq+q/GDACGhu5PzfLNfl
gmsynjWkki+Tmue+2biVVJwcFpftgqBL+5dTTqHFr4vcLEK4lqiMIGhc0PiHPkITQm4WQpXrVUM2
X9IibdQP9gcqC82qdPyoj85266+Yju53T06IcRpXJ15UrfZLRQXYcDJmG/tQbmlQMFi3F6vawtqs
+fcs8hWuXr6d/1z9KK7YoHKIb1CQ/rT0dRNLAife4sDSgxnQYLaanjPxADW2vjN7AKch3K4XWFSz
23PkjFcHZ+yhkZ3RsvBFZzUdfpzn8SKvYriejoBXPpipJAre/xDsBW1dxZKEcWP+PGFHbCXfH0ny
iFcrXKJ4PwlAzy/98vDcCn3k+Tg+lJB2i17ljwVuvSLbP3XzDCBV9l0O2Z3mWPWMXdGxIMF2pjVE
GcW+1YVZ924OQbOpsSMtNa8C6RHeIGpjRF6BM4exiWjxFvCs5v2ryXEG39Ntlbpz5cKK6N8wRYbN
4kFyqQEEYQVtBytgSAzRM5NaHWP8dIDe96f6hB0T1LTnur+HlMS0w51TLXM6BYcvYnV2BfP4+S+l
p+0l5/GHjeMxXF48Iuubo4aFkklF4TkGBX9DVbGVO23zheM9taXMis3PQpuLvu6hgcEhuOWYj31W
DxvlkgF5HEf4wlTpTgLBX1KySNIc2dGDcTr5LsXL/fbQcfFf0mkeBHHrwwggPmj1Ag6H7h8+oWEG
EZx7vqcTx2O8nT0eg58SxI1x/ZpqrG2lr4yx0JaQ++AxNOA4JVYdxnCfhinwHZ80Cr1PgtnI+GJI
YjXLaMb2CuiTsT9Qu++94tLozWSdiBx2raNFbt51/+bLoSR9om7sjqFEa1DJ4/UQoHv9ryZ97yXM
DCeLWZ0pq+OrosnHzCTCcMQIgHSJhqstw7oN89Quo3QdiuquHhERGOIblV0dE6tr7BrxVGMuoypZ
3et7sdTQ5Oj7yJgwGt1prPXv9k11SeWEd+oUaci2DaS98j0nUJIKFRqhfHXJrXxq6dickzcs23n+
QcYuJe2vPF/xdkFEdMAAeS9EUllHCwAMbcdezzSo5eDmVov6xMVIDUPz0cB1kTVGhzqTdAX/ZyJi
W99Dd3O3VQNfK4nPdWLZHXi/jDW1aoxkfcMc5aE44bxgl4xste4QDbx39rkwmIoleJprf4NtMr2L
1l3rgHuZGbTrEbq4AyiEqpl+cn8+KrMpAoqBtXV92a0faorBba8vnu87WOSxIweaCywd/zmefr8c
PbA2tgIOSctmsZq8swOGdY4tltVOeSr2B2YkWD2cEgUjQxbYDcPpky7e0dGECguYxcKzSfc0Mavw
qsEetAwiQ8wt6UajYeduydPeSHXtCwgKGh2QvkVCFo6SB7d0fb/VNqq/hXavVFNWKYqKZrFbYSya
24jc+liA7VxeCPGS7isjiROOGlUnFFW+nd4r7lp8xbVRv3JEp5WT2CEIlMugTZXm0B086WuXZcQj
xtYWPKfNyjMuJykNHMDSPP8Qk5O0CpN1UQ0xm73ZTUO0HQG9v3ce6rvoA1AvZIpbCDFMZSlVb0aH
jzlgdEFkCgp0ikGg5cEGjh93T7atQUYjgrvOonUMzDbIxcjnN6Fey8AxUT4+KDKdOit5K2+BCNBs
p8UX3tpdHNV0eRKWJAovJXYXQ0lF657UKfQZJGqgDe1ewJp/65VKKbvI4xyueokMb5Dp5/tCtg21
SZs5YYMoyNUqC451hXW5nZeM8HgcgHHIljvQRUWXjNk1bLwHUtlUMIxHoHnO4yIYpjOR2gy5iEI1
1/oLhsh7A8s8Hkk4wAdtVf9Q97gn0/4IWUphCY520WcIYYrxxTl+00bLejh9COdhnGUr1bxEWOyL
H7RU6D7DWyNw+vbKsC1/J42bcCeupGsipC5sXU5dU1knutrBYA50qCUMXnvoyFS6Vs0725M9d3hc
WNmc40PaAFvj5YT2mOWwPvM5gEqiM1lWB/SM033Lrmx3uH7ftjITMAilvd/6sBSGDHFdZCiuYyx+
JnHrY3Ex2Et4qkn+UhM1ahMU2rpJaypJ0Vw/Xsvugrov0UfuAf5b/P9CjlKHz5UgwIpjLo7kVSyN
5c27GoQ1m2iNVN85E41bDrQL4xIu0d2DJjyKP/vzBk2kHGOdAH5Yw9T0NNqer7z0QJW/gkistswz
vGXXV69mj209md7C5B0BAF3Xoge0ynB1KfqK56JcpfgYLZ3W+qWe51WiWUuAve8A7SeaiOTT9jf2
+PFdum+dp+h7cSAUKOpQYgOsFw042xZ7xxaT/H5UlbXrPKO0DiVzi/2X9NZu/CIXs1dpbyRWJTYE
xQL8jvx3aOZCY7Cqc5ZERsc06Q57MM6ZX4KitboYdchorhU/09YzEJqltzhzTdUXj7WoMnbFo2Fy
ZUo1TxWzFVhHKrXN/DgwfrvmzpXBqPghJ78SlzvDq+3wXyjcCn+BP+mLWaAAUh7RviHZq2Z2reDF
7z8jEpgDy/pcpAZ2MgrD0fSoikwfi8fxSa6QhfYzZHAmexcNCqPas9fcPv2gyDbw5y0/BnfDaNp+
qSzI2Gd3GWILymEvCOheTSjZpXb5e24Eixxx4U3ievPXyn6MYU5B5fbuaj1A3F9IIsh/FbNEyYzi
V5YbC4L1mwXMqxwboXcm/o7FK+itGPUUSfPJNM0GF1IA6SiThdY6JSHcxdEMTwvR2FWXVCGmEp65
3i3DGRyCPY+Wro8lP4Zgf1i7ZWMb+2Oe4MJZIsUOtyTgrWjuprJHdfEcAd6vo9AOne+VgFG73sjJ
CntcdsiU75GLeVSTyezr6NqZx1vduyQTeK6VZvtgqoCuSaP0RxJmC+sB25oTd/r26CSje7CghZzy
giB8/ICQYR6s1a6vEs+93yU2tUITXzSPIJ8O388WqtY49VRQkWqxaK5Gk4+kMtQd1Mt1GtzQlp/6
JxT3Xu5Gi50saZUWysh7GH4cfcLxFBsSlH/LBaIrDaORazPXpfwGtsE/MQJKxJDSIrhtyeGH4ox/
vYdfg07T1jCd78xyRELQwNuaMYgt6p5qZo4ju1SpwAlXZJsjpNMeJYE9bljZ0oECxPqMLedASiHo
gSTTwSA59xWevZoUVp7f3CnGI1OkRvbvqQXdKG44E4oL4THtjV4sA2Af2I1P4vYv7dASxkc9X8F2
ZLsnfUXU6ygosWrrutJRKPhvIt1HO3iDl1kKTy/D5tQG5UQrRzGKR4xS/4B5inXkTGP92ud62zPz
0kZqWhHc2xjRBckq2rQVUfQHYrLBMPt7bqDceAfCy7uch0+4e5inQ2UnGzmvyYmUMy/uDHmyu3Mp
Nuw5nfiAM3/wGZYQ0O5r4pyzGJBoeVN1WYBiUKiMTCP9keI7DUIRKuMSlDXJ8rrKdXwmRQvaO99Z
OzwULEegaTx4eYhPiBI19K6cyqUkQ5FEufkFhoktKEBp+QEd3gUsu/1+/95YM50Vyo03slzc1ctL
OkK1E4y2zVfoNEFqW7X7i5JKssWPT0b3ZStxIFjsHS/AAcWILvgwpo5jfH/49THqsqA6W7hvfdlQ
xZBM3YRRhTR7nIo4+MUqswc9MViwGuRFMvqKts5Oqi/J3EeEBI7KRTfHG/M0/p3waJyl/xXHc7c4
FzC9zfTHbrKK0nk7s1PYUfhFNPO/AzuUPGJFmOO606DFm9dAyu8OrkVhDhaz5WiyADXeRyQQPajm
CcBTdgJf165CxEQlFfWPgs9l1FUMoleiu/cyYks8DO/iV5S3ShPZRVqXJk66cOD2GHRqHC+E1bpF
N78UynNcGUy3NyX5CPP+U5s20g8WyhRtr2Vk2scpHaeLZJM/DS9OHlJBZyQTmIOeP2mcdQZXX7XK
weWuLCoxDM72y8kmCDIvR0jg3Fr3F0g9Va1bQsiZDpkoS/IIkn2wo4nE8HZrnGCP2+slrEUV1FtK
sFHUIH+7/sb4B20oY59yG3I36uvQ+nM+KT51ju3IMi/LPzWcBMc8Xns6HNu75fqUXlSwqTjAvgoq
cmEQL5+F2r1oi5SXLjz3Gm7BA0xOl96BWMiyVmbhxJAcA8b0ZjxYKwMkAxTz6ilNfdlH9yaivxlG
LWBlME5VvolP5V9AWsgydZ3m1RKLsM8CQTFHNp0Hs8EkFSzsB9ndooWkMJUEhhLSJsjPRpYfuNma
oM0aKEysFg2kgUVyob13V/lr3KP+Zw8BASwMlPc8k46JFYdIvB7vad3nBkSgEeXXuS72njalQEuY
8pYcnDDWmypYCIdz/7dMjF09G0qVjch8AH0k2yjUkGFVG/91VG+dC36kCs03Bm22Opm5Ou21IO/d
57f9xso5mKDOopGMLaJayYn7lwgwC9Jnq2S3GAfio0bvy5+F7iuaQw9wJ05bBKOI5cM51f4BEwS8
IpT0qvuVMWDWBnNSdNAJIKcdkrmz8GMAThNjcsIvFukidANfw6v+LTpYC6KxzEkPYl0xqYaY1xk5
5b7OFH5RU0CNBq8/YjWr0sRUx+fbCTyI1oS+YLXOSPmVBzFmsgMkUwXzYdXgnF8lz4rdRAhJRB7V
ugdlPPaCHYY/9JxbX+n0WbiRO7ttuOkrpPkFa6yzp+n//6/d38r4Y8nAEYV3XqzrP32nHDtkMqbY
M0zT2Vy0qNLuBEWMkJoSgDGjg4d4u6tVJkEqxWHBnYWXAYZYm5rdaGKlbQzGg7hL1pxGI6x+dclz
oILQ26onhnvfvvWsG073h7n+GkIO+qIEc2fFsCP+a0VujBZLomljUyYDC2K3jWYcARomqzGh8WAE
bdhKox/Ti8fMJGe0TUarv+yqxRzzzY+f7h7Pwhj42Ey87aqrJ3QKztXc5uWvCxsmPWvDMCutuSmq
tPbJXheibpaWtYf2cVAmo0oMjjl8ZAtSiEonqJmO4VxeLDPPOkpsokH6Za4IPTgjjB6Wi8YiM55K
pOJ4+de/wWTMzMZmhMDrBY091uLA9a6pTvActtl7UjYT3tUCPxccuOnLVsg0DqMkiNEUVQPEjBYv
B94/wb4ZD9InUvNECTOYG471LAvVLBXzq/c/dKnAdLNdKyhlzGs0SGusrwKjWg2mRIKu+CTyjvxz
6+dIHdlMiQyOkda0XSJD+KFXxEyFmHBlem3HNHk5orxNYpKrtZny7lWi43dEtH9Z7fmJ3fx6MI1q
mmsUu5HlNVYxfbQJTkecaOr1dd2Ma9mHyCWrzisI9Kh3zjcr2ZCdSfnm7doMOwv716+4A0PPX+C6
2Dyg/LK0uuihF3S1dMcBbNusH2RkK7M8+WIqwfrjnuemJqCgSSO3Kmdzs80ovHNTEnABSzkFIewp
LcB9CcvOc56BuITIiOSZiw35HEFGOyMMyyEeY8K7pOZ+bkb4UrMNohOinXTExnsYAMvEXBo6EoY3
G6644eImMD8UWSh9CWFn1j+X1FTRxSxTPjrLCvMyMGTgU8C8L5pBmElodTEb49vf4HtYDMHQcuS6
dJ/U9OFjGcpht7ugqjmlkKpSB+QoIGBWzp1Ywtqn3WSw0RcsM5GV95D2VXjGckhfzhyquCRtJzWx
Zkg0LZ0JyQSyGgDvUzZL+r89wz2lY8ioxqhgmCI4MGEg9TDn5DVd6xssBiMWDaxq26N8RZf8knbW
p4Q81g1y0aVWBqZjHpwjUIKQOXtVLDbY/X+sYXwplYYAuJQmRURgc1bxtdjYmVA6BR1fZEoLokRW
JUd8Wx4I49t4aV3yjCVREVwyVPpqUyXH76fyZ73VDtjW4IGIfsBlnP08P2zWOHBv9Mo2OPiR+rbR
e8ZcKhXVB1kqu6rFfFpY+emm777Gy4irNx0FHjnNlOTjPJMbJAk5o29+80cHZro+ucOExqoQ/MAf
+tW5ivx2bG05lGpOI4P0f6qH9VuCNMCvw9o5xIQuEv1yZdIE0uRFCafXdniI+SyGnPYh3e6Zogg1
S5aHjs7v/Cp28TQx8fQ8ZvKu+8IOjiNmEddSngcOxR+485RXrx6ZPQ20w6CGCZAr71/s8lJ/k1Pt
1j75GG2AY8JmmYXAQEpizZNIAG7JDHe50pZPNW627sWzsqSDMc/1czaTxNL1C7NeAxMTnrmbCz6U
1DrNP8qB4PVul6q4X7ye2CDTWcY+Ygq99afDm1TyVaPXeRLZ1UnaIHA2HKtH6TlqPEPZ4M9zDXw+
pHuYbgjM+2a3k10W9rrC2aJMfsdq+o5oDHauE9s01abIgDK5+X5NpSstl0pamR2b0oLT1Wjgm/RB
yqg2P9WSLyJNjg38uoALL9arhoaEGn6HJdYI5TLt+xHPFbQUtBDILu9RQkSF5f7TsA4SSsHPiSCb
awy+6GAj5Ht/1Y/ctQvd4o94gskdanjiHZY0oE7/W3KLTo2awE+Bi3pauTzXAkKleH+QX/j6cFeA
RnSVfNuqaZYMrhSYdB0mm0NjydtXcW6D5gQxId8magUadU3klyUTAHdjMROdZdXvKmvonR5B365o
qqdYZIE+coGbHne1np7igBd9vHBHyr918OUcj2KFqMywxza1jE15va8l7WwZZAsnRm8BALQWz2jz
zK3qHRZP2rnKcAHe2xy0IUEl247qeCgaSTV40IhoeLigoUZnuFWYh1w7hiz2RmQyUA8rl9US4U1U
A2WvR6dUuALBhyqCqWCWE9TML9kvFcFsRbGD8y9eTX5RNkyvv43ibam8QGAzTIrAtNM6gHIonk0k
oi4MHxz0rEnmg5Neg9J+udT3lOWL+vhko+eossZSr3tUdrC3dX6hL90A9MikCJxoJ+kCsrpcninI
msJ9gM5lWhcBknLxFJOpMHPVvaQ9Lq6/mKtMB5jEgpRTnqSICY7ipeqq+GxRpDEWv4cLWbYBQTB8
CtQvnU5rShmHXwOVO5HRjjxZHKWwQctyEkNPa1FQPB8uom+ie+FkYG0bECO092LFvYwo+443Bedd
Ty+nTk0CYTB6j0lCRNLDsiHXU6tpElHOKLvQcBSK213PkHqDzco0Kiu0cofAIagNNWGxt9vogN6T
On7XOpUAxu1rBfpfP95qfIRcWL6VynaXsV/dJyoFc8rPj/DB4QGV4sL8dEE0HhP9Hrp8miuxjVXu
HrumPf4eHyzpNouEh10r1hOsSQl4XXihphbHF6teRMRFglB3kdFRNrG1SJC/LR6dXz195P3XdtdO
ORLnOgcgTtlg30VWD1C3z6Dvt16M2xIlzUsNZ66rcfyKB8vznz8uU6hIh1aFiusECc/2gFUqFXnW
Y1iHuFGmjmx9f+BY4bn0dsAkNKNZn2VSuJhEndi6AYaWI52ifP8SqNx9To9ZRGcskZEuDsQ1eMRY
r2QgNHpu1S2Rn1+YhrYjBTCO87SUex9Moodla9fnyK0g8mQM7Rix4sbghr4vEzbL9rv76d5SJjUQ
bqUp9HeEn13OgBfnZq++haLCw2UA5hR/SaJrhcHHxlkhZZfRocIdtJgz3V4iD89A+g+6hFOT8knU
BBgbrws579ceRhPOUMfe2IDsRRg/ndQwsEPej+8EMwJnuo+nFn0El1imGhKigz7aff8UbNeH+b0j
07zOp96zupAc6kENV1xuv+dmav85luKODrA6j0wABEnAg5P/uRtxx5ONhcfJdw/7g7XEIosFYHs5
/6YF1dJ5bMib5v+8wVsLNsd2QS+3W7rhqfn+hTgiPX/soNS41HAc1+6wbbTPaWVqFOQJXWYQTVYA
zgEYe2bm9sR1sMOevG+j7cS9n7ot6n1wjghRC9wONKOnKwtgwrQxISlC/CUs/qsNnEwkIY0ZE50l
sgUZTqX2cIjmNnxzrQ4vnHvn1YyhWKqexAp/s6ZKPMcFCMQyy3I0hkaslV4qY2xk3/ugsl/IQhYD
Tp4wWaMdZl03RYYncgEzd3yWOj6p2PwKul2okF1s7OFMBU0RIRGzfwTPoMKiCxhq6fxUeVyEnxNR
7H+3AqIb3EJvUlfQPL03WhlCpj3vez6FWDFxR3IsohpcN6+X/grqnyr8b6li49QGadvrKLy5Lziq
0vZPnBLl9TnQ0Sc5gbtp7FqBsbxiRGe/WGxZpHVmf6+TvzqNsAMEU6RLA2rkMccOEfGpC100an3F
AI9U5ewIaC7gsytmS7y7reY5T/uoiJ2IQCHp9O9tx7hTZWDhqReKyt6MLJcc4f04V9lhMnL6KFr/
Ue5zwDyKQX/9p+m3JqMvM8ZgtE4WDKGx0tl0xkufLnorB95Ot6w/vWYD0xJw+YeaI4CrGEKAz7yz
UoOsJ4ZWWKAwClbZJCIFglG71uk8u2z3+BcgowlJA6se1zXZ8phJr0K+muwLSFrvaQGEpcd+Kg4O
hILfj6Mv2oWtpqOjH102n42sgRh682DdHioRcFUrf76bZhDFdGKqrda9n/ioTUgyLPZSH+VumJv0
wJiyghV6KPT7NbWmtAsJS3Y+dkooITzqXYxAfoBcZYsdM38ifWs0/0FuKSFnxYfaBwzbxLM29Rnp
3eqEg29lV6AfxGnL3zBKRunHuxPuzjQU6fWJpoWyLSkkwZ5x+5RiZiP5oMGVf2ptx3P6KLQwPP8U
r70xyR3v9wq7QSGtqFjXFw85ZZWTr6gpp9LneQsEqfAHiJ7+6gxZM1OGt7VmHEVyJwT9tUB4ztsi
w8qMFX9MPwHCqWyCAXRHT8pqoBb4SC2PHdAFAFm298T04Vh2AXrdUACqo7ctQ0E41/RLlcQQve5M
XeAJ3ch4qcurwlZQ5WzhWAhGLnoSKCGQoCkrsJaU2NQ5gLaqkzrtx3zGZyWagAPvDqfoRzprR4OM
T3jOOhJiVTrT3cDteg2PgEvbq6mRBDw52VYHID/w+HaLrjG5wwIH9YQiPGCyXBoBCZZ14iNNe3cb
2FbWtsLeDqA2DeV1lon7qOMe3GumVocm+/bYkNmugP8JJR41i8L1FoIMDYaVoe8FMz2WH2CM4h01
lbytlIwqASSoilm8HAiiHY/rKJIUuQl/tTy6v4YMs/1oMFwfHFzHWA/Z6hk0EAfx2YSOtDncMo67
mLIgDH4ndRkhViKgow8/QmN6dBZ/mGFz5JRKrgqkje0oe+KCNHTKlDPTMJ7gY/I8NUVLhkiVnD7e
5eGrZdlL0Xa6YwCCbI8DvYoO5A3gbTxf2V2Wei7g1Bn+w2UIKVnyEpwu1bHH4ofHwKcO6cdSIRxx
nh3f+R1M0fKPjXQGT7sCHyy0crxXLq5hNYQylgw2DS0pP4pF6AXGt9LRZdDaV9pMoELpid4K/Y42
yrscuoAnEIi5XqGvqqJ8tDOaZ52C2mhuNmBD1u0eroo6tjvvwlnqofRMwjsm7Q7gl71XpMtUWMxK
sujwgqLxtzjDvn9Pag1mauf8P20hwW3rBHyLfRTbZtXXM3XZILcsItYAN7NQFcVcOu0qTW7jE2k8
HwcFl6VZgvssyJ3FGsUbikzrLFPsdh3anEwPUVvE+PQWNxHRysokhInpO/ZdVCabKwhfnbcqvkKV
oYHNkgWT/Ku2nOHWapUzmWlJsiuAIB4HgJtMheX1Bsm2pGkqyJrxc3NwbyFqn2ZW5dGh8ISrF63c
aDq38D0jobUUk9qXpGixutC0zhHy1ILcvppqUn7C7J+YiYp5032j7VkHs5TqAxlE/ftMmBSJPN2n
jzN0Fq2ojo7ZsLmqt92MHPK0U/FtDWTUVKQNkPDlE1qB1S0wvkCtgZAzPpfj45T3DYprI67oDvNN
6lQyH9ZMa6RBmBFiThzFjXNY+zSqxOC+fEljuelqWrF1BjDR3Tr0ybMneK3jNo7alAcz9x4brStn
AJrXMXjeaPQpL+I9mPJSro27INTf8Ag8EYKORPvgjc4pkEzoU1oIs04/bf/RN2XB61iv7MzfsTKg
eFvd5GyqnkkrdUWOg55/MHnU1nooiPPeKwgfcMaXUWfPcKdvrwQ6hAefaQwn6t7zW8dnJMAFaCtO
vidM/v0CUwlnhHkjsu08W+1G6Q3qBWyqYbREtMUs5iUXoBq0JCzFEbor8BR/v85+HiOuKMbPANGl
mpH026XSlL8A5GS5IDrsGI17kMY58lNzalDtO7x1h3vFrtIetWXY78/hTewTOtrTod6XcO72vefD
/l8Wuua6p6uhaSCrIBOLPwRP/BzqVjtwCkT2Do5Wx4q5chVodj592NwY5xiwNdM1CMnk4p3yEUBF
6xSL66d5WAQvMEuzEmQqvtX7BDmx1YV9I/QH4AHD5bRLCqpCmUyHb0+QkosINNjrv9UWMe/GJTl/
IE+bo3EZ2ueI5gd9OmhsBuqG84lt8Os4x5n/UACKC4+sJlabh1eGKwZFazHnUZkHuEkYHNmFQlNu
+/C6d4wQRrwHGn9RlMs70M7z4/DMik57x/Me1zYdj2aNZPd8vZKESMiQZZTL7AAa+S3+CrD82eZt
fh7FPZmUfupghbWhoYmzLbPRvIc6i37CHRoyk0cfSh/YXt6QiOzpLpRKMvN0g+xEcNIzyJl8LZL1
k6viTIDT9AIcPEuk8TSwkgfWR6vHNMYTWVj3138WwKFgdPKrHBQRV/LYERExtf793AMsL9fc3Ukj
Tlfo3fRo9zn5eap3n6Dmf+q1FcWGRNrVx1eRD4lYLMTEP4J6tZ3UJmWHK9tDqMCWgUbQnT7N/rOI
cZ/OTDACFsCcKAbWx40zssOi6uB2LT3O14I0yvASDXCsIUVcyZZRc/i+nxCr99n/MvQFDK4Lfp0D
77Al89JGtIVmfwhD4NyKzvFc3OM/pEKQKK1Lt7ANSYRx3nsKD94PlpIlLZoLwaRKBSLKP9RDDPYN
FlAFE8qiCwf2p3gQM3pSFLwrTIST1I0Hkgwbx7/rzkIosaimYTnHmMSWBJgqr7F5/LRWFsnPUodF
4rikz1lsTILCqNL2BHIKf5NjruupVMi3fG8EAJO2G/F7w90GMQmreqwg7mwZa+XNl2YekhsYjkmv
DA4GL30szM+PQ1xtHUEjuehBxl915tgELhUX7xGvSGVIHcWaf3wwO18JpbbCUEcpXi9JK6dUtvta
HuZge0ItG+jg0CJPpSsHMm31n7OJC9HBxPTAOJdV2zTblL+NKvY1v8FeXflHko3tV8h/kCsDU6Un
pRr9BVnVXg65IJOD+JOK22LABCNvr/eoU9zqoaeszKAd5tPJvWlqRIMYKlYFy7/0V+KxfsNwvdvF
E7MAZpnSd4qBwpJv+WtP5zLRO39A1Imf65hxEE7Q3j9dOFhP3vDJRjfbkpD3860oxfvPMglklEku
y5NT7fFTHTIb50QYiIMlmA/YJsfhv4sL5mhM0PbNZ0YZevH8hlHxzjzWJOykkfK5oPyobX3CyHP/
22QzirtPEzqWhsRpzm7Lkit5eQj9kPRU3kpz4EhDirUc7OqQ9x6dBOuhrp3CAlh5ifJGn64WKU4U
t2/Ron0gghAnAQIqmc0P+FxQBi/BT9UEdzzINP6tY/p3gfCEQ787zi+Xk43pz9OWLl3cF1Q806H8
2OFQakU+lZee/6s0gFVayZcEzHJ094wcwkncf6SLtdM/6EgCY3lwOAHxRq/Bz3c0vnjJPtMvuZcG
ZvNWV4zKoif5AT8DdCM7U3XTcWXc56kxA8S6E5o5EFKkGq1IwurLeIabwsFD4NsE4PYLCx1hlFH2
S19BpBzBezFU/a3pr43MXUBFv6CBGfAaYQ7uVK/B61+lqw+7Z8wIrNyE8y0iQwU5HSziXqUm9XlF
48aTUZg1/MAsQUm/PltsVAHqTPrmc4tFAWN4xKTnhNZX2h5rygHBYlU8rRFnWLPtA7wsh0MbjzQ/
yy8DLXR+WYT02fAeuk6A8sEyLgpmtyujDAmcisNABeOflZNJDM5Dh9QKQn2MXTT67oC4I9Vrcr7e
z6Ii5ssUoaFDqGTje5U52ufMWM2AmknT3LusFgX4ww/eeJAONLlZwJgoJ456aOOYs0g3uZMde/P1
q3rtUsfqP15kAYjpURYiv12aKE0bk/g+Szd5/fhCG0/BbiWmLdPlA0GzPuoPtaBszVlv4hfTIc52
TCY63nwvS+21a4ZpZ7u67uPRifeQnr1imP/tLszYk0zPfREjd78GPOlpWoTSmcRrd5KRZVI29EVw
5VRLD0BOZBDoCp9m6pWIWzE/TmaXZSYp/TP/sOvnDp8HFsFLhg3BeYzurPK+C8EF945wXaeSny0T
xoBZTr+ZaYIeYROM78BzuLKUcgsk8VHisnZZ7uANarXGXUnAedgbRIQDIeTmkyHL7ycWJkkXiJ1M
T8km1sAGnqGr2XpqJOUBpe2YhC57Fj1AP7k/s5VB1JTlkA23S8zVC24ncu2LOCrHYe3SKCGcovx2
JhA9st8dLiMj3V2rQZf0UZC53tJtWcEsYAwJCqjEzFkxw7mcpuyYUqbcyTUItTVk6iAXu3US7had
fKluzO4odYKc/gcDfIE89sZN3sfLObadoGUW54dlXUe3jodTDotl5I7xh06bZv6RiKqdcZAJRpRL
WnaunP9jK9V+WUVpA7uerVdBYprqPqi0vhgs30KHilZ3slprNZibqgm6GMtbA60e06suniOJ81/l
6PAtniXKkOFyvlIsu0GGX+yBAZhXRrrI+Uyf0L90Jm+dRW8SzCTnrM9TDE1PqsJMyA3tdoarsxX4
UkZK+hY4B1HgHIFy4OFOUwE+wv2Zd6KvC18Sf0RcOQfWMnjQFoN/EUJoo1gOomfCVP5JzoDgciJp
24FoAQYMkiUoTtlgpBNrSOKs+n6CdGimLSkQ9TZZ8An2lX+BMzHc/2lK4SqRP2pinvYYW+yYulXI
nX5wF+u/l2JFlDhePs7yvkoI1KWfX7IonY4kkqklhsffahb7l4r3gmCr5sZI50ClaWa7WdYT05I+
O9ffjITdWN9bdgiyEjbA5Dl8EA5U5xpLn8dEAI03xljMo/RgKYgvbwEsTXppCpIlszVphvRvEnFK
2VM/UtvMJRumnF4+9bkyt3Kf6M+YqTPVZl7gvBg2XJ1rK/6D/m9zBWo2mbNTs5uwlwSz/iUIPMn3
lZNEEkzoB57oN3bjNG2izW/zLVgH0b3dyOih+PUqfDv8p+8fOBlYs3jsEhX1h2QJXKbh/K8sYLVp
lDUpYP7u4EaNHrYPstV2wicqYr3xGLEaFc6iUbaSdVLD72zrt/BiXHy32W06MR/QFrZ9q4Vl5Ftl
9s/QxgyvPpDjx++AUpVcPr/KPIKH3Ua5RoUOEZKIyq6nmoOZYfJwWolF6wChdw5vCfmwYf/fbJwY
3cm8EmvkFuM5b+nFC9fCeLqasud4xxSk0o90XuZlY6dQK8jGatEvTzWjSoL4RVwgFv/qT3m1QINK
G4oW2WX9PUEhRGDd4UNvSCgmYiKG1stJQ7lmW7Fum1iVXRBAAWAB2kgXFTjrAWH864TM/LNC5v+8
1/NL8DNmBXo8X9jP33u2jxQAGNzI3QqAQNVs8gm9tEbX43R8ZZWAXbIMCO/58cuCZlDLVC+R11jE
NRfVc90y2Pk5YaWlhXlzGoIJq1WUC8PyItcZ0vQ6xYJ3F7rOpjNSbHbIkBjeK6zDCWE5C4Fgxb70
eyYVywaI5JP0RFh7Ly9G4J63ba5ZIxDX8i+mjmW3hBQJVvLFfM7tf8GUBL8gRH/g9ih94gDjAWQJ
1rKvO2+vHabJ0IbkjZFfOOTpP7LvzWj/eH7dldf/EQ0AD9CIuvy3SH6oHv10wLku7EzwInKUQ0Qh
QMEfIY44PGFaz6myPntr4Jh9GPqK1EAXcPrAfzqFBdwTpRw4Cy1Pc45cOHCkssyBAOU5dY49/FjF
kxLSYVX2DzfLBhPXogp9KViiRl5ftmqBhgxisbGnAL7xNEWiPbISHhk5AA5YBawovs6lIUIwJBPO
vSjpT0XtcBb/5uvD69aNEIgJ4vnhC0NrPbNy33MVxtJMcDrZ+fS9SqBqZlWfughtha4LEkiUbi9k
B8xZuvOqnR+tKCv6RMPqA1Uv6NerSe+LvYu2rYYXizA4KQBGCwAFy4K/XL4Ej2FwfRr24GsOofbj
w1rkybbmVZ5JuY67Erz6yAPm4ka6szylWVx2NS9zSTZvqjanhYxczZsBOcL5bj8a3z4EqyUzuTSW
TVbo0yZOpdcDkBhX2nvIkTojOEBxsindtH2Lkeh/WHxM1kxFclyRMHOoqUr0BlQqjyzx2SJQYk/+
/BDQybkoSoQ6F7JWdof/UlueIek8hUKvg4JAO8m7MfgFKDo13XIeyRKtQuPHtA47/Zok1EA+ZXqZ
Ua1kbj3nPfUD0b+zOt0hZxhbEk1v90N4AKTGOsH7wPtNXcdDLxUA8gUHFTqW8V5W0rWfZn32+ePp
NQEvnnQGzgjXmWybA0SRMAYP0E6EUuJislqZa1xs4yJDtMAhRRgtZwlSxgGt8HZ/dwAWEv11QFwi
v29A0ihYDSlwyJ9PWs7vhdiWae362shdmdFUvAUDCCPFEPdYjzximXGWuMcBe1pUujS1yCctfvkJ
kMIA400/+mgEMPiabuV4E+1VEje6usKFnCgKaNZ3R2VXB0gP2z8vB8QU2duZ7mPgpxN3t+g8I6/u
lo/3zDH1Q2mx7DooKjdWr5EJSanYr8EpXnyNIJZBzMzbaMYC5nRPxX/RwPCDGiWgfUgIPmuf+oan
gYNeWXsjg4/r1dOfOPjDQBCUlIEJZeolPCHL5LvxnHRNj7p+ABhoYgcEJY5FSJWSKSrcYbYBaGeU
UKEAE3RkedDaZkJl/bRGJ1L+q6hKwzSQDiFlsFOmWRCyKb/5IPmBhyJrKRaypxPV5p9OTmhjJg6W
PAKrCurMulYQ93f0JRvUwpE9qMcWnBV7zfJ8IApj2g40Gfc8oyLz7CY1I+CekSHrZ2GrOO5lseh0
S23ekxmqwDAd5adVitN0acrS6q3Z5GkiSzkAKfq/8LdgD74YTiw04F01sGuFxAAS9QvLmj5fCDV4
P1wnaUI8qbHOS+/rCdhs3KLQymcsLA2zDrUZnTBjusaXKA6DTygzMYVOu48P3O+Lt1eBEci0nNIO
qHtJE5AHGla7DVz/8qNGxWXnlQ6Wz8rShjIxIEN0AZl/lc1WzpJ10xzGJLe3mHd9+ZMBqyJqbVG/
+B79qIrjt7UyOYjM9L1wFqfz8L4mYiCXo4IOqvlgifOwqJlhjtF51hz1egKb8A0saPBoxpWDBq0N
uI4itj7NNVCzWGMUF3+Dz9HVqJ7aaboW3KJJA43WL/WceJD7YnicGrud+h8ni5laafMaYOot6Tzo
xc+2BI8CHJdBaD/DadKowFTIMWjCwBgVpLMe2IDN9hOarcuKaqe5/wXgbiQ5TcfVRPBPbD9kSxkv
kSZf0RvWOsR44wClMB38VR+tBbf8NLc9LT04M0s9jD1gKD3/XUmKyA9Aji/BtHkDz+jT9IS7Nmlh
5GTZNZUNfXs1N5SBULNurCK4xdZ3iHKwL6Ctr/uzwuiUqlkzbAbvgsAUl+aEcZT/2ECE0WSRUXVd
BYO3gvzNMPaSrIbzyfBbdrfLe3sLo8xsW9R3jJXR5Tlr3pCsVAvkWpqY0kvjfpz5bwkWcS/4BwIQ
MkhwYfrQGjEDqmXPD5gyyH3RG2Vz//O1uLdTeK3eYY31MwkYzVLuh44JVoktshFceD8wjVQzplGc
11fdIm5T/pF8B6Ku9g2vBJAEbrpmvZjIEzLS5dKLGJsa2RV2tB4nHtraU/8GMsyVFm+VGev8tDLM
fVxFF/dUlUnS38LLZkwVsLKxnTZ2hKhFg4G0cNN0JyJxSS0/OYkID+740K6eqQ8u5/OH6K/83/xM
UUkzs4QjIeLChQig65A5sdYO3YlggaHHthO7ayX5hZJvTyYKaBykncDxDZhwQtJgRP4gLkGzVPGS
VpaUqjyKMJTIJ6MwC1HqCSSvZnkM2ZDp2T209Sm3Sv6pHNGPZIUNGY6Lo9ovlZzPwHMd+qo6Hcnl
6Ta06ulDAOpVmUvFURHqz6FWFMua/OUNerGscrfq+vXODuMl3OFGmeZCHO1Q5lWjl02nGLrz1OBU
ktERk0iROMmtFXbCI8ZFUwu0m/UPEHb9t8xxlKMVM6l6+SXxxgHOBBas0xG3VhPX78gwxCxwFqUk
LcxX4E+x2YyM0nAAimI0xuUvB5bcYZf6HYeFHXz5/JCqOwIPvVV7B1MXLDo5y44xK6w3Rz3wD2FR
Ws12pSETan8DciX2Lzh4WW+ucHfCLTdrgXH7ajMmqt/s0MeXTVWFTGEDZrjrxoNCAIUzU62fVg9u
IRH9uL7YWdIUEJ9VCNGss+7ALoLPorq4pmKtQY3ve2uU48TFI7vZ7uuNS9wMEsYkBA1T2dBKuWiT
BF0cNyPxUF+YMnnlULnzWYGTrH0iN+PGpszmhTE4b8qRXzIC5rJAZpWVX0zdIbNx0gA6774rXrRN
W/pzCMFBTZcZRfG4pT97mqs74IW/nywt/NJkYMYvw0fnzfeA7vP0BVwF8JNre7xEx4G43dUN1yN5
+jrBtiJnoG/AoCe330k78g7ZsR1qs9QpnkK917DdqjiqGDtnLD4IzcIrYOYX2EFXgLrCW2X8ZkWo
qK4b6OIBk7Wim2d92ye2Vakia9ZWQLlN6T5choY/hvUoXNWQH/U2SlhhONtk29cnM6MO4eblpbr/
yk3uocLYrrPJIdRLBih32zkcoOz6XxcYmVyOvO9jYczkBB4KpJgBtpDEcl9mU308FvgL/rXlLR+M
Fyz1gH/EZ1sIcOt6LDujvyIaHIrgHeSiT06l2tENsGEb3rLp6hzT6AAeLF4FxYXUzb+qaYKtYOVx
Vs27G5pVfTc9/B+1iLwE/GODBNaF6RfMf2k8W9fhasD9yjMkla/4OKyGPbcoQusPodp7jf5egKX1
p338/Vu4hYJ++3IMKysD0Llp9jWd8YxHO7t2/ZtLd9RY3jT3wxM5de6EY1/7URPXof8aUpt+hRMQ
PqEagrcRFtyMQqfoFj8OyGpBk6D1VDs862XBvZEdCRoGYqAtdKGRGZWe4Vk0A+260sExw/zdOsp2
8w3nF3BsNYsXj9NzYAjSYrpzlJT5EiaYi9AfyjpKIeFno6zXh/Nsa8wdy37x46MLw1ePBNqvZTaJ
rb9U26mBIzB+Xz9dPG1y32n8hnM0Iq0rXsiHWX8SSPjD9/HjCet/5WD7h0cim0FJCyS69ZpqsDjX
D1Q2d27rQxrxn9NX9KWGdEm2Z3zVKjYYmJ9Oh33GNsAL6GlrtN4FotqLs1O5GA3Lo0GdLYalJmDD
rdvTR+j6zGocxt0C82FJgfUt6K5O9kVMcK8ZZ1vz0wlfQnc+H75go8kL+N7fED3M5Vahsnk9qbz7
qOy4clv+UwYJE5toXg48t4jHqPyGX8PqIRMHWaZ/fBMVJO4ZVrONZiWzxBm2AR5EnFWidjXMcR7L
0OsUf9P0Z99vfSjkSp6IKL7G87upCRv/Ymg6pxkC5rlDqFn0iOFn3sxOPyulSW9DngeR/0BC6CMR
WkJkxyqTvLgvNbTPBmfLQMHb5N0Z8Ur+WadIkh6S8mROm6yhBuLLCD1TWpLYXAehlg4Nkb7KR4lZ
qHhcSxTRRkoUIbbzbO8l/0EgUzhIoyBXyk1smfumHAq5gu0EYDG5kSu7r1KZ941xxsGk3MtRNF8d
QIrWEq1u42ssauJndc6qb3bZsmvPpfwcWk7otYSz4lRvGV3dGh+GlEkVechKR1R23/XPwlGFoqsa
8Z6uPkL15m7MiXnsxcsLwUtx3Ku27cGM4Vnqegk9iM1gBcEp8bsyMt3feNcIhfZSIZoXuWCSRFBT
qBGwbmbCxE4TfXbG+yaSD23oZ/1lb6rrHoNDsAY4KfuMdBSZBkBTr2QUSTpkz8758TnMUelkQSH0
TyhWD6bSaCL+KjV+nPrkza/k/k8WSGMizmxm5uPmPGjbHszT81eBWtrHm484expt9jAKtoRVSyba
oJhnfyIyncV6I9MIJsj8wRvRCDDS9IAgC+so2Z2UGuDy8l6i/BFCVBxTOBZeI9aXRrriMzAPPTZC
W/kXzUNmnnAhAG0xxRTFi0QLNa9y+spppfoxokwE3Jh6OpZrwWVGt6LXul69CGaoSnfmJfOJ1SUd
oksj6g2tf2KktMrcZQrnHprkBMUn4nqIDce8JMznKM4QQUUsfcrSDciBhQ/GZ7kU0GAdJ3aWFLDv
+bcd6Y5dNnm1N+7ZGN+v3SKA2wmqUhgfFRItJzqCIxvv4Y5ZobTXW0QqSXi9CHzrEkYbWjSySkao
4BEnrYmaVybHW433l04Bgfyow1ouB/9N6CRBZqR7GoEMkAqsmrIczVOMIsMzor2/j+bxx6pLktMh
C9yhMvkPDnDdECRzXBPdlqndjV188FtjjQrr2cl4QhuXHJDIctzAgzOgs65D9kYv2CUtqiK9xFse
TVWRcBWk141kTGH7vmNQbh+Im3/UsBuEjI2pu1wOQhTsjRz3touFWXzfSWXm2RzFM24VFXbtSu/H
5twp+oCuQiwOen0PHxy5qWMNaby1ytqlqYjyxDnYYvKvFTugaut4bB7M285+7IExVfWe+jOyALBI
wv0Q0YWZvSxw1OQe0+nLxVZ9vmK97taV06drQTuZy7gTwMO+zV+bAGozNwKWi2JbuqBeXwD7P56W
Ghgj5VGgpTifLk6M4LrQHVWiEUrbIvdz1Xr4l+Iq13qzd7Hj/SlD2PShVIIJwcrKw+F/R0sVjbzy
1LgFEJRZCOGokKx0PXs0ILNkdfG7ugj9sHsubYVZ7LZQ3WudF999HI6FqPW/T5lCaJyvOhI3ajjs
NKddjXzKnPN+37oh6Yf5GUDYciMIziONxHvJYOHVviNyjNHlYLs97CMVAV1bMnVH4Js2tEqOAiBk
K/CabrX+h2iBCgv6J7aIigQmjJWBeqme1WIverOQskkTgy0ShkP7Gg6rDS/DjjopLtvgbVj2/f4I
ldyiyKAbEs6KtwlLZxsuXowss49Y1J//pSlx/KHP5ufbb3r4rHBt+MvGBY1iJAR5xH+73pqgBu7T
4fSvNcu3R4597EbQ7ZrCMYmiw0d2z2CJDR5PpCtO2ql5MLTm/5Pvz/oZ4XvbsmcYBqNy9mtyWZ31
3hHn2ls2nCMLCGefASGu0In1hlRWnPFg90A5+s0YzbbB1l+W64GZFJHSVESN9NvOU5f2651t0VZG
aUjrFF4Xk24dr1yCh6zzuzBYJrhhXfBm8C4kz8nc334C1Divgwki59hzRk1/s2oljXKC5Cdm4Mbp
ZBYwMXhNzTmQjPnYZKSSEB0AYUg1smiERxi85ashuxzwTzRlzHrCdWc/D27cnF0WfpeDjJNCIS9J
HH0d57oL3AokzxsRrGGkg+haM4uXYzwjJTwMLeQu2tziW30Cf8lsumiMmYYHSVxDCiY42MSEOiOJ
8pR9GXhlzSrljUjmniUNvOqALGUoylKDR+dMWpZ/c7drD34pFC7lEFc2+sK0qpTh5ERlxPg3+brI
7n3XoEGh/SKh7CCNZ38awCgfQEEgeuMH5aXlAYdSm7lW2zGeKE15Y53o/Ic9jtvxAWVIczIi+5wF
JzclyuvH1pLhN1L5IIzLORZcMBKgcVkDZzVNdNhwPrXKGb3bPqgvSYTcwuta257L/5S2Xb8dYhUE
nUeRru3iCQo3uYtpgJWxZRvgEGTfAu7E1dMnAyAIWPUV4g8XBy+cd5ItK8G56fwlfE+B3OhsHIwC
4paRcIzNpUQ8FGbSFIFOqaQXMoPusqeolgTco+TJtiejVGcO1YNQ9+vB1SHdTzZ8nVfZql2PEl2F
MGFMCbF46Z7FMzUcCYJ04RcdPVxg3aTc9N7ZxaSzJdCHGrJpB//xAr/u4/+Ibp8g3d/IBro125LM
JuTEem0Abpl2s0zLl4UXMKZYZF1cY5EEzK9Pm/vLFki+VfoKGAywOH1CNnP2leGr2cgi6kX5QK6K
iy6000wBUN3yqDAGVaK8j6WtF7wTDU6EME5/8/wX3Z2aa4Gz7yhwjcHZjc1cz3UYCbK+FKHl/8tk
4Zg6R9shOT8JeOnvm9OcrtuKjzMhzS0Cmd6zGXNAkHe3IeyQ/G26G8pZum+wh2OXfCYxn5ZqbvGL
qj5NZ4geRtywqHG6v8BDcB43lN7olTk4L1ll/8TGogYNkt98q3IqLJ9ot70JuamX83HTFXbHE5YY
cwMERKDjJsqdgfuJdSF+o0gFCNVnIaUUjXN8YpuR6SYJn6i8QS7G2M/9/JzRuXnPuugCmugdgP8J
ke8c10wvEfQp+kP72MABaQpqg4HJTFnTw8jDg6osSSDDWTQOdBOgKrd9nToDx8gKc9RX5vhFO1jm
bdJTMabF5ixcql9RDPB/K/yeZUenKib5hdFJFdIt/FaUmGilORfKIu069mC4kRj69VTzNCH5J9qW
U+MA37B3GjAVmGtVcg0ecxmtMYnyEweXTxzpQ04SqoDWWRMQF03vOY9oMn3WrlM0/FM8OffcCGye
rAJMY3AzdNmdgEPiH2gbImELUrjf0Z3uzDkRbEig5xCwDA9T+apEP+ZQOCG6PtCqhYNREGk5RcjX
j7kwdYifHod1iNEom9VnDEXI9bigtE1GInmH89SFUBFmDEFRrcHwDmnpsleBArC3l7z/9YvP4urM
oEl9MSUJ2KsvUPjCP3c1RMdTQ/S/BeeMWaaKGKHBic9rz1FGqSAcr5F7514mb+NINAvOi5d3VQn8
qNcdy5D9Eh9CMmUZ4F9dGs6MEI8fNNi+ATKdcUdpy72Kth7N9HkADq0Bi40/w682tg8Hh43THW70
45DyIvTd5frd2n34ytGoI/Ci78Go91kUGRsqruGFNoGjAoy3j2bUs9gT4g15S0NX+/mKPXPBIt9o
KAhWVitoyjXCoaE9a9yziLgDrUnSO+5BROwK3tTjntGX+NbgEvp1y8jQLWJSVmfCTd/T8mTxT55b
+Xh5dVdMXX5tz++3wUn9OqjYZ5icg1eV68D6h8eRqWbd6CCU+pYhJ3yyYzwrMtOVCChHloEdMypr
N1God1G9MVVNtMVgEow66uBnEi+uHhNaPqJhmo0/WcgS1CsK9xY/idDrimlHodM6HigiAw852NTS
17SwQo0XabtUxknlgc1z9H/xKjgLZOTV5eJiWA04zEVe2bO/21+GF9ZbHHhsK+ZWKv4s0Ji9zsZg
3tKrFhR7AeEZuosFX5Qrx21iuR9SLwgvFK0hK560H9zLvJYmXyHswUlIZh5YIMQGOE17tUmuQzGm
Vx9CsdJhUJgAbvjx3CWS476rGs8h9DHov2GnPsqMfrDBnSZrRm4YrC31jKtCxepcQWUfvRmOVKcO
eHMQcMm540eaHJzratSOHlhYb0OUmpVJ+QpD/aGMjRzpk0tbjvtF3w3A5s5RnQpcCDvXT8XqUcOG
RkY166aV540BDfSUp9h9lcVqXy99UrOZd/jcMW6YriWfo3xgPU0i+TJfFM+rPsDfbwhxINAF0Pdj
TtqwCCWd3OfuBJlS2/5TwYsZpbTwEA3ceJ9Hd6ISljpkQHDmXPxfOhvC/4I/Ic+qNwZLM9ZO2l0a
VCp4xn8SKUzvygK2rq2nq2gIfVFzz0E9Lh/GSE3Styb0la+9t+95lyyRihlpvgavp5Tj1ihvn50D
LbfAljwaTPWja1Vhbc6z+cmBjEZxv3/AzFVYqGu4WqkB4yBSXs1jaKcVxbrx4wyhO9+ms4BeRneX
4Dz0DGoi9DGjSGzAb9PKmrzxbIm8Ve1RXm7K+6VGiBZzG1b2gSCtBcJOUaY18siFOlUl5ehhkqDc
ph26tMBYhnBDiwqE0/qfOfZPF8/+omxy/l8S3+qQH9LOJqixu6RL1O+6u5I6Mh/Sh+Vg0boZrxBX
s1AYiOS/plKk9qa5YaNTI/zFji9XwyT5ZtyjdDig0PtKkhhkEKvK1FYA2SdA+5thdQ9kZKC7+RH3
EMXCYSCk2/w7GNfB8WhK8jDhmfh15imjacUNyy9AVHZNL+fgRame87pZe8BAr7fbDqvh2cbLaFh1
j/0ZU+yP5N/rjayvRyLStI+gDUbyheidNlfKAFXJB/QDKEmn12HaYs+rmYJQEzEoau0+2ABiHEhf
nxVn1zpvI9UrpUjh4hYBK8Cuu6oJmfHXQ37sA51UpfaUVvlhr46jSwFph25KEHN44uCpKyvB78uc
1mQm4tHo1TRVl2sFqtlpSdLd/HVehh6yy8gxf+ToJJPhuOG7zTEtwR9WG1uFFfiIjlQwDy1f7kaz
kpkTXQn03kFDqboM9tO2wr3l3xcYU1eeA58Apn0pv1SBNO9jDAaYKuvq7C4fesvaiZXa5AKUhnZv
B4Rzf3rmLyEel3/puzGtHbVca/NeeKL/rb6nI8P5+Tcqzf8QoAzli8KAFcsC7db4ibuhLJSwlUGJ
9SPv2dSA23MIXWcQdGbFgxas3MZSQWZLFTfRjvRyWiksOiDl3Wh2f7mR1tZ3PRt9toICTE4xEA4G
22uXBryEWSQg77/+FCRQICGPAML5lBU/gR6CRnHcTWBgNcjv7NC7M+GV9wljO4qhkMpLS1D9AO49
CGdZNURhOj1OIHGjkjYDgsNgX2V3/KZPVnn5z/mXJJ1pksT2HLteHMM0VNzshhsq9ev0OJFH/Zep
UOcJFQ8rpgHQUAnq/B4DqbsIDM72O1InUCAbVATIA5CDy3rdiz+nmelZFS6QpDMsBRUhgIIyxMPl
0LgO6IMlnrSUhqs7M562jpSavdWX6RbAybppjoeDY8F5z9iNa2ux3ylBD+kI7ai6NJd7/pxSfaTh
oPkQkn23B7L6t+EXQ7+PSc3PJcQYO3AivVIpuHhoF7dDRNzEECtD5p5ZIQrOe8D/gVjD9yB3npa2
3/GG7j7I5Gy/v6etQfzR1DXc0tMWR3evTNqCSz1giZ+HywjYgNlf1TRcHxi7TwasUJY+lBPIJPiX
jwKL2Srq6vBq5eJIEnJSOdLDb4QsZ8LO8ReZOsW1O3Bqkcijc9kSZ9ULF3LK7+5+y09IHHbcMxAK
fHX5mytkgOgI64EVKk/f1Ctd9scEBzAv2qBy6nohrrsRGJX2jNeEdzSxdMTjD/yP1T9mPi34BuYO
Ncbu+mN5NKchjhq9GESOKEOfWASoU/fByU63YnqPEvekuxVb19G0jBkXnjlVsDuaT6dfeh02zhjG
YR2qKiYdPFFoyFb55DTAej4l3xzXBopB3ZgvahS7tDwM88SEThH9wIObuiDDszF38b1ygzNAbL4Y
pwHhvSnGlH8TcRyDqgnN3n0ybqRhSOiZXzsTKPoRd6REy6QC4kkAYDS27JwRKjJiPBFEiOWzYDot
RefCv/PaZoAHwzExkTymRX9zOlC/DlgspgFXXtozjDNeM0hdy5tuzCm95s+tI+mmoI4LBtBaAXzO
Mu3CUhI0OLZfa7/YL7aHwElDeaEoPhYF8fp/svuih3q6NYhhVJStrBmCFMWyRbrMdxT9AgtnNu9f
UEm4M+3FjBN1I7Md7kLicywzAp10PQCXQ0aVqFQWI2hkdOw9Pen12MAlXcU7RjYZSC9lWQlGQ1gG
6mmZFaYz6jHiwe43vd2e0aBAqxIn8agooa03Uds6UmkJxHWFGgLjy6d2sQW68BBLwWO0bZZmNXUv
/hcFAZ9Lix9oI0Dt+RkR7Q/g3ACerZmMLWXzcNWJn+nUzh4bt0i9cfx9D6m5NvjHPnKOgqAGCR3Q
t7n4NiU5DOG1PF1jBe4zv3sNdb9eUwyxT/dlpuow0ftbDl6/0NdOZiIoSJIYzni6jl91Gc8Z7AD5
hBmD2hROBZTghW4TlavhRLueFyHii9kf1NH5QS6Rh4EAIoIPMEIQotZ6fYrKY4XxcCNlRkZBiEcR
eMbu4BDBvkWiEjNaygo5f0NPxnqvaTAATqCQ6vXaFB8eh1dzBubotOoOkAt1UmiNJkmvzj6E/C1j
Knufa/vDxTu3BPh/97Gp5BVe7UPG/Ra4+PpovHo99MUhHpuSGGUbeMRBVycT0Wwpm1H9DZp5gPIQ
QO1GON8sUc6xCmPqLwdOrNwrwJsCYdCH04IDDJUAVHb3rBVg3KmNLVSdcQi7QrlbHvrvSATIAWkq
Qm4DkDEdmIRqvUR70bUCWTluIezCBRlAzbavXfgH9MnN3xQS9UvU7/uLXLIZSIkfeOYqxGtc5f+F
BdIa+7jJN7S+bTtSLUPeLh3FfnSsKIlG4p/WFiUjJ8duojZk1UjhVRIgd9dEHxQWVhx/HzR/4ygY
q574wbHa0JuklCZxd1qQeo8tUXBBmeAjWFvAR8jvedA34S7zxnySxMV7XoB8ctpJ/crTXddMRRfO
zn8w+K6hqrWkrCbFzuTSxwwldFr2/yTFLw4TEJbVwAf+Ezy1Ych9QNnZMgUKmj9sgJbUeztvJLH/
OdYgYsH4oywLo5tzOzu0r2ZqOe6/+WEOsfFyIG9TBAS2MKYWwUYxsfLH+H1EDLl8OuwmTAIfRF9e
IBsJqxJIw7/RU8GzqHc1aWKnEkjpOJujzMfeKLw8RQf4kys9ugJnEPOPU/At+/tyDlgeaVhz4DvG
lS01Y+fAYXoXrkzX29VuVvRCrmMpcFgfNXPBCUmZcC7hIcYOI0NDQXRiN06XbXFKIVg2XP10bsQY
wv6WQn6Iw3HMfR+D/qOPD4R+d4D67qMa/xJhOW7tmBGOcHmuUL07fdRkfMw0V3wUP9nCCfG2iv5U
WsqoXchnxGRa/DYBRKN6BJ3sd7mnCsShjx31Dd7dFogE3XI5VGbd4eQtYIEQIuIdNYx0TrGqR1hf
1oahOpnEBt+hOXYaKXbEDpNKG76OUgPSYATNr6f+7A3HJpjeHlUmbRNZRDV+CmwmTDNauytxuTNY
D34jEeCOC0bvfXuqYt4lp6p0aU5IkSPo603d5O0i36GiGStG1NsTrQo3ln6UjpoxbrG23U6kO/K5
qPjBPXhb2kpV5Z7rb78Bk9sYl/3e8wy2xIDWqjEhdngyKrUfVyurF/+8vHvfTji7BlpsAyN0T70x
0g5+9IQkajBsKFCIxWWWQr6101cS9zx7DNpaiHTOX+owNhWiBse9tA5s6HxFG78Ki3pZUpmHqxVL
xilbrpF93WpC6IfbsMdelahTPBFUBNyKuAjp/GkTZi/vC3SnNnQL0IagSI8HLUkYhaB0LUEPOSeU
0ConSj4B/whAgo5QvZ3rF4+1/OY1MGkyEXWztGd1tiEFiUabSIxEtLAtQzjY2K+MKIajDtFppMSb
INU48ha30fTxJxkMuF6Y7BlQ2LmpHJ3qULt1+OA6xGIjyblHqNzFsNqosqdsO7WGSHsgn/Cwzi3w
D31RywaD0kXRsVQE3KYEdu+zevVm9tNf7y2B8W/0pu8e+bc8RCEl61DvgTGYYiXfv20D2B6x/fiu
0GtKISw+bHlHWzDSqW6FKi77MnwpltB9lEuU8qkz7xhyZwldoLhfeCHcCavpjk6Srrqc0oVxBk51
D5+IBQSove6a30fUNVKgbdKSQIVcLcX3dnfzanW8fAL4bfdWc0ybExrHiFHk59mXdwpvuogWliMl
QZqLVT4MkIaumwgTU1CEfcLf0VeYDtvQVJU4M3CqqdClauQ5aJ36QvchcbdDDW+h9xFe9au4ZN6N
gtxAW9UA43d5CitD7jItWX9lvBi5ZNULoHvVBSbBlxjGm+gDqYUlUod8q7+/zQEjvkhM3W2fKEbX
WJx0whtq5UZfjgEUwVQlOxyq/84v2g3AuFvSCYLEUIaHVAe0fD6PcehJvLhZ544G7Z8syntpJJvf
M0ESTP9WefCjB9GdDjcE3HotqXr8rOe7ED4Gl38zsHwOou37ejKlR5gtKynXGBi+LpDQZbCNK/N5
omqs03Qr2oKeZsNkyYcpfItPIE4HXoTdadhnjB8In9zUNT72mzWONMFj6uVG/PFn/XB5WxY8P6Ew
jDVg86Hv4rEhf+3LJ5vuUzauBkCQgVbvxcxRYOOzUDD5AzaIzkqxEF7nzkfIlPZsnpX6JzTIUB+D
ZAmGPOq9C4NtaqpN6hOKONI7ZL36FAgbNatl9hftXwNngy7tEYe0eHNIcC73f23SkgafD+SvpAgr
VYXzyjFYqk0YBpLTlvvOHBuFuw4xS7vvNHTKD1uU8IDQskIzHElIbBDOTu3stkBOAwv1uefFYr2/
reQ3yZb6jxslXCnCsZTNN6ZyIF1zbY9jIJl5D/KVxbAfvbeOzs4F2wzBLRiu1FrYGZWn7WRT2Fw2
n/ok66QDPRMRTMTi4VeLo7kTqGj51FCf2Pcc9818tDHZ7pNz9jfNyWa/Et4wIy/n6luHze761khi
0Sy/MK9zKoXKR5ZWzJl07k/cIF/5YvJ4L72+7SIvRNPtGprZEFjG0tLmnB4XQ6ypBWFZU0xPei43
3YzniHDBCS1thFv4v5/2AnNB+j3+T6U4UEBiG+ZlHVm7q5rp8ienaiwo2/yFfhSsCS51L9yN1en8
vpzaOVTwxlcT2SNmV21LqoOmfO43dPNzgPQPQMO5fRfPKAiojt8oqP/Pr7wxScIy4fmy1joVai92
YdUDdrybcezDrH668qQtARdJWDRepze4Ycj9F7cBd9kjdQz4B4JqhOvRXhbAYxjKMlMtZFBfFJMn
WTAj/KowSim1pk2VEuAz/CqoeFNmj78z54VtLKQT145h5yQgE/Nd7CevrXerjVGISinnVa2mU5ug
DkKmxN9j2zFkfZfqTRMMdlD52rdxz7AvR+A0paY9MUNC2R33qmtNAjI2xu/RkmHhxsfHpvJdBRVg
QN1PXrNaWE5zkXSMrH7VckoK2hEXhJfA3vVZgj3dWzuTfBYG2jramWigf9qs/ZGRQPLQ5QVuuMaO
R/0Yi6VcnP2FBeENY7wDt6JhoQvYIiQ0Mwy/UDXuAvcJuKi7Bttb/pKh3VyfPR/IKQn1aYFRXfIJ
quSGIVk4Pvat/vyJZ0Xy5nk/yW1jWRpeDIp2BYMbDf7gPZl1zQ31eHxRuSkhsG48XzBD7IlW3Kxx
1/VsxGxeOIy5gR457jOIKB2/FhREzJONIc8lsFl3HSPBLPO93PRHEMBcrvKz2bYVLm2ciSmGpKCK
vJy9Xk/wsvSb3d4srKh7EmCb8kMwFZDNGtOdGW7Zx5pD5N9VYfeTqfu66BYOyJS3YhNTIKsLD0Mf
rEdSfdhxC4et/F7WXveFCY8yMv6Il+hTYTNijeIKupYVo5bxKvO9NW6hdjUoXwJKAega/4l+8cSW
AsQgkaD1P07iVfvSYCvNv8HUoFk7GZrqhFSv77q926zW6ziNjgQXRNIvKuOT05z4ULs3x8ONUw90
7OOlgchCHD0LeA61T0k+rccVEJ1Q2BUhxnD7ay0QRDx69X207xSdzCP3p/T8Oh/ogJ2wEgXmIbm6
TUSoPNXIFoF80Xa+g5cN3CG9939SNCwMlZXxF0/iTnGlIB5obuBrq3zfptmARFAQiOUpBlYjDtkt
ay2Z+xNff+/PYhoJh4dP+YUBzvGsOSPBax38YbyiFys4WGlcbzqDTF+CcH97iMzMWS7dDPKWKkTJ
XNg204ZJWcp9TnXjjKbxtjBcee1i8HqVcJD7hR51G/rT1eZCmlVRpeHNZexPJPY+QMhEn4w9ZmwZ
Rxo9XhP5nCKXIW7UUIFAoog5lNS53RRDh37xnmmcqJdFYSUCtecJC5MLTTnW370FcqYqIGWjWrWQ
uy6ePSLYnXth+ULNuf8LmVvL6nQhF3qcWVTQgWU7PbcCmz2AKlAe5Y3oQkEOQCdis6+fBxJANcri
vepAMzdNHzjaEHjCIL8A+K61xp/5MZ71EXC6oDv8qDMBI8A4huHqf8JUC7Tv8r4O0opb0OG562SE
VeO+UjsTAQNxP4goahxddNGD2TM+ecOlzZ+us5XtxQU42+d9V6kDAPyETJd68eXUIAG4gYpfGTU3
ELvaiF8s2pZ39bgdJp5f4km+tiTRHpQtm+YUHcaqw/ZQiZB0webiVLFhTgomtSFcQUpanRf/n2AU
67qULHyvzUM6htJ4nkL/vSISDqhT+s5HsVzV+knCgL9Zmyp33HPYR28oD7NZQjf+HOYsELqnVZzw
QIs0qi+nk0K7Tc8f1Y1BZPK5WvE7GYcqdwfZuhtLvvPF+zuAytkIXhkA/da1ApdieadUtqp8vOmX
HE4bpor29luR91Autxk4o1ExfDLE2iBEqgUurQaK08KnobOR2TrbDl0tnwDaf1q0+aFNy4kii9N2
ELThbQ+ktzgLkCHIWXyCHwMs4iFNce+vwyK8OOWS6hqwxXtk2uYgR4iPSvwu0lAM59aXGPk6ye0S
aw9yddZI1zElKVquIGnImtPmDlqtgtAfU3EMblPtP2PZufMZK4xadNI/iJYgx0BQtNbqL7tOco2x
dpapYortim4SCJ/H7Fpy4fWT/joxoZ1+DIvYpkfo3sreL0Ez7iXrp84fpzeSMx6K9mTwk8j8ekBE
d3eolsxZ3bnV0OFF3oFbf+SFHxeVVm1Z3Rpv6/jQG21ba0j1JHIYzSPYg2R5saLcfyy+4810mOpb
3Lz+35ebT+X4nFAtIzGkbCJ6HUgWawkBiTMb/WRg8W1vtUJz3ZmXmlo6KtvSOg1Y8s/R+bGshzKS
DmskrAO7nsZwG6NBIB/2DRSMHYtSrzhEtYIxsb4QlNR8cTF0N+2OcOUctqwDynyLcbVeyaeSX/7p
M2RxqD/KbnTgbM3w0TcwlJiy/WEX5aLC0sgKgH2cJReYJR6fYE2wohq+6O+iO1ktDShUfihnSqdz
yvY0Y+jNixk5HPUpYzOP1ktOUXtdDKTqedOo4NSO6bTmT0F9tUpXZRli+1nFHudWPm4H6OdHN7eu
ZD8yHXdDfl9K0uXf+ka01uA+0DrJyuIZ1xaPrfmWmkdQJ0mBGyMDXdNBCbeQuak1C2FhcEEd37lr
gL4aTEbP0HuQjQrMF38mOlB8EqKBaTQHhrzPu1vQC08bkZiU+Qj6kaE0Q96J6nByu5u1sBhkyZ5q
x1PXR7IMQuLNaWiIdIl6KhIZSoqvB9cP2R5Nls5AmmbT1gv0YogBpB/j/XqR6+u/xkw0GjH2vbKU
EmfmKncgMQk9cLKKPRohM0EvGLNAB4bgjf71UK3cZCImFMnZRiQU466xyKPSG3yEBhDHORouh40z
igB9M1euBU5aMXPmwCSZ99Mx8PkHRLV3F79d1BljHbib2T9zPxfCxljBL70wczNlMjEt9dqxQ7lw
1jPHNX2Hn62nGhc7foF3XSU3GXcBKdCQW1/qYlkJjbmbGV/RXRYRYDltOKHiyhJJUZFTKmPPxxIN
chfERZ+XZ6ftEqNGcNsF7sLiAndQRRBT2lDbkxCv9YMddeRIJQJr6h2OEp3zm94hYo+I/1KLTZr0
GLnzFZACWZ+BoGq6cjjfAiAGUdqLFrzD41AjTqtswibFFGgvBuwgAY+yL0voEmD3FxliPJTAyokk
yiM7jl3H8IME2D1ohf5a43gQM7JMJLRNT5pFZjh92zcIQIKsCWHlUBVdSVKFE0/pu9qN8Lsc2SLx
vV+K7pmjALtQ6Eu8HUBR8Yr9S9xqo6CvD6YRchQy5oeTFn8HxoLrKHTQtMsVtB8dl74FMVu1hYKl
MsmAVyKVAq/CMSL0r6lAxD3ihzSYdmoYqZ+b8n1/v3TGXmA2lvY2wZUQ1DtcGHs5J1NOpls82SZZ
Qrk5j1mikqlnPxz/Re1Ska/TZ+2gJFam0oqqm1qzU4Xo6EhzzMh5eoYtYNFtoetQv2ktu57p2o8t
fVtwrKMCS00Zi5QIQEhLKjIWgqJuND/0olbWaSYq6JtaEuZ2zrzS5cW3F8KwGJ7jDHQktuFGAhC+
KAeMBskBszu6ETVgqlLLpljjK+XGZdNlsF2r4rKRg7HJ/jR2qQ1FRP9Sj/xJwu+sDwHbsCSGcdQT
jbkVSf73YMs3RErC/x3cp0y3Dw1pQM1SVfmXj8wwsPnod5fmRqyE4Bmyoq1kjCSEvkolrFM8dr6U
DxVIv8UCqzclvzh625OTyZGIsSs/j0z23uV2ZH/Krv2viUnUf31BJKM7fYSu7LbRGFq647hr5d5M
vNHXctNXEJX7RnzQO2yYj3dtRao+u4ZJzQLvcUCgimfZf15Y0ylyhZ00hhnHNafAi4cu25RfUWJP
TOpiBCxIkX7ZdXoATlSzCGjqcdqQgMuONI4Q4HmmWCP1XelJEoY265chw2iwRohSGt5QKOX+9iFf
N7GNpWP1LCIIOcLZ13++HCdXh7QZ/Ujc/CgY5+hDyygyZ4vkwSW7Se3GBW0LdqyYM6pRkIYmciE0
8L+SmSyqnHc1Mb9t04RxjpiLX8EqWEcY6H4NH/CY9QYc/X80QF6ZnO4ehC/bwXitF/dGeL6z3AXe
Li458aQPlTIEjLdAtHMREpu3Jj1e5Xvzfe+wDNPFSxxjqdkm6ZtF9jjGqPoHJw7pMvK7aaNNhNGy
Qpi6EZF71C2axCOCr64FIOJKFXXOTdFQd0vwLLYiQQQ5YgVLvNNbbKWJnq8fczdPwEUXC5+nIRGJ
XnXgDsv1LE2trjZ47Br0PufKrc+lIOwZnVzHsLQnNlsd1k0YF2APCRZBcKWiGqKFLPKM0qfNeXmC
lS+aJTA8fjNrEGDUNY8YnGEEtuPiqKZgF2d3NuC4Y5cY6wi/39qTU+KwzPCoctLJFC2YV8pYK6xR
yYoaViaLJuu/qR5CTBiGJjF9GmpN0lVCgba9rIsS7aJ0Ck1Dgmi7mYRcduNgJ9czSj0aNiR3CtNs
X4VtN2jeH0HtA5QDw3shvClr85H/Q074PQbHuHCZ1xTRM540GtEQZOcwIziIPhQN7edzl7orNBi9
x8IwVcR2Q1al5mdFt+a5tha+cbogSYy3dwMfQRM5PIbCoWSiyy33pv489DrRgtbYM2VdTb1sHR5m
eXjRA0wopa87BGNzEp1XmLndyId+zLmDVGIco8ajghT1tb5nl7Ag4YLrCznUTtZsNoWRkxgnonuF
J6II+qZUPPXzEaGgVuF6JGYdvY8Rz3BLUF42HVYTklcgh/tq/u2Fl6gt2PZv0oPu9CiSri3Aj5V4
0xxFaYaLbd1hm2d2XyHGr3fg31HIlV+CRZonefWCWhFKBMiz5xXsnVh5tn7/E1H5mz+czi3rqDUj
CMoZ5m2UYsmzEnJaR8vuLPpC6bUV1NrLD0JZOm/4NzQsg5+om2gCfxTlq3nmc8IkmNCLdI96UeZ4
22QVMCIHrpLvDOQtAXnNs71NAcnuqB2YttopkOBDYjBjQXmdXJUyXfoNWC3fI7KbFFsxMoYh6DEf
UX+BrcNFP4mfZe3okKT8JabO7bNazwCybPGp35P4EN2rNmQ3lUgm8lLTjSI3839hv3dP3cOJWzVP
FdZfJZQf59A0bLoe+RpNDPHDHNYOt0XpYNcwcMofLhKOclbREsBKzhmTWSAL6fFh4d1OtWRYEmFZ
MWHZPEid7onWW4DpMITbnUlucrQCe8vyVMB7vTJBFe5ceIaqwihOFVh98y2INMkHfSE7wGpvC7Ga
UMtPzrExWkznIviPY3icWZUUq8cycbGN6KGTYX/kVjOgebZuBnJnpjrWLU6EyU/iUCIotQQGJtCw
JGL8cvRp0CQKmYlayECtVU84o0Q5fZ1c92gBGtZNzY6dlgdXYOUQTHZsBegI/YoNO/uwNmIGeD3d
ZnQEsH1iDYZSa+3FlsT5H5vYnwSQWGu81GaleQCOJ94mJiGYJ3ZGjFrCtD8H3XYkbM6iHJrHSBc1
68z0qvYorkbnZRqkdIpvVHiHJjzIjIExVUxcaZyQ58GaN09NTB5V3KdQ8O8KIrQopV5tLK8zoWJ6
ayFrKmJlS2zmBFv5OObtxJ34QyTOEM35h8yNI4OCRg7af9DmP2xrsN2fKekpQYHv9dNtLSdtdMtT
SL0j1YxEyOnRHnq9woV82UBql9s3601C3peBETn2oclXa5bpKaBA8nPhSaRf5XSpQxzANvbscDwp
bVheRTpwOduBVMittgp0fMXycVm3KUYonGqxJKytw28zJsO7VYBpGrUtEqMpOpjiVgQ6JKfXYWN3
+m10lCXUGXfyuYxXtvZ39T7sh+qPldTsmMWgChScP6pwEkP4LuRe1UrlweBA++bZt116/yCATc4F
pCJraas8AD5EWQsFfahSDWAUu39eRTPLJnSc7kRVehwU1t+ISflYDw8GIGFO7VKlxyLDYzosNU0v
oEzVb/F+SkQzrrONyfZPmbDMUbGvrHd1ZPTMHDPOHeT/ekbQ3Q160benmWlLX3XsXkuPJsAjv74f
8hrXnZl/SQnuMQEdDVcfs0/7E5ipwCzf289WjXycPiq3S9hqWPBbnNmPrEckVHYCQS56x4Gij1nq
UT8oKFN58UIPyfzKmVGUXugADhrF1s6gbX1k8kSM8/dEYSp5gOjH81uYOm8Oj4lJl2KG7slXzZVz
ugrh5Xkp6qffHIoEYIrgqIHDyjz4MjlyoZbNv8T32EbNaOqneLKzkkwDOLxgDdWGlooh0qv0Tj9g
09+WB2lxE65lamuEB8a5dtS3apt7AIl1rc74ekGWqrew5SkXA5hEf/CMzkWjoqXuukXpje10HkDb
bA+fLv6gFRt0ExHQkIeGsS63QKpMex21EItCEAowU/QhQEAutg7X4enZzk9tn/2liNn7zmFJY9NN
8tzJ4vz/+ZvKuhbu9aH+atsfHFZT4h1qj5pj83+/j6Y8xNjhjcPfxAJ2yXhptpYvBe9xze1IfpUo
ReCT16FStSixm0JpIHbwPEJqVr7FtJsDiqS+2DRqPZn89Tsy60e8rLGr40NoT9BVgJJhGZwyLbHJ
wUoJf0oJOZ5I+EqQ74y3628Vkw+/X8SkfMNBLCibezvasBsP9kSxXO/NQ99H5EnXF6qFE5z2OR9Z
4DRYHzA6FUm64qjQl7Uuao21+e+7kiwgRAJaJxZylvkJ0OZ/rpdac5dQXdrUNw8xFl4DDJUS7Fr4
sb0FKzdqizBENcnoQlFma67CJ3kdjTQttENnC9bw2Lr1jV5Hm1Wa58REDWxj2x5iyECOLMHKjuw7
3/jyBBOTsmsZZY/QLHJiZpubwitHklllfITUqlXP2e9Lmezdbs5ip4OX7DP39raHp5tfK+kyhkVX
rvyd9BB2jiUkCEKcQ2xOnqNkzJ4oZbt4tT8zIQXfm0sFCIUATVzomw3vpt5gSxzmzjBCF2rtKdwG
5hKIgPmd67ATws7MT5jmjOCZRd1j42aFtNUI9+kTlNziQdYMeWfhFF8UMIOy1ktDL5A1wj+M3mOV
mNxm4Diisdkjy31WMkTzD8r6gcocyaERAVDDaANwUnt2NmlLqQqLryCsOX9g2Raz/7G2VtCCH4st
Vbq6SG89GqsX38c1mG2xNAYYPTVgTX27u1Emq9ynY4MNTqPaQ4ZMIMtpkLrGh6VD43PnVzkVshtA
YFTe9vWXdBXajDcFyrG6ReYoFKeQd5dFT7YI0FMe1yK02c6+x6p+G3M2jDWF6nlYZaioS1sceHfB
R1dqYbxfG5A5wxJU6lcde6cVoV1cvtwb1U6OZcEVrSK/ULihFUngLNQo9zo4bbfMuRcDlSyi7gWI
fgDvoraw+x+vGVOOeEIVpIGAQtbXVw+93z3GL0G5TKvdq6yLTs7/njNJ/KfOojCGpJCoTICN1y6w
KYGHgZ8rNVFvt9UJ1G0RWWpCaB+CoQNo6cpSPEVNG+duxfRa7A7SgKBqJKnVdg0Y/enPS2meGVKm
NY1ee3MioYw22MiT2Y+XLr9X8tSn1uKevvHn4OTsFyxMCj4ETBl/dLePaJCFZjG2GZmuixg2qiRu
kOrzj2LGUEM7fQxhRQHJy9GmmbcCCXRRCS4sX9n3MjTAmzYBC8+ASebXKAXKL4vZkWZiWysB15oF
oQvuHqgdVXGVboYKTkVav7jnNJKqGuDVUQNSU/LyuEPlJfje57C6WtiLRB2L+nSmUVaqZ9/+mC9R
BenQtXulvVIBrXbw7cJzhRWqyoWZkujPkvHkEBg+skvVoMRP1ZmbXwKuqONIjTkQFt93eGzOvKgD
ukpIBmMdLXA5LOchZO2P5tsbk/2w8Wv43cyRY9v8tH3KEDArBicOlwymPz+dt9PEFek0EBJxOjm7
H+Hd6/uBekYSXYZ8J1IPymZe0S2DbzjFs56BrAdY5CYPzJK4V3gaZE0X4g4vD2mG949OGSL3YLfu
III3jkjyYEAfyuYsHFBucPDgXIsc5RVxGah0Fl1eR9vQyqWhtPHsgXIs+w7jBl81Mzb/rwCBhfsP
vI10F/xWzTZBMq+KhSjMtdUYCG2ihWdrYLkvhpKpbShhNjqQpCt3e1VcaqG7I79NGHTKQucRze8b
F924fpXK+E3BU9K7z3/2VnDorMoQO+EhL+3XqvpqFqhuInqgKWz24EgUYBIu/29NhLX1alO9420b
NYCqIq8yd3TblSQgEPX/n33KplE/tbATtiLa2W0bDo5BsXuCh5kgaKoD2vm361telPNZyvW+1K3H
MaTaHTvDnf4FydkCn53/IJWZgb254w7wfOYeV9QyT21JlyFCCnHwf+l74fxxFoqTQMsQ6X8FGtPn
CH258IQUNZ8f7DeETebJA+cb+h/zN1wCh9vfJy1qR1kCTxFFsBtx9FJgOwE7g4t7W6oXMXSlkrqF
E6Yg52V2+FUwlpsNRjerwnplPdP/C0qZJK8HhNxRVh0GyY4BjftcsjZAocxIzNEpdzG4mMwc0Xci
GNEyESTE/AAci9J+9fc/pV7+bHAj2BSi9Lopo23m0b/WGZBz5zP1frrTEh31F+lIUN2iKiwAZD7d
UNYdyxdNVBa25hkFZ22aXdXZ8PQ3Akp9gof+bKrELqptlaAFGEmDOfy3BqxSGtd75BT30HqQgJO9
1mJa6kfqOW/UlK+mrupxXm/BrOTArPTk+/ZpuPFJ+SlAFFoSUEM596vqIJuyMmo481759nFVCHhP
zYhNzPhWtLGpMrlG7utzXjj5gyvysKxYOt78Ekvql/b9f7rcKcCjONr8XeBcZJ5eC9d35A71f16J
J7SVj34LfVb6I+LsXrubVDtMRLG6wu03dvZ1RLyxpLi9HGeJgtN5RSIvsPy2pi4/eGIsmQ91AHw+
dpInRO/4Qr8IrY42n82DNYHTPFa4KjAuUZrXHO5RbQJHGKnZmLvPDekPr1AFhvleay4ZNsQpiY3G
zwdblMY9BqXimOPKbgT0da6XyNGxswo7zC6YKQGv1vNs27A8DzwWKEBtO7KaOkeHlUp7FOy8VkiY
43kgdsNUB7E2ooOHipP8MM/K9tTt5+Gzr2UPw809tzSsGvM8qpfSNaTc+fvP1Q6+bpyzEtGeZYdS
KuLcHCpQNt7U3bC8q9se5DUBxiUVA0KJPvmqPo5t8iKf7Rz0oSCrrBEk8Ol/qXGJYCYl4JHQBDT0
8pFVt7uUfQKh6+gGjfeHbEkGZxAZnrBrDFoTS9vI+dK6WsVAJfosS5qfz6UeuCl2Z+jF/EyXjduD
ylEiuHoT+gAc4VP5Cx6xNXPcA2YmQMwH84UAh8nViojl2GO9XgEoArhqWTto/eraGfNDJpM75FvH
7BEFQwazeC4BYSed9QtLX6j5iEpK3vSC2tVAILR/P63XxfSeeu/D2z3HLoERX8tGTFtr+fsgUwKo
uy11J0f3MQkwb3GG5jhDnz3amMBhaeBRIBaOazZmGbvwwqL+DW6oOvaOhOJbyqfsW8IWhoDJCSG7
eU/2KJZxotZe/gEw/1I2qUcmPin4q9ay9+Ja9IZA356NRYqSFHpsJRditOQ61tFzYBKF/CLAYDbI
OiRzlpQ2WQ0hBbMFY9a8w2CkrxocryIe7e7cdQgd0crx9d6+g8DJXPIUDPpe87xoxLw0Y5yLv5ia
5a+PML96SLTQ2REmxvVEjzAOk82Gkd5uwlN6DAwG2bvuOWkqrp4WWx7deKILLKmHc1VXxRaVOCu4
rViGBhIydzK3ZbySB6o3cQfya87XzRWkoGglUgy7ujWKHG8xnJ3dnwDktaA5mVfyiEKrfnM4+KV6
eYT/DoIudS6xOXL0SF1nCJ2EgPWoqIZZwJr2U8KSqbRYrPtSXycNNPXLJwwsF9rU8MWsu+fT/z/4
+HZk65bu2U4xN5pf0lPjbJvICoMAT1f40v7kAjSIs9ZVjrY15qJs4yrqoNyZoNoiAtipqo62WsF8
tKEMQRiH8aJRpTqqf7368WVKs4Gyi6gT9t8DJNzUYkaB4josNGd1upMeIOM0XNAMaZdzeJ3awLyP
tCwg1BRas6E+wVEBXFeoXIm9KCFH3om/QaBBhyFMBDw3MCT/bGGNM51Rz+m6uzVne0Uy2WrCVggu
RDt1RWvGEi84OiyywkFk5A2B9KfFEAGUEegSLuydNoLv0imDjATFy0cH/fLxSa6GdXDC9R7Wg/4B
HrUrICKzqQWhpVdJ6V5VPTgPmkgGnevMkvgSk8YY8d3vh/q5KPkNVWQNkzOy5S2dGBqnm4KkbE59
6o7ruvKz+ZfgSDNQd0dGXcsen6Mm6pQU20o/r7Bo8SQ070TmImi3mzz14bJPb0D826cAybvoFsql
ABncXUCQi7kPpI5kQ5dkOKl61XVvT1qMUgEBLqq8LSQs5knu9SH+2KfH2JNs24BSkvs+o23lPwIc
JLtdcUXBUzwyueMqk9EXUAkJrqsafGVhKanq8n8NdVPGoxD1PbnGHO5a3HqEiuVtqo+uz2m7I6fN
Y/U/gY27xfzyW7D3nFAuaJ1MmURqkw/KamjUDWVl9RlgjJEvx89fCcH11zPNGrk9sCMUbvT36w0d
cWnG1S2hKhReBx6YCa1ZeKP2pszhoZY6RCkSfmPJqYIP/OaRIhT0BCLkLIuQeBikgpPtwU1ldY4h
RjiLgswIkGYCEGIUEgZ7KGHuWs6M8QCIG/jviUhiyrftaBOJXFv/8rHEsIWBAgDf/RaL/GW7v3pJ
PiOUVjnwKJl/21dYa7XACbEZ5fonBaT3j6gXzq1GDJ9cYk5X17RobNTBsEacw/bUlXRMOv0ZV3K4
zMndT4BSC7gO2ci9kmKK0nOotvnT64L0gEAn3Tn8UTsUoHv20R//9aBe2BeRf5CdDtdRJmB77MC8
g0OuNlRgsl8h0Y6Y74GxekisPbzScPb72vcO+/o8q8ESM125nTWbaSwPwrjEfdKGP3oQl+6yqCQU
nyJ+AQpN2Tistig/nv8q+TKt41PW+k+YkuDiLfR0o+7KyC9n7bt8HUUelQ6W6aYjNF1pnIGYgX1E
I6bPMvIhpuRilYS3KNkadjKdmAs5Y1xsKVYExUaiobgytVNhWysrspHybKXMLTHQ1/wq8QOiBHXU
VKVEEg0IoNDbhRQRJ1bjoFTBddoTpysgLIR5pXRj9Yr0lP/Y+Lg3QTAarmUdVjxasJF3pDl3k/LR
MdIPOKjO9ZaQrVL/1qRpUBRBgMnlBtgsh03K/5PaURjfm0RkgawPEx1kTkxmwyiyqJ8iC/3zbBme
gJbfSnX6ocLy0ZF78oezZsf4c9Z0ZRCNYvqxND0dwOO2oQ+J3l0awl+CX9VOlewEf43UYJvkAg2R
NRifj/Eifu7H7q94NpiNe0BrMU9ZyeDyvQ+kBeUAhZcwiHQPvKn1ciLd/oiguTOmJ4y/X0v8onRc
N1OGzdUfASa9Flxld6Wwr4TFEZ7dp7tvoxJ0MqYQdJkSFOCZOkbni+zOORk0JoZEQulfSATavfa4
bBYRG2HnElwec5VC4/NxxxMO320yV5fDmyNLTU/vlv0t+1LuaXna+tU1mq0HNuq3AdDjNNIiz3lc
fsMtpNjtaR/kIkS+kggG5fYobFcQW8CVxTSidoXZo3PAAIWIGiw8SmxB6eT/mQbI23fS+ikDwO/8
SulInEVgOix/toOCD4N+iK7vjbQoQj/+Dje+RIJwMDQ49+6vWpXI2mg+9Pc7e3cS4rtwYCL38CO1
7naUfWbFwRlFrwARmB6XSNGa89LzqDxeQ+UjF9aMsVS17+Scz5Mc/vL/b/ZLR6LIWZ2thUds4/rM
Cd0Z3AIPwc4hyz6iIiCc+uDepDtM7WcejjAMAEZbnl8ujbD7JzeSf9oIXr3m7yxuuxJdiad4+2ma
ClcgtpcPaL6wgT5Xzx4VE2P+SvVDmeeqdVW0avfnTlL4E3trmx84KPpPjiV5ZFgWclqFzksiwSNJ
zkMyYjOGZWLk2q/aqYF3eR17d/NsBDYFw8U9hdbhppshZf++LYr847OlRtMOOrujhnulG1sdFjjI
sPZ9dxhwCDPkkD+Ms5vkaTera8r7Z39/pNRpr2wkBeVxu7yaZ5/0t/iA1aaCmNbFPSCIPyetI/4/
GQztwOmBE62sUGOD2jQq552LMNjoJija52kCsXEZihhN4ksqxx9eDQmK9zH9sCIjYqSih7/slaRJ
riRYUIDo/YnBdGA/fCSzoPYMk09f0YGUUoVlJO9OSsGMoolozOCvm5dkgOO6kLELbg7nBGMDnjKe
GTSd82Kj0BxyMFXN4d8r1PLQSLL4avW0LUeqEqlB5sQVmr4MQSL9A8cBagMXfZ4YZ5dxIB+86oZq
z3P23y8+EQ0b3cMa/24ruENiK/lq1WqyKa96JFkmbHsypj+RjkNn4ioR+LB5tQf5h08ehfkjzyog
GFKio53elA9vob0YtQs3k2ekBhgGI3bXS8rTAZ+Oio1QjkwqIuXMa3dVIeypPBOL2i7YbX7QLpGC
NI1BAcH/Ezwviy2LT4ifaflYX8dOpcyMoZhz0AYK3su3kOWWy9kdTpZi9eK9nkrKtSe1tDN9aEyV
UYeE7Zx8uurG+gu+GxlQln6IyjinzjW1NIdhQbAMJsNXAlXj6VwS4V05i/piBPwf+4l9J/PiTG73
1MTbFEHXbozNx6t52v5T4zSi+7mp3aMXSfozM6USRz4Cgx9j+0OpFTFelCY1sJchD0Dw5KKuBt5j
MxU7AYI+mNafDNm+N023Y82v87GNMSK0fTFa3/euII/1v56QO+TMrJj2n6U9ITXFCV4qysTA6I3p
9WIDh63R6eeWJUEDd+xHWuZECHehrMJe8DLCnkbaDearF/berOB89Kj2V3wA/Em6hS22mMb0viiX
uh7cuez0uAAvbkBGozNo4plljKfxHojHjkMtVYCW3GNOgH2K69F0NaYAbIaLrN9MsvhFboBmOUSR
7E0Ep3tdfACbRz4iREPuwl6cRERgIC4buRhFzqHWVeDfMVLmaWgwkoOx2INoN0HaXQMrKjpYh6KY
sMI10woCXlgO113HCL6K52MlT+y8qmLwHoGdd7ktGsk9fycxBYrMTZyhC6kX0e42EJd/ENf6b7Wg
1WSmT7tbwPr7FxTTzhQP17C1mKXCGmveRcUAvJNx8rN/rSiXx+oyje2mpEDwF1R4aeQCYq0wizql
LfkY+tUsMsueTBueG5xmFw2TubEvt8QcePCqZoubrlcTcwFKLQ6sHGpUpFKTheoyuqLEXzHST1Rb
97w0Cej3iafdze3yuf+h2ugXBVcpF8wrOIzacap3YGGzckzeHS47p3QWWHk7McRAxLeDs4emt+dS
btP00KsXMvEdC93cVbjhnF2qH8mbUrWwHTh1dRtyMfaV2uggksQR5nd0Vut+UrlfA5wXuRS/pe8s
GwLU6dVq2DNyW8tv7dSIwOlwL4EIyA7eiBBiHWW9EB0yUxMEw8/AOE8xQIzfuuEf2rgOYjG9WcGX
SNISdFF9MoQMRJn5/cj1nh5M/bnIGnBGJQjYCg+Pyq4pe8tbvErWNeyi2Pv1EvVTawZ+7npBnKbh
D2/SB+NEbiC37ZGxbPvXo7bi6sXOkP4XxuivqKxON6jgBV7M+Il0By8p+mLpbYlDf0rduKBYKrbX
vIxFUbA6RYxCIT9ldtE+/8ng9A+E1cDe6WIvONAmF0yEs3/iuYPX3RpqRWGNHwO9AunrACZwgwtA
47FpxQBcsCLlbWvUnQkl1wq9oumF9ScFzLz5OjGBD3SZRPfJVDGj8EJ0Q9hP4Q3/MNbxatQGL7vh
6Kw2UvxXfM1GHDa7dTbI0WQ2jTI9RUXIOMzT7Y4haFyY2rjtJqhoKC00EDj9wQ3bii1DJ5XYU5Zj
qrJiR4rFszut5cJlh1Uf8fVVFRyqUTNmzLlrRsN2BK97BD3GLa0oIIYhjQXey+p9jw04pZN2VUnw
SDBQfivhSxKIX1mP0q/ELSkkP7XjHcPGyR6Vyc30MuNmNLGZkKHVkQZoNgKPbcgp0O5aILgSwDJE
f7ZMgKJODUtBVBOLmzQhVRgZCImypzVzck/GqzIClRfDDNp3KeYA24rBiiQH25l6ZfTZAoNzSJMl
QaD3ev5e3ILLqXWZlM2LlZnLwYRxndgYGBKQ7Jr2yE1eoSu7wfaqky1ast0zWzgGVhBBydSrgms3
qRr0WQOFzwUKKGqj+y2iWEfCwY+4EtOeS6KtWmsYmK0DjRw+dLpqAPU8LFvOtBuCK0haMCzr0tX/
B/IwkeXZGbdlXuzvU489JiI/9+Ex6KqdjhZuyVMuBlbkUNMS3xe4W9yluHwWF/JAIXMNP/nVd2C7
0oRj/OBzWcXEdFY4Hun4+7qj31Bv74cE7d8DFgmNo4gt28CH1ujVMUtfxUfJUaB8hBo8Zk3AIHbT
hGhuiwLygMPY78oc5qUne6W0JtyPFhxR1tdAxkAEhhp+a+anLLN2sGFASaQqE66M9Tx9dQFd8ptf
drIzppIci17qeA6+nuNjJp1cXcLmPzcFI6wbE1hUwFIs7EcTYJck1r8qU+nzzVa3cWeWn5faBvr0
p6Ws61oQCQ1hGdfJCpCsCTqyD9AOXCtcOUSYyRUoX3mkixZ8ByPndm+whSjsppyhvYBMGSzkphSR
3kqHMYa7ay7gfQhME8Ynsk98os71Ivsjb9UWdNpkdSbOKmn9MntUGGNlrzjBriRdkt+g86C+zmcA
+P93iRgUU36oZravlSpEtDOMts2Ol3x1l2gu3Xn59Lmn/5iVx8+95DnyM40h/LHkNup++0IbRNAx
uIgyCcZxNxhqEPFDioZDePbf1gL6oQOMBroKhx4PTu4tr1MuTM/y+QVJkjqFTwYZCHTpjUqpUEs4
bKzwxld5+OsOK4kbkcg4eyzBhpzmfz4YlGsMrLYIRBlLl8Lgy2i/r5HjoXBzIssxPcnSht8wNlhe
qZylr3P3OmCACtFJm6Pb/vGz83J1vSUV/pwcUbOLvrz84P+ddn0dKqplSa+mAyHivcKS/MUlcN0A
sYOHQ3N089DCd3FSXZzaz/7BR+Z97+DZvTXk7AEp/RZgY8IUfi9GpCI/QdgI/XWvGf5p1N0KxrQM
odUVH8JgL2MK+c0o70ShW7Kq4IebJCLSrh4GbGGwusVwM9vwPkRTWeQejs/UqayEPf/wstRaiq9j
SG86bwkKmx1DkQ7aOk7Z+i56cj1ZEQGdaIdNuQuo7VMd7DA8JgabyCjyBtZtHe/MJGSoyfhvnCXI
H9EFLE+9KgJQgE3Lp2ypqwgSxi3n8BembYutg5PYAHL7TdWjyYPNYW5FDRlUFR43u8SOKjIzZc6M
XkizfUfQHr/dQBTwkeBT5le+LnS1DRKMwAZo8D+z8hZkqpkNIbrvoAYITdVrl18qgwBMTEjwaa1/
mv4snyfrYX5T1++ruHBnogNld67+zwfIV7xwG3iJN79XqwvPIVbCLSLCdpJfF/DgZ6ME9pSzEKeD
UD3Uoz0Z47vC3goSvLydy42lzT3iiUxlSpueWBxqdLT8dOPi+W7rgyE2MSozd7qgTHw99tr7NOBk
BbMOcnjmsvexPuEeOzRcvWcvBx5ZQWPbPlRObs7M9ju5Lu5b/Y8KErqFrko+NLcaPnCgRgTuzjp6
6zBb9OTPu8973QnGDiPTgrpErESKxWLrlBoo118ujQ3Y5NMzqaP1MtwTce5FkANEoYnRY9KpOsgx
6/WjKGbfk9vL8ZCAa3iFnkog3xeM2QilJF4b/g0o9jrhVP2a24opJjqsMKGo3Hkc2TNdtR0ZzlIE
jDSoOA2CmB06aeZI5QZDZrZ93mdnfBIsuhqR8CQBfVUJZSYbsrjAiH3dV/lvm5YsWcLMc8+MUX8R
gXIwraJKwz0gSkVMieTVSz/KlwrB3CEG/hATWeZZDVGruANdVvgg5dIvLL5g1E1JB4fHv0zcVBpi
L8/8hn89+eYAvgCIWx368koDUSLhs9aRigGzjR621pZgKW09xMU5IATvGntdl4Gc6h0v6KDQQLe6
RkR/f9izSYaZWXNpoX9ZC1+CmwbFwS/r5rpEar0nlPQIBBwXOMZhU6crQ3fVJ5+kxon3FnFkNXwB
hxy2s+DHwsbhEWpxWlZ5+RHqMZc9Ejfpy8KGkFJwBDFKi6otrADbz3H6queiBwmMTiI8QxqYJ1SE
uBYh3Zbq6l+pRY7ddr7vGlcbffPngUW9YlK2Ubjy5xM2g0m57FyFF9b/e9j/E0eShhn9UqlPixUu
2YHGkkOpXLCy/a4xvuo6qCpWZPQhDfbPP1gDQk4qtBpADYzHxxMhrUhlQamTUrhCX540v3XIgA84
gRthXwwmSDr9u5CPwnQs5uAqTynNKk0Ocu7wAv0Ca44zyzrhceTEmfvFk7cq+pjSvsAPFTiRR2a3
n6TYCw0sY0n8CJTl1tOXRQdy15vp70Rk4DVl9qWl648IDFIuEbsQSWUTtW5+SKlGFU22oR/Ny7jd
Kw4k2HUM/buRgggFkzOkUaD8akAV5vPPhv7Yfn4zLD45huFqfYI/xhzsOvuDyJcj7fZVEa95ZnFT
WQdDY3Okkpgtm1q17MeiMh26roSiSyQsWfFswBsuM2UOhGTDd2H1JQj+Upv4F6Nruvcmz1n36Ihx
roWbNilPZSF73B4mVCJLbZmlxHmjkkjuFIQtDKhqhe9/2Z/2Hi7719xU0IC+Jo7aGjJuxMLfxSx2
F7QzxPgZuvFE04O9s7lgksAe/ooonFdsjPTqd6sLrNSC8m/9IOc+GR7p2dMJXF/gbmWhZwt5n6P2
M3q+Ooz9AgConcZ0bnpBGT0CBD6H7mPCjJsQ4QKDJ7DQNkSGliuz7bdY8BT4B5jQmY8lzeqSANX1
4rbJ5q1qUr7rJr6+fhkokZlrx/B8rIgw+iw7jfqqtst8wiCRq/verP+V54YGe9tEvMFrH2CBEa9j
VR+os1WqcD6OgcdGDF3jkG+Ktcb/H8hPlXa8GD0BJ79tFf1QDeGAlp+9Af3zeusZNQkFcw/6R/ck
uiMrwDvocW/wWFlXvBloI5PAzQYeL9TGm7R+9lTMD3e5KpXa5Zlof0vtRvD8i42gVY401MUTB5bo
OclUwhwkBwztLRNCz9cbGtQwKMfq5mO7BrsHmza4v++CQk61nUpUMuQeNaLZi4YiB5JDSTeQbCZj
Z97u5X6M/1bNZxGh5c72iyTK3mt4pOe1CX+dlV+ctWVYt9WrMKlH2od2hRT/ikYQ0KST0CHopfX3
tJH3XqyL0mWaqHio2RhFT1vQhN2MskChkXiC021pPYVXSj+HAWQf1d57Lu56oWffr2yemVefe0vt
pT1CA2JEssIG/s0dlCgQc91e76Zv+IjdE9mpvVM0IKF8l1TK089khNnCMjvoxNARJeq20qM6C4WW
zyRaq+0KJi/WNDWehLbzkHe4lsRFSe5x0Z3bd4/ualsnIk6jvlTGjxT3JrFMDQUjIUuydSqwTO5m
IhPfVM5If8d125jSMTvflzP9vrwjNHYrurwZiMwlEibXljmTFn6/QCVuokcDQ8vN0tDGuWrGAGNL
Mt0SOLeAPDK9MACYhRAE3FeH7ioYL1LlkHs7RinsRgrrGQWgzExhm27HajtdoByCtP5VGT4EgIK8
gQ8fJzx7nKcqG77O06Sb23905fIHs2J1t0A8+k6KW/VMYFqWDaWipmVxpCQqdw+TljQbi/RaFBeA
Ta/g5YrPWsdF6AagvYF2oVtdXzLF7YQ3Z7Zd1JjUnvGgcScilqfFnIeIwlkn3oHs61xKBhp+x+31
22Y2AxpJZUHTWEByY0uBAIQ2LZICwPMpdibEUAgRqyWlAURLuyuF5TtC2cEOOCMySbgc5GBYyvbA
8WyMtg1g/SnybqyBvvhl0mzXOxNaJeG7bgpq3Exe8MX57xtjjSpXiMi/egUegYtV48lqNXKDdNVg
vch9rkk/WFKVzSTrvHpckq3mL/zCad3UKnY7c8qRQTAjvwTfR/7cYZRwn5i4300qLjtubNYRKwAd
5VSI2HXJMEyKde0u6a/M+stmjfAj8179W+OzYJMQU0/4ca+j2HCLTb3+rVvYRDSZva08G9SpGt/v
GAOfw1LeBzvZghdD3uLSI1O07R/NUuK2n2Oen/7PaNfkmu1EqUN1zEMkzBP9OhXpL0AUxETI5Zpy
9D30RdjZ37PeLv1cwv7o5Zl0211n3ewmO0EQlL5wWr61y0pRTdDV8jFORh4YIfIqnXCdGGKrCJqI
vk42roSAV28CagsMRgjaTEW79FcGImEJ0eW8TSvyrGY17o2iBoAjwvPbnmIt+hOWF5be8hA++VOf
gXlYwZYR1CVPseM7ykODtqLkf3T+VDuUYtAgD9vBlptkKehwEobYut+MWXjiHs0oznTuDdHnKkeE
qZMrVGig9lVB6qdVm6IG0WpvmCM8gu3IV2UZ6ZIwrPJpe9yaxWNfKDYbMY7Gj5jRhqd3ahQ/5udg
b11DUgN2W5kOCvqVxz8G9BhbFyEY3HZ26XI1PG2921VqNRUTPA/OuBPGxfQv4NLPlZ4FZPodGZQo
JZ3lsIbQfokyDBoF+s1XqeE9CjQUnkxOJZ82PV+wLL6ZLYnkW0/HiJaNjVdvMTmGx9boLcb+GvTR
D4CIKY73qYAP94n9lwTqqZlgjTl7vltgyYM2481Vvp9VnUTNb85hqIThw2NOb0wCM8wbnzgM5F17
kDuDQ3VQY9rCQlLb5NWEuqUfHq+OZgh/v49UG5QoP68xszLPiVjcQzIV40M6ak1yEhsHA0M2Ylrq
CD+xVCg2rfiE/idLIANIKDp+bLHgJ/NQIuCeP9LGxGG8Z8IL9TnfhH2raB8WXnAhiI43xzkgJHSh
+87QEhLS/IJzna0thF5VUFN+ici5c2ukLccs7/EjI1IVG7nayGcFfckoGsny8JV87WFvL7qSrGJB
w2egm/La0tlCHUA0L8pJcG40nx0I8ouBA9U2F6Kea7IecFGbSwHTWbkRlwXDUGtMsJ3CcPM7ZUwr
SCeNEoCgcv4jV5HplotHVUnszKtYBojPsvRPd3lU6ziy3NNywUR1mKFmNLDupDstFrwsbrOZP4BD
+M2VG7KVXupx8c7Z+EGaRG9DosFkX79tSaLCz1m+2G8P9eKPdWRXZ4zgU/vuL5HJwJIhapZaNUIx
PXXddyYjotVbPWgHLBdKSaEA5FSmayloo60ZoaVzhGVjIxpQAHfmd4vEvod3F30gXVklOE9VZXOt
64jKgF+AzhUYaHyzzkHo0V3ft4hExa6uaeQxCoepC9GheSvXAYH9uitBCdGukgRZujrQeK/eWiZS
GMt6B/bR+pE/slY0zUfYA52jZG6MDddHXMnePFRA2lXeKds45tAhGwgNF869LvwK/9KWLtjwQIJP
Psdn9tgd366aKrO7jUj7VhGJt7OGx2WcdIXihiwVEaSNA1DlUx26iz3amtx0PFcQmn9WzdfIkhQz
u8tVgcFGTigu6pbi2D7TrNsYhN4ht2BrSa1rgZY1606OCy3ih0GWHkj7ciLCxudSsKZSb+ew7S+I
6OmE466AprVAesAptAvWhmN97CPExK3tM8hDqa+7kvw6xJRJ3IoEeLBzwvDj8GAlY6CzkX/BVCG5
Lv4XOMPKMgvtf9GHPzqUi5/CtsEmOE0vaqPJAfDrDvDZoPGBz6IuZ1PgenfHegSqbPV57E98yOZb
tGyQpcz9TQiGMk/r5Jpe08osJ6dQpiytUWppnLYoeeAt7h7oN09Mn6SH+fSMbiRQuMnrkb15O3SY
03W227fD2rjOSVLYQsu/dNdAKoSM5abHHxydTAJaz6q9QroPabI23NKiY55hL4qnQ1kwjvNJF3ah
TyqG3/jE1Yq5q/MJsoxMA0glJdPGeGSytU7kT/7ltQOhLT2KFCFZ9CoKfDXvMeFFLTFJTIxL/C4d
KlMcHDEQmR7atOdQq1kbxNEhzjn/Efv0ebjY2WaVkWZ7xmP2mtZN9NkM9vFkdj4J3IYR5E+1tq5y
sYK4uI7q0d/7FskuaP/H8S1nf5Jr7J7WMsJFA+KZ4rzlIQ1lhILCBBUm8xSv34/au+F/B6ezV3Cj
2KqysaTeSGZUgAjr5BKFQuiWd35eeFnchztonKn4cbvtZYn1ysz93IwWgDvjxHeJ2am7PaRTBVi2
1VZhOf10tK4KQUOXusxWRgRRv7UhB7DXi5NxJ1q5JcCoW6LPcSiCKxRb2r3g7TWzW2/grGqjgrEE
7UsLYd+rXfHbu5/Sl0ufvwm+8LogKEzOjNxDAejeMI0lJ5eg7mrPlaCHdXrd0FaE36PMP27lzpV+
ps7zfU/9D5QYO9BpejzY2V2WuvPTs0O+EwMPKyeVodKMb0WQVBAl5mJGBk3W6Qu0/LijnvGP6oDU
EduCeGcZOU0VR1pEwldLv4D0HVoYiW9QVFFjONEXQTdRvhC7LSbDmZaY7fMdncaFBc2/9d5blb5A
5p5sTYdqsq82562xNYvR2H559NpJf+xbby0bClYsIhkUMPJOTId4HG4BWwCt35Y6Ev+o7KPUMcB7
Jk9T+ZoAgEGSFeltXetgZK77lUxdLzkv35gOzxHq5Zlg7TCf9cYfh7PNdRQFJW4SLmJIraH97Cmn
uAbl7BFcEFmX9REtVmCgutGoDIHZuTlpa3Kor/QcFHZL0LktZIRq+ES4Em4AABwJLg0ViKXEI7Xn
pqC7M/+SPPp441olsgE4rzKfTpEpZ4U5tX2capD1szCU7u3950oadgs6/0HD+CXWhg4yCSpHQWHd
2dDE10xIz+/RLegnn7de+hg7u8YY8pDHWwOYEF/228Felax0LnyJSHprQ4oi4UFJASiahLx2mgJJ
tl79a5trjtbeJlS4KR0Hy2eNZe95uYanJNsZHYFF0zmauMugZfRux5eGNGH2ROQeiP6neG9+0z7N
KsIRfCsDuH1tVwLqYtZV/2ycTHtV0rJWeaQo8H6zwZ/ipnmvQVIho+QCPjEok1tUM+W0M3tM/qfQ
IJvaDSuwKAVxZe1Cyav/h2KD2yOdFL3j3PaAtYR6t7J4be/PWmq5PMjKG05Tz5TNcdYALKpNAOXy
AXYicjP+lAtVdYhseXvjWkE5beeLD8wD/aNoEj2z6Ni1j3qGOA9ts3LLKN8cw7cGtSzbpA4ne22G
NfjnG3CMn8agzMl3CW/x9MYO5QsMyKKafuuImbps/GbnLgmB03L+A7WFcQ29hDDWPh0155eMG02I
8NoyjgbZU2WV6ih8nK0rrOo3Uq+7kzdeGHPnfyEwAzBjm3+kWeEEP6XxUY06JLel8DNDDm28ho/y
S/m/Rojcv7+Ms4le4L9gpKA2MfNyIOV7yzswsBzqJSeF0LYSZFVvhvo6f8COneL+7F918XQD6JzY
hYQ185q1LqmaX59BDXWBHBoCb+oqDb1l9szg7JFM/r7kEISa3mccodvoeWzh7imsBS7ytgvYMOUP
42/M0eoBWJK+GJQJ20PcATkiyQmrZ2OXT+4N4mLO3XpYtqCJCI7ldWHgrMACYHwE7y6HHpNm/eZT
QQVe36c+KiSrWPvREacjYS22goFBardMcvCgxudjM6CbfIiXE27Qyu7PsDhMZKd2c5heh38N9FJR
nESlWpYVEllIQ3owiBQ8PLSx1Siu5ClwxkjBHln6CGyOaQ5ejbm2/TTUQXWdY7os/Dv1YlqFpQhi
iqaazjN5TdmAxez6Q9lxoIqv9QlSZ2jchGqrD7bg9Pv1ttUO1Rk4SSGo35PRNrLkUW5M26WM1+YM
7ggcDR9NugwQiyfBNXoiJrJ4LH87DY429KAooOhXCmDBCs+7/3REeQuAtt8UKgcVrU1aHVmQ55cn
6+OnqBO6fv2gB9y37ZVRVtgcfCiQbzidgOruSQmZsCUQmkzXe5IqRtWUPevzTZcofgt6l8RMh9D6
M9K15kL3P4PtpQwPwb43tdyjfgIkScDyrx/N+AbvF1Ho8+9NOb9M9iUEIEn9dvqtUyeQN5a+DBSM
LiUu1eWREEr/MEbMbADYUkdN6bgVmhH/MJ3VrV8zE9zbMnDCfo5/3+tNxWql7VIasQX5h+Y+5mcT
WrU+TyZFKmyo0Qfinb9W4X5ylUe/72YtOILN2l6zFY1wLSz7DVyzmTjo9jMEKPRJhIejAb+rO86R
834ScMsqr3T03AdSPDcGJMazIimnr/NTc9mgIlycaw/M1KDIDBhxdtIgP8MS/yNrG5r1icEy5Hm6
1TUyuKgw+R5dlloYiy9mLJE0OcvMTW5naipRSUq9Pd2K2PIVvkQ6O3FJIZ3xP8VGij77IgxOSvK/
myK8MgwHmWmQt1bbH24rWMmCHKvFxa6l6wys2T6v/+dKPiymqrMinB/DQpy6ZtCnVOgRy4hAQHf0
0CKEil3+dk+C+zsd+YwcmpVCxS1bmTkqMu5DcsVrQ5o9JkcnmbK98oZxNxsTNXAigutmBTNEaRb4
B9kae390v0Vx1h7SvcJ+bREc8tEepnRpaT5in2t7re4yznQMiXxFZqGVZYvto8iZBx3C3wyr6bi4
1yTCDO2kJwpCzMeoXBYNMwj0g6SSxQZViJVgs/VKB8dovnLAblnZVRjyJq+RMsLCT05pv5lfwwE0
WlIgkixiENrTpovJ7w6pl9iYXGw1WRWfRNaW+t42L9hVylDF5g/Wc2YtUC89L1dz9A2dYnQrJjZF
ApUIOPXVRaUs4juI2bof9zyKZg5U9huye70VSxQXWbp+k8kcskl/E9L0veFCUWXmYL+ft5OPzNSI
vynLSzxbGu9DkGSL3mmqBk+YE4EZ0XN1vmynPMep0x5K7oP8CT+xVWMfldLkEMmhEOYr0WeLbFtB
5vLYG77LiNWfsx6zYmJGzq+bcw8p1QHcl7NCuCelTyjQZOQ1kmWtT4mrgE7YOju1XBiAe4+GA+Qi
FNHZrRPtrXQlAz3qmrRqQ9eQwG/0HpyC5/Ddt5ui3I0Dedl+mv9VSFXWGi880ePyU9YB/y8RLgJ1
QBTg+UY4unauYDwnd6dIWkSegmY3Qd1xKzYBMvcNjphsbLWIXRxXw6eZ0ER7apfM2T1SzXRpLYTt
slgMI2eqPl/jr80jGuPWvZEK32vbX3UqvaKJD/ObBPbkWmN9qSWRqISEvqpFsiNWR5wkUoUN37d6
+wYhV4pQdovCXj5tAO0TrarPSA5Py7JT7TiDBQAFX5w2B0cBzMZFjjVgkvObm/ijHdLUQBIWnbJh
DS2ubzKqoSN6Fu1jLS/eDX67df7gw5mZZbVd68Po8lKi+XA7vLOt6FH64ZXnmFGmAh1WN36zWa4t
1kuqNo2h3I2AKqUduH5khgFO+vMdc/qxY57WcJtyD+soopnrwdenWL7NW4+fxunqYEsUu/ykin47
dG6V5RAlCOqvNUG3ugPCPN1Cs4j0prfaIVPlUxdB/YIERBQHCwILKiNBZj+BenRWoQX+Ler47//D
VDIiOuqN+TkR0V3pQXL5sHeyLGrcF3Oq1vBG3BhnUnSptU7/TG2eaf5ARhVrpWUaxHJOjLtl4Ny0
+lQK7mUoLNeq59AudMn7GnVH2xYBQYimrZJ4CNkjXcaP/SJimiE1LIwcHQ40CEnNOzAV4OgejZH6
EeXtfz2lDmysDNhqe6lwqyoU6LxuCKr6egdafo3Y2S5azxo8xyhIzGHcff/9V6Dw7xEMaIQIb1mq
BoAiCueZkXHUW3UE3xVuTNY05ky0aFppFnsm/8tfhWSYvDxchI3styTsWuNP83u8uJt+r326jKAo
kHD0UZXLfvL62JJ4xoOjfGywJLSYq2MMPUH0On5xEYnTMYckzZnd8enKZUqoRc7QlSI9gYX/zXFa
5l3a8tqvAKIj2Gg75utVimFFlqOZh+OW+HBswWDmYQDZFUdvg/2VHc1hBxhpJBGjj6vmN24joF7J
FdfATEAT3ronjurNQYV6Z2OqARZrPqKAhUmQ06mHuqsjVtqyM4J3oQEbeuIq0Oo3zjEnZDlTqd+N
Nr1BIngBEl3oYKlLpyQ9stMLArtiGqZ/ZOSHz71f6VxDqGVULdfDN2/+8teLLsiPWSptPKk4S4nT
OPcO7hs9wqteoXunWGeQEIJnuJOSSFEojHwpf/SOd1p6zSpb6HfDf5GALqbSk6teB1Zawv22x85t
w9OpbEu4XF1/dlx47SKK4QrqxoQHhv4D3huxnqF/QqlO/7Flrh3sT1Y5ZbCG5xZCzwCuzbutFe2/
EB81/Axjlr9PNue3snHCmRaGOAgEh5W4hUitkzeqi8TCWZFXvEPZCoUXa4h9k8AaPUE7K2Tc5s+j
oRvHdKvlDCQLLiYY8wcdwVPnf6lTwcUCaQF8Axc5dlEVhyEpkj1rKodFdlqhS0OV/fPAzkAErTmE
1dKVb+zDYwL/zMXGd35koBbR/jzxaVwqAZG03sCSSaLaHloXlYCsjHm8yqud9HMeLlin2YOAgH2g
m8KvKz38ctNioUPbpZIORAZMF1TTypSiRJybCoejSIHruqsQqxHM4V9JyDlPEjxbyMLoVq0JkVVT
/pXqfbIBMpNWwko7EPw/bF6Eza9KOyyRPk0UO+XfOzf860SfJqF1Fb0EqyO9n3M9IkDmRIEAaK5A
hTl7QWvbZnbQqyHwmeW9WdeOd2bTSSGXKdSRMylBiunNt6UqI8lsBrmEnIQCmmVatYfnpeBgAbPV
zXwHOaD/XpO7P7Hsdz+Lkx5CNOUr1kxZFkW8wx77YIjYwtCMFcFNKKbCiagaNiAbaSx7DnVMop1u
sY0Z9kUPvXySMgEWHS/ZDY8iGeqIVXMSHcpGXQitMTv/6qw7lLqo5xff3T1kE4WgmZKAM+eQzTjW
8es0WO7Fdu5q831xpFt10PjJ9qsFVAvBDFvpEvEGyet8D3DjTgIzAYvsV69Yb2sZTw4aFqUH0GRP
Q8OnPHhr9P/3fHine0qtSUHnJEAZSlulxFL3ZC5QkANSlcCSUVpE3mZF54HgqFH3dbRoh3tpLU2T
8ybQgn6epoAqnOZSvqN9ct7059+HDDqhkJQOmSm/C99u2DIUztjKjdGzA+ko0HLj6/K6SynD5jTF
JZCLB1ai2AjihyJyZMt9wmZG2r8ZqV0McZAEm5Sd8GKvIWJSFuIKFc7Y/s+Gwx4UnEek1KIFnPPz
9Xk3rEQUZIFwxrkXCsZGYH0fyN4JkqfYF8MwRL4AwXfHTczGThihoQ3fYg1FmacUSt43FVT51jNU
nZxqFzTeulldKPrFhLvLxiKjlMr9t2qSSW66dAPMsZjeJzksudU+Ua/B6qarVCxkQXAgFRFCQRl3
U9JOnSWTfbOjGl4PEvD6VthzxMeBP5O/S5J5wvUyujGBMLLs8MZSQy0/77mjwl6gKwmlA3CDq4Sj
9QGVKt/JxMAIGtXiwiHS109/qTw8Is26KTpOxrQTbrSN7VhriUJE5x3JaXDRecr+psQpCiZ+WG+Y
qncFmxt/1Om+A5zpB+FkYkkkpJVaR44mBh5TCtGQZYTGrfaHwITB2VOTVIzKSOfWf/4AKsY0ABPu
+uXCgj3pOz5nS7X507C3cUgl7YhfJtNwH0qr8oyr4U9MuAN/Ba4ef65HFj3llDKAVFqE1d1gzj6l
pD3dp/iwsly06nvEMjwuWf8F5r0SuyZFXN+Fzf0NQqeFGmc3DuHu2hg8BgDr3UurrZ4kyktocyv9
ZyNh5Z70N40xsOFsBxDudl80kldQ5Pvr85LdLV2kE/uMB3CW+E+8r2eXHFYm1tTbvVOjh+1hDMQL
pD9WN0CVWtP59WJTflxacSXEObJrZ6k59NNLk/i2iJxLNuv1pFQJGxTaCf0gx5DcH/BTuCnZPwKH
FrkLXfRjg9Pwbi+ww3VFgEanFU/Ih/GSxYgRvNSEgiHOxxKeRk2BZyR5nBR/YIdq36vaWtWyRZH6
S1z3nBHQchyaxYbVjT5vm0/fbcge1yImFIF/duUWPUg6dGP1FSjDy0c4tEZMiGypqO9Mf7qt3seY
KFEK+9+Ba76XQL2d6hCrIJEFEkb6yAw6ZYYxk/0dHr1/Zo9zRaFsHXCwMTf+gVYCELR2H3kh4XEW
ASG3gOcXRfPYsSbVivaqeGHczsYo2hjxBg4gzGIzQzeY/WP3fsC4QUHKdJlMLtCucb7P9HzCYHb/
3HLnG6CTPEKeHeQcAhGSic0D3Tcdkpbrn21gFd9J0aPn7jo1Z3JH9fpcvvSAK4afAWUESbWKkjHX
5NAX/5J/iMU0bDnjUGpb4tPq80Jepvo6RaMHQCHzhFOaiCjDEoOc54sM7iaNChgI/IEcMgqjNbZx
1rIB7tRDakRrTXFo5+n2dKpUOAeEs9dTxUt7UWH2InB65uUvx3Rmcu4tvUQrL6SnemJkKgIktCuY
Mx4dTi7N1r09goij1+VXD4dGJjOTBuVYHBOz26b1s7YIGFKAWt9Kb4Lp+OYBx1b/pQA+LsPxj0j8
9nlAUYlbAHHA7fnXvPJB1+IXKHqwHqnqQXFrASJ8IoK5dVNuTjJgCP6TdRykHvvfpxgUScargzYP
J/ER6nLnUjGbRx1RAtbU3Q41mS9JRdy1IlLsE93flTioyEZYyNgONY8KxeR6f+sHNvDYw2adEQP4
jLoL0NehqDmMNZEux4SI+BhLYTDHy/o2tZek31p+C36SSsUhwJJ5gI6gOcDuf7k1Hizy0I7b4t7F
KmLKgcLtr6wXD0SCmxmOoI8WVWMq1SAW3N8Xa3/0osD93nfaZ9H6KHOCf0gEYO5R9w32gj/M3+sd
1++UlIac3qYk7E4g/A3CwRaG20rAkgrzbr25N2Q3e/lPAgzYDg5mlrSoiw08atrRJOGDyS7fuO9R
KNW6HCvvF7jR07IuKWs0W82K5LxFNY+1CfWhFGNVc16Wp3r/W5tb1xoUq/Urwi8saKWOOc/rKNyp
FoQG5SXk5Xx4EOg+/KX1ecDZr/pZF2rPHFYM2dqnUSb73GDI5o0DAsEYi6coxltq1T0w/lRNhBRJ
IHJz/mVWARiBJ1h0vqaU7Nr4L0pqIhSaV2x8/Cf4DzwEotWTJpNwu43aYFEojeWAGGXcO1Xr7YTK
lDpv2B8pyp9V+mQbc+nsDdVP67QGQmKHCWpQXUox0QvSHLfIPzJppwSgg14TXmrQsSIIdNooNyLe
aEvUs33eE9AQxFkZSkrdW6nU2OZF8wv2Rg/kUUVGbvMevNFnU9SOSrgP1oYtKEy4P4eln5WP6Ced
zkqAW5YcDH3y4Eq/6A3nEluiuXegdBKCf2+ARWVdtLNe+rfiitnmbbuyIaNzMmVGCqxoX2CDfASx
j1Aadseh4UlaTNrlWACE4Awavo4MEjhekR4qU8jad6D8FqTi9WLqNJotzJ7GJKd0ImIg1F4xalWL
apBC/iz8asmeN05XvTe0586D7ZtKNkPzcGHsmofksR1NnmoNQEi9qNv8XKlkCW6J1tkrCsfd3PA2
0XwSM9manliIQ5tPtHo6W8B9Y8i55jkdc5QNtT5DtJKNtIDFg4JdaybML16kVYJehvdRk4M63tmV
UG18RQWffgGNusF9mZ//4g0rah58c7msq5BNcQS7I4GyZGZZjNqv6CwkN2nLVPhCZbuEpM0GM6Nx
dEiLcsLKVW+TrJXh8ssCgWTLg7rlN0FyS7XPYY7WXy3bsczrwl2TEXrvQEKn8haiVDMPKinAUeSh
jVIKDHImUFDIstFDE/gZTE+ZU547RH+dqLBISAaJpK5YB4MOa7gddK+8AhbKPN1RvPD7Ib9MbEiN
GNQcanTxKOG/QhopFe3WIjhD29bGTI0l+3ubwE7R0EPSp0z2J0O/SLa+W8u1bvy75SViOL0eAaci
irZCY6hdjKNLusg+hcTj8Aavm9C1XluTXTXJMn/qAMCwq4U2jsVW9ryUUHk89vqVuXv/Wa/5cECP
cbkgJixJ4bHyOknWWUFU+8y/Wu5dwv4FBdtLebi+lwNGtxX0zIXLQCK1/wpD3vqsuLFa2QKUssL5
GJ4hkBVSJGFtKmdw4YZG+6g848dFynEAAiAdjUvrAgoHIFdNwOWM+RADOMNk/Fm2WBYTVOgQtUuX
YieTHGTjJ5l0PoLUL6S5Bm7LvuIQQZPlWAx2tKcMsfivZ1CHOn0kGcjREclTkIXADRkuJXSdmQpo
xWv8RsM3hlpHyIGPKKjms9HyPp5yMXa73qGPsgK3/dTiww7oCTkSjWOP3h7wKbo8ysb0inWnXkE2
dmiuxNVEuBaDGChs9ttWg1NjI/04LiljBxWdRJNumwQwWTTj813vhSvLfLQ1AzWegDMfu/ofWmNU
94hPkBDlYE0/cuE7Qe8l8Ak8prAYbwvSJY0w0HxTr9/j24xd9qVgCi7PMsY1oTiJJl9f8Abi/Hfc
VyI7MrwLtT7/E5fXaOgQY3lXGAFsNN7EpA4zbsDS360V/fLHHSbhOQwoQOaN/Nd8qg+FmYGhFVBL
2wrjB5FDaSnIPbd1vWlD6G5TVxLAXdJW+STIGL0bfk2gkr5xhL7XaLuvtJjCvBfPa/NUChcVGTEM
eIm6I3KGMdmJ6HjbAnIP74JBh3WPGxoy2xEUCzDO00eqCmPuLcqbgsxpbTMDtrcDp/xm7nEhVPcW
fKtYJvVWUhH1e/Kgwn+h5enCzhGREMRId5VbghZ0gTER+vOGzZCH2X34yQCVuUSqABmNBrMtiOxM
4ATO+/c5xYWKFxuU7PA6cSU+xWSrAPqcTcKePDmAxGxVwZE9UjHIrW9Z1YqpRcu/LrGBs9RWXqFl
xzjbgWcW4rGR2LPYsPA/JcWqvk2TOqmx+R//pAnbiHwsna3vMY8urT9U1gBlesgWvraTSljt0q0o
m824PPUMWDT/Q6ThsPwg8uM3xmen+/XqGu1rPLIPSt4OIU99kMzubfUP71LfMM4eBcX1llV1AHX4
CKdZiuM0jSgV7Up6rCVu7S7VzT5QXhNCZ51NKnQvTh96A4FUBTxDkwnv8PsUxEdN9qL3e9zeaPCg
M9urjXGeSNXAtjdI+WaeTkLL/WFOdOmunuO50e/4qCVJnv5Jo7lSTEI/l4mQT06ZQasPqMFgCZLD
6tZ/A2Q8q/gIpKBm6nnrO1zykT76maSbAicrAkaraZB/3s8l0sx/eorSkAwR+puHnygSj82L/rrZ
7hiGUMU4uYsXc+KXsyOfwAabs6N4myjaPzIaxsqpnkud13dozvob1ShM3kR0Cn192INiJgQpV17Y
QG/xJK7rxDET5q2hGFmgO9RCBZCp5dcsbRanfU8twtbQIqrJJ/oNBeQy2ijRC/7ScPgMQcm6ZR6X
Ps14Z7La6XrWSX5IrPEz1ZtXfL5dkCAsJQYFUx0533K4gYN34A4C5N/hz84A36FY+IgvwN+wEbuZ
ZEi1sQ9kH8s94vgRNKEdrBaOiSh/tbItwPpCVyr0atrUXgWr4ta/jw0y+BLrN26kmoDm58SHGdSW
gK/JpDUw28wX/ACQ2xeIvXXrZ9EJB75461NFx7UpAW2rN3T8P16fpsdcQgaTSN8QweFmRhv89anE
e4u5w9ICTEzQATwlBf1jKY5scabMxjLwx8jIWSGQDa98bLvlxJfrx3RbqnRxITjeUCSxNB034o79
zphZRPZ684YP/H9XXUuAhcTUxoMj/QLmfLxvcoeSJ+gxhVD1tJ1iqpLu+UnMu8h5OhKiNT3N2HLC
V8Y47HTQGh+0elPstKYYBAhhJL/yzADkHPJTUdyBgI1v7kxdH5VWSaCsLS79tIiPQ563X8j7rPM9
UZCE1jCOr9bmkiZz8D8AnT0ozTWSflk8LKkI0YVHkaR9Qt9oI5W+MyymbfN+QEututBf/gFcnI1s
1nSmpUJ6fkwZdA9EKTynFyXedm8AoY2sn1zn6CGt7AA6QOANw8L0cIWlY1tDjUMUv7GqIunhdPQh
iYgQow2E8AFR7xCQukOpI7EY/VIlD+XX/QoSUmUNtRcU+uehPy2hIJnIvb9//QJIuwVDwIHNYweq
qCbm9X0g0bYNgZJP5fmSSCYSYia9cqySNqnnlgGhUPdB9f4WuD0QIjMIZT9BnssaJ7UGzyAK3YkP
nun5VIyyuajoNrPm2hqUvVq1tW6lK2doB/+81uJc0M5JrRML6+SaXPxrBCSd17a2nxfsn5RnAYh/
bZjRdMQjvcPFpWn4fBcU7wA+r2ehU9SovJfYBZ4WM2zCefJNSdvp5hs8xUk0MO8pfWdrDCYMv/4i
7VFPazfupaELfPlmSy3iBVS5ZK4uDONaPJcNf0kHHHqUPTID4iBTs3snfxYBpyGYtp1z0aFfC/Hw
gM9Xe5w+qxs3p1VqbtndMoKYQk20eeQBEoqD6IemNX65ccjZ359h4pxFvbTgs/LTDzo7QvgpZxEt
M4af2eP47MXD4UlrG4wr/SpRJ00bF5tlSImFt2eZ8UewDUzdwUPyiTRwnOc1Ls1KXOa9DF0OVN9z
RU2rYznNZdD0SMHq0hmnnYEsnh32LGl/6h2QlpykL1k8Sw4Sy9rav37ShvVX/6XdimvbLEHR7Jef
r+l02aXTk7dwQAbcS3yQzLlTPoB5+pFVnsamfK8jpjHDhWaS/s4leO1VRyiv4fLDAdEFfcDxLG3b
dhQNZSy9yBzwqXuQbfWEij/23IhKPt64kZqwmiBu3rBaS510JrVGX94XZBD53Os+2po7Yy1y8bKP
2tagK/XIEtmAy1N2qUn3CmajJ9CnB0l5aAdL33AhWvSlcRp3IvIEzrDVyLdPgAGeCeEr5G4mCo7T
s58uS5RYGCfCfZ9x4lMC5x0fyFeSgkS+dgFfwh3qYwV3prhO0Nrx13tgpq4w8ULEgNNH0/ncFOk0
EFMdpE88HtfhNI8FD3FBLCNyTWLLTIHrqumTFviPfVdbJ+vCTxyadzit1GP5jm5su2hO4Bvzo6EG
tVv12HDtaZNKVm+Suxj6VoG8bsUnT/i4Zvpk/t9m+xFW/gGinZonjDcBsh2q77FzfV78I05scW8s
bSH/5PsPmuqBgWmwAi0tCkrTiIOQPDReJZlgoNmQ+6+qdQBoC3TMZ4tVoWdfXOXFpbzIReOaqbga
p+wfJS80Tq0HKxT4LRcMpOhxgiYIT0W67G3YiWVEaFRHRmAI+8+BoWV3nH5bcaqVVSU4LvTodFec
iOPS+TH35E1pEgO3mZzVmFQKhRYPyJKxN6x/6OpUHWGheBdWBqOWE3LJtN/FtjzzsYKmPz0BaVn6
Sy2RUGevZfFtcQ8PjN/UiFfZKl9nQCeItVP+D7Kv7ur374YUEAopyKRe6s6m3TeZNpQKyh3sDnJY
U0Dk0rjoBjvzAnoGErCWDaKIBF+TdTiJTiSmkkOquDKyZvNI69uS3pcSXbUOdwgsCLEc1OilDfet
ybMtnDYyNecXqDx85hQc+bZgpFmc2NaH6rL7eNVJ7kcOMTDxbISWc25kcmhsfqpMPXNj0iSN3dCn
z+Q6AUFLJNj7Ix4Sw7c+BDDcIzmsw4AUYgx/jLgnasq68R5ok+ycIdDqmQU1IrlPyehnqNY7nAOD
xgxZ+WxXF46vi81jIETPzXz1b3WeUcEuapNCN7/bSz0y2gaQ3E25EC6VkbenDl6fx13Y5NF12soO
LcFvS97CBNPix8Ea1Rpbvvg+38NwQDpAP0ZUeOqHAEPciRLT74L5ozELxpVWDdoyGM3P+3r0Qd8v
bG8oAr8T8IZ/aPtikSWEPN0HtZYhvDZs1fmGgBk2Kp+f/0+EpzgwNe7tMzkD3F0DkNfJnlvk7yI+
WkkVwDf+dpSk+n3W3OzjHyP/FwLa4pObkrO/27pGpucjUkaYQIBWVK4iJrDPHW8pxqGo93u11oID
YSTYSmd4Ssfk7QEOe7OpRlX4fRvOvMPOrtpZo2b2EnWr1wRiP4sKiDAlWj8c8jP9g3u91xjOgCYl
J/8d9+W2tFHr7azuURRj8EqYcmkLEE81ILm97dMo/nLQo4NQnqDw0hk4tBIlVwjngie7yA8fd3Zn
8nYkAEPj10zieYjKO+gh3JOlMMVhx7Ul1R6crUbaeFouNwbzvm0+usatWE+7Fsp5gW6ACmDvbija
dUzU8zjoukuwqG4B1HUvlmgiI+PrIEXCD/AxgMhC9HfdnYrIqwHgo8Euh9klj1mDeQp5Lb+NZuh3
EjUHwgZj6+XCbr1JnClbO5KLjOmHCwFmyeuVJaeP/gbgr3XAyiy0fFXGxmhlcR+hPpbrp7RTNS4d
Hz1teyt1rq0CS+z0xExglrnZHkE5iV9NrDZcl2cdW7ltkjZgMVabHZj4WsA7/WWuaNXDB93nzxLF
uyVSGRBzBPRfwC6VMhoT36hJXZkZqhWrs821O72F+Zl3XKYFuch8EPv95/8iz7pgAYU585kvnBmn
3jmshkDgmEMcJH2aXoDESgUDG0UUtw5DWzGdE1+F0yv1L50xlO907uC/68fVLP0Tqx4zhBXUYgds
MR4Vq2UuWh78F42KtRBmkb24Jb+Hj0br9sRK9407pH1mJkvdc9jpEcgC78cthadwT8feZ68uQDCI
/3ksdLqunzz2t1HSTBvCfO4Obb0+NQ16HjzzF02zneaG0QqdZaNyySDDQM5r4WZT0PHRbBZYjXTP
yXSys6D4vpTYL/78KewMUCOs61MG8a2DwKenXWeNgaOeb12qpnmbW/ayq7iKa1twOTStcyqQtEK3
+yw6CJwVIA8DUDVS+BbaS2CSvc2rCDgp+Mik0vBK84WBJBv/mfGRtbkeniK7aerAZsqjoddtS4np
qIzoBYYtTLRPplF2BAJWK/Nc3dBjgkuS0roEsDSjWd4LQylzoOHLRwi0CzPCdUBHz4XB7LCKFjVX
/bu0Fe3sDd56IcyPTLunVSyQU3LtkEcSjpwbEpEog2coOzfs69QBJwYDkAuT/4QZP0sqd3kx1XEe
+BbPdprzZ45NAr72rMyBg/QmcwVhQQ4I9B3ELK+JYsf2BpuIj2tCV+D12F8QAc9PCKWnMnxThtwr
WsxPKftT31igWr3ieS8IPLuprR37qAExbLmc59YZlpqop3BYHEYa+a71ddjYou8eQv0LCuUEvflY
2p9lNusjN05AgTxXksBBbxL7DfaCXKRnuCFaCyJY3/yLO4H0h+QAYrenGsfMJvRbW1amgsGb206s
L3qAGiA4DWvTuIfzDFK8SgP4DdkgmlZJFSPjvFHXgG93E5E2ImhtE1JF3r/JMN/EEeA5rfqIp2+B
xQZOW65pQQv65a5BtsmPiw0XbTVxXpkB21UNRqAhKpKmyLhnFv73VHMilr64mrlVr6wPuJXStU9/
KIVak2ypxU1WPIjT2aAlUkUqms+H884mHB7+grZMwuGdYD0i8V1YpOm5l6YGOfuyoKKJOQLYCwvQ
Y/lPUEQ8nmifedXfOpE3/5m4R49abAFbZ07YcUfA9EgbDW+fOId037LRMYX3IT/tAbHtIWptrLXX
sxJaGGOdEU1y59zBumBWdgOeANs6KkaMahP+I8+jcgSTy8s6YhsaILOpks0VqH3d5qg0WA9KQ59b
kFnc7NkehrBBg0I/g2D81Bq1U00ogdIxXGGGote+yLvNWkgqO7ih5WHY8uwImBKTcLDejeecgRBq
pEObgtrWUBgXEvqEuVrdrqTd0HQlGosmKg+om5sNN4CU4qWHHpkJy77LLHKAHS4wCj7fF3Y6ziXm
6CNtmQBvb57J6VdkX6cgbIxPeN/05c3NAB+KaguYtOZIIyClrEpVmXowB/cfvoXccD2CFa2mFJJ3
D32M+HmKHXDQOpfMIUlDPfP7O3JCTco44gCtSRR0J26KSkfrdNckI4XjZFBFO1e3i3H+U4j57gqz
6xChpaXPxM2cOoUuWff3d9Jokdx+JX3ORjmLcpsBiGNjfY+UW0UmiGcym/Hy1tzZwTADhbI44o5s
a7/SQkkM3Ikn2UBtvMGRKJAE/IKx1npiLou16cgDq4iKSaFSLUErH8XcNmiOg5TTJF7QMtrWPN05
rBmAU4LXdIem0TJuncS4D5aNB7Fgsq1Jf71bvTppAOOEl6ZlTsx5SNMqCgOhJ4PDKzem6NjoV+T1
awSeGwyjd3JcOesuvH3Bx4qRoD/5bx1bOTxIkRGTkPZCyBh+yS9k9Nwk6y/7RsmqE9jFs55X6LDy
UXGcdpPXknuUd0mCHysXXp97ICxPLSZGMfZz7oHVxPBM1KA+94WtCFkDU8kLZDlyQh2KneeeXL+D
skbllw5PMjieRm8aJ2AJ+WNUZIUcG6aqL0VNxXhsw1s1CHyQ9Foug4W117r4hf4btkwk3uPzAwYV
DcTGczeETr4u3FAMdPu/ZRNeqwACBaWWyvFxWmWt/QjT0ioHS0J2I15eIeu/luF+isqUj1Nmk/l1
PCeIoEvOLCF3Yh5x7tTSC4FKemoYON5dWodGJJM5AkTEUAAzqI0VO+xvKU57Jje73inFkGgjnlO+
54B0f9oxEj8RxOYujRgg7x+gPXH7HfMp4y4FxiG47WJf8MA6OmKiYwowXmDr+6dB9J6zgHA41q2L
vvtjs2MJkzguqJBMyiFZ6gdjq3MAXPPp6eyxhxLKZ0ZrurQpD9uGnuuQF4atmEhtCSZbBfJXLQ9B
zUtB8n089lkUNDeonuelQcctTdEDObwrDdNp/9D2TotMdfnLI86Qpfl4h7oCFrzOOU2/1dq8b+Gs
DuM9EgujEHIA3ZJQkI0bVEVNL5fSNE8jq3dJ4YX6kyWC+j4xi8oGQCXELrGqUG86fzuivIk6gYZT
j2qigGNbM3KGlC1cGy3yuSTABhvU8ptga2AUxW0rb11mjXo906UelhgYV+Pt7a2TwSt3WCOb+C0r
5SSKphiWl9+vCdV3HpKTloZvMGD8hQoSjNwj4cscRXuP01BXsl7LbxgbbklTyidgFvmnP0uzpSlR
4VfyKHMozzmiKy8vqHjN+wWuJUigQJy6N0jVzZxnMcekcweSQ13EWyj6XaOztfJKJbltmtgrWvTY
MZf08MDfYB6VQ73Ze/7rlujXPS/uRieDe+n3Tt7rnOTtK7RzS88b7s2lgTWd3ni4ev1i3i8e4MVQ
bico6BX6kST0CoMvvEb7SR8zP+n5lwNkZ9cFvSsG0iRc0Bb9dnWzdSFGdtp55MqoEK52nemnMfJN
Wq63BBhgXZ+Ndw5YSucpRLkcaufzDgjaUaVTh6wH5U67QbMecjIFMjWd7mKdi+MVeUwA4QKF5sua
r4reRH/cOBMJYTWg9zpBWkmt68//BPCNk7WcqU9sc2BWRA/epbfU2RJkizkSuE3svoi8tfIKpw0U
P01IrZqJoPvtojKWE0SPm207celLNJvVsPR4PLmsvQgQf5dB0ZtURjSAy1s6TFn4m0Z80WQRMyT8
r4m7TPM0Imd1+3mGqBySqwZsQvsS2lx1N7lX1WE2dXx+OglsH1wVuoPnju5/p6AqSdcIL4tYCbs1
0G3feH+rVdVNCqvTH6oPpoy7iyrHkf+hj4yLUE+J4EtKqkU6tsPUCattn9EA6yYsBdNEsQrfxdq/
LXN7AUCSICGR1254Se5Mk9hlWPlLW+6kuOtJMzo8VDt8lx2yRV6NdfEPkg9Ee+gWXBAvkH+FQ7va
/DzJudS7kqqP8hyDQnFH9D9fUZoEbS4yoQ9DocFja1RHlqP4mJQ4bYims76YOpCpNqvZXPfuhjD5
57gOFliFooJmQbDBy91Qgcz5nMzcHhpDo4WJaKqlisgAhudzv/4x87GGj5WatpLvVnULFOh2HW/Z
tg10b0Z5jddbnBlbc3VbkLwa97FAJPZaj81RmQz55u8ls5VyzEYcEUj7cF6DOrJN97w1MWW2fUxP
5FOAY7v6aVQBgsR5AhgTvm0iY9st/gD2o/qhfDYIt6JC93SocIZoghwrH5Yv8XySghobIv94Awhr
WjUGvdjqrXQSTLIXISgBoUctFTfISou62fAjeFXwOOb6Mv9B7x31KA33u5hc5svNumPudI8Z1FIi
YpwvamsTteKbRWUaK1PLS6ssCfQdbFxJwv2KBCK1ABC+RjZVFszndHtLsuG3afwP5MG43LKr2u37
XVpR/m/cQV3u+jLuICbIcHRztfvdVszCurfrWARwVOpKlfKZFjcjHbyy3pGWe2JgHEeCjcb9Od2M
1U90VOSe+vE8BYCaU2E/CdhVSnJgkuwJl6oXy6uf0XqighBmCXlaQRNnGxZ0rFDRWC+Vzt180mwP
fc/6cksVDU5EVE5hEZc7znfRdwWKTddBvvyuYNA0hua25im5sMxqJjZaXavPMWo/3wt3T5RIc1NW
Yg1Q4pPck3Vi0VZFv1fvslQcrUWsJvv27umVIcR2cmnc6o12PVuEAOlRivMeGS8Mgbv24dqeGm0D
DLbi+UgCa8lVQ64GkjhSqQqaaejxVkvZ996ktnO6sXwcLRyTKLSyEfQQl9iEZeO5I+Z6UUf4eIWU
assenL0YtBdaLkg1S1Juf3tCmXyRUWNbfewMN4m4BO1Akt8YOrFroGGZg2GLjCyO2hrT570WlO7y
OqAlMYq1ek9sxZz8jwC3CmdR9+icGwSHeq15qde9evSL+CesVj6mr+BONYceSICtRxaJ9mkZ41D3
19ed3WTCvs/XbmOCQhhU9r6KBtOwy+9WGVN8hXssrVXl/YEGJq7yt7XG4rdt92UsPyW2f/V1ErQ6
AI+6tgzW39NZhzqVu4LUI7wa0bPmqTF2bFpVLKJy49AyGh+2Wu18FyAChsBwJ5JSfuzVHnN07E5Q
PyFetvVWPb3DvJv3u0LtyFRR3PMPHu6DbjbAfQ9X+p1f3xRx4UE6OL5Fm9ZZgfQUGFTeaXAwW8/4
AOYSVVFXxyu5eKGRMIjL+F8Ez9aEj43iHRr1qjYPCYJVaNlzzTWvUkySXybkqOyCRwg6x1qt4n/R
Yz0UYEBZeB1tQgYXljbKI/9rKlSfmtmEI67c7uK3r8Bt0TvO5dmFQygy1PkLL4EBbgHa4a1KcKrG
w1s4E8XlqvZMAMZuWvhIpCGgWGxo3skGFGzu96BJ8VAu6DOe4B9LOtffYAMaRjwqtQz03cyWK34x
qXxE+yEYpuyeil9MR+lRKoaJWsDmyElIJILIW2kLS3kTIy5jtu2IqnsuQBVYMO+EMpJv8iupSbET
cIHLheo1oCAzwVomAnU1z3KXOinLgof0o2J627vF/1EqIx7dyJ4G4X3wIONI9mfCFpPN4pAciSUf
hQPF7KKExZ7PD9E3YYkTzg0erdBdmwkRcMfQfU1mvxZxXhu/red6DCgrJy261zOsWT06w2dGCpvJ
ghoPEzw1aW/1k8JdeMbti436Hm4j9FJxctAJHdUdvRoxLACaWj0EkxvGRQ8ZSI70m6CYhK7AE6pa
7wJx8hSX9g9goepJW/j2ThxtV7nLJrC7aSVDn25Bn2jMkk8eDqW1gRcNYDAxHqdWmoePfVC9B1L2
5SZCFDYvGut+Y0p/W6FIHemkAfXx0NKclnRw414rTmX4Jlc8UoD2UzcpQ25GYTMy354f9RoDXrML
8Nruzg13yy0LnS+O+jIw3B04nz7Af5u4Ap+zZbLGqVGFGK0Oh+eJHbxs+mJ8iRVzByDLnzF3LiFe
rOoTk5wRHMVTR0Fgpwo+1yNoFeYhJTC5Sw/wM0mbrSz9p57IAVkohHtEizVIxg40ZuDN4jZTFQC3
dkzk1Wh8n+yZEHuPJhYRHKSNPsp9iK9jiumlSvFnLPf/Z9j854m/YUbYq2U5XnkvQQ/2lBkhRg/i
TUsAFDwebN3FtdJ+RbwxqbjaQ7sDT/nQnaqP4peTRBj/Uasvp8QLQe1KzluUS4kkH72S5/X3U69k
YyD6+xEcLUHgqVKGtChBbLokhY9/IcuM9KhIq3tNARZtWgTX4AjRzTQBQY0dyyU6tbUj3y/AMBgW
9W251ZPeLmGNlXfbvbtBFLkOsjSgfZIvnifcbSEtQk5g+LlnIvE9iHncWalV9BxdDpaaHiJqA83q
k8Fv6Y8snLK4bU4IDn6kfAzXibwxDG9AmJcIzvPOBh027mXZm0cZsguiI4LgTjG3JTaYCqPhvOzS
tB0uz3nbD8RZYITU28OJMIIWoSenSSVitAjgCDE2nrQ7tNo1v5hKfr8WZB8B6SO18D2PSc8ma/Q2
HNjViupAJoqySwCzZYfVE+nd2KkLvJINal0WNHkXO9NTVUri8kYO1omfVp688HxJ//jBCIoOKIPV
/5nmSaWA5I/JH9gBLDPj0br9ZdC9YvnWQLHzJlZ3jlPySA2gDJ7pD8DYeBxX7BnWMegAwqo/LZda
qqM5xVSP6P7j8IQMKtA47pyep1nDrZBB/tnxnxgx4WdYE2RoeiRxxnOla1dJoXknrAt5nmt0bx3u
5j9oR13UIP25Bu3q4tKA9KnylEPGA7HKsIvqjD9yrr8dSNYOZyFNidRAtJUDhHWJspVfHPmL/5eW
/VLQUzVnJh5YxJJtGlJokPwWf4SEgFPfuqISFkHpEkOLsCP55hyn5rywRsVmJEuR8uiRFj3Xhw9a
ArQ6HXBA6YAd0MNkOioBXZ+6tOpCq6loCl69FGHMcvOOyS/AX8SjSWV1AW7EXFC4zmhdc2dOnLf0
oKO2nbe9sxnh6EEQJ9p7s6lxIl1hW0hnJmdEm7bcxoKpFOyyN06aRAtUfzd893NUrP7IOWpSJ992
bx8vVKnavc7L8CF704lOI/20Cv9Abakp/tq/qpqBYfUcB9m16d98I9Y9DR1swadD4KH7nesRRQRt
p5hc0g4mXstzO7nQkrpndKuVIZVxgONimgV33TmZ4mray9wF4FC456CVUir2tic91czZIPv9hJju
wKHnMigr1hSlmP9i66gA3eQE5WBYvHNeqc3KE9EYfq/vofd9xt29+aVrBvREnwQ7UV7LfpXOfGQz
MArfk10kzcYNLS+S5+rLAR7EteSVDBjC/PhDAe9O0JdxtMqxrbrtrN7pkyugFsJT37RR5b3W8uUd
LlSwrqMdr0DRX/S4mvWHvcl1ZhLCCrSZqUFDoZa8sDHOzGGyiFAD4NZrx8oOR9kxBclQ3fp87r8F
fAzC3LaM9k+heKOYnMNf7MyBJR5pLYU9hMNf1ja9ieX5DcphE9rVJuiL/ogUpW6KALsEm8FrzMmR
LHqzpxWD1GHAJf8B0jetKLnmYMoC3tg2+zTsjVDXN9fitL5hmrsZtcgE5lmLrSQXMlWYA+c41L/E
E7Rn1FMpPWyx1z3L3tF/oxzjB8SvF2f7FgORoFFsykEevbGW1AZ7Le32SxDdyFy7kyQALa5Lww+5
RHWFTJHo6yQNc7igiovXhkrUDXm1XNkJ1WEYxBQNUMbA5fw7blMxzcNyRLYeFfImXTga6szNsZs5
WGYqCzyGohvuhel8tsijkFYADzAVsKcVDHHId9wM3m1/5QcqVCmsTeFUa4uNnpAUMnxc0cPKhM5Q
KdG4Fje3i2BPshOCF/+D0+W2qfNMby4mA1JGgCfNBzcgEqGtRygKrNGEkKgekrlnCbW76Lx81/oI
qM4EinewGJ0bs8lkQIXvSiHhgKevNiDS+TrozXmHSyELxFyXSP38/HehDeOtdc9VYj6P9Pb3OPT3
lv29gFfXVBDoi9jcpRF4tCmC7Dnnjm7eb2ICeDA9Oo5JVr2W7BOa/hK+XpQRPu7aHSuMuAaWSCE2
iCb1ellckBNltbR6+uSuV6qZUf6PT18ArJK8hTU+oITvWaWTu45Ra1Yf1AUmP6FTTz1m/C9uFH7Z
+MXAjcxx34YCs2CRpne660EH+IAo92+FHkx3lM/wIHkR5BTGwQGrVVgIkT9NibJpTvaSkJQyspJ5
R97SrMjHMXcYZPcJFnVm5CaYUE5pCLmhBmTI+n1lsQpEIyNnC4THvh5RLuh6LCeDUOmW4ppuLYpZ
F/JJcQWlLXgIuU2LPTO8OS/kmzVP7tool1HhlHUzEyAHW/klLNqKBfzSH27HcJp0mBk5K42/spFD
MCPjLtal4qj6ED5koSJn3rl3Z7ntgLAL0H10L52PdAhyMUFmIn5h1XHAQpWhixMaRjnPI7buW40P
sb4WsqVqdu40IyFy3Bg5UULa+WHZwwo8g85wGTMkxBgRVA1cXJvXzjaDjDi+zTJPazR/DZqBCOsJ
K2NsSnwBXP7lOPU1jWtDgc8Dr7yTgd4vidSlkeaicAv6Lfu24GbDW+hAJBqN5J2I+oqFvNu3vX7W
ucLFDJn3BV6bmbKCqyeAqpmS8DsF880sqAm1g07NcMtmxxlhyYhLtzCMIpSdKv4ZGuXxfrEVGmfb
wMtiY8dHNaaGbydxKN58dq39T3E7L3JgNDz2ob4aUTltOsb0tDNXBnv2XkAnV85jswLSF3WsfwWW
QNFC85kU50wz/3siWOL/sWaIHHE2FHHfH6XM7gmLdy0inQQ2ZFkXSYodxgmXObizU83GNvDrFYiB
T1IlOxPIIGxTgABbdlu0yESl8YD8mQGfkC7UH6Nby8apbVzEGRNGmLHSGCIxJewUre+CQbhR/jXz
OItnk0J4HE12PWIg+G+0VRF4nWn+/Gi5iU2AEcd52rfOS+ODzS2LkLftPHqlZp8pDfhZRSX+XrwY
UTWgcQkOniCc/XBM0Nt+jUPYsKgJFlHGL00sriyu98cdm8zfD4OJrcSZpahaKdhsHacomLr2DyHD
XxS7TnP1Z2PPnQSQHDdjs8SImf9oof2C4MUZdgOAv3f25R0YgPZaNechJMcemjuX7U6I1UnGgaBp
LubYNC+RJKSI9cirG3IZqIJOsJpx5u2y7nwKcRuA0YEtWqJDZZkIfAWmL9Bfs1jHZK7XmN90GLZi
BQ8cfQxWafsf9Uw7vDviRWG2ZUapsKDwFGT0BgsRsc/OPQQU6JEZyRqdOk2puMBXmn0zozfWx+l9
HQJr9kdm9J24pnwW4HbhxUei+LrG3PFIKm7nKqh+fIGI3E548QslV7Xb8GaaMeJyHwAJmBke/25v
LtVHS5HYAP3WGmRB6JkASgE6yPFvXLwd70/70i8yvIZskp+aO0DxfcN4ufS9xuzl9zncqHO+D43P
wzU7kwshXtmjlAJTKlaL/d+2WlNxUmS7g+jGLX8KIna3XiYjAgk20UD7zzuSKYygyovVD0OKQBGM
WOxz8RJr0rnLXJEMTZhaODV8lABstQZaBHMeOojdC7neA1NOZtRqpSPHKJW39ZwqCIQ1DMYybmaY
FA7jKPHsNlZPvz1Fv8L99+ihwHgPkLF2UzKOnJ7sqdbCoKd0dFr8sADNxHwTtV6s0TkdWjJJQVeD
1MAyWJnPm9GW1oYfTph9LxWe26NDLSH/aC6oAHGzXUn1qFOIDumK7KDJATjmK5mM0iHhQ+7bHoRc
yr++mf+7NT5kTSF7Q+r+QbYBJo+cNmO+Y6ok2fE8uxrUR6ZMPam3M+Q/2pQmXEhbVnqWbnEVJhsp
1+YIJaBdvkv6c7rP1TvEP5iNcjU7iM5XRSG2n9aJPH6VfjRG/5VuAxtN4LUNMd3MlORs4kkoDfcl
whJi6aPYr+bsokJt83STEXTY20PGDfxkY1QUrIWGqvQOULgv4yhggKBoXyR5VA1uAfP0y2LzgFuA
z05v77oLE6MIBgGNbKNDP1ZzUKkz+UA2nXMwLvkepbtUHqsLNolnt7CGc24yrL8WCRRwGk4JcCDm
fp0X4KqmKwv5iFHpPXQNl3oW4X3dmiYWhmHe7eGdw39R15D0RgP5Oy8vBEuW3opgDNw5Zx6MQoB8
qUymit1likGadKoaBZMQgyqrVrW0SYuxFyDvKMdhuLrENwLvXKkxSmYfHXMtpGXchbJYjrwrFtpN
sEtzSCpTAV4Xy5h4QMJNbF7vc3GwBeyJ/qjx7u9TTRbuSWM7Dewd5NwRNxAcLat7s6FgG0xQlaxK
Iy/JWxu8di/AuIlkdzxk8LlE6UD8av1ljS7JZCdT/N7MFlzk9LlhUyXJaQgTrb9Tk3VPflGphjZD
ljkTz6W5QNuZdgY1ZkmhGpPEEfRAZ0Gdd0ptmowTbKud7oHZRFD3HLBjbtBn3uBzdb4LgJmZspLZ
+wnkmDxbTrCis5rAFL1gqLWvNOuiEJ/LgGBakALlo28X8gCnCn13WAggWNDOevYF1GwiDxK7TdyF
g+xfwqOUULPSARCkAYIG227K3ZBXE2FP/4A5jM4A+4Q+clCawXk1dc1vY+SlO2/N1hboHVQ5JYib
ruKl78luI017WG5Rl1Qu5SpbgfsSq3bH80vw/G2gKhPY+/bBHDW4v6eqNuxXQBN8S1738mAxXBjD
Qjn04tStk75yfxo7veVDTDw7BtY5fkuFlX44pr045zYI8Z2ypbt7URiVgXR5NbXfk0bcSHz3SnO4
CfLWJkH48IHXHZ2IAARH9c47/mXqM93uyk0xPQemSoGKzDvmvrbJqN3XiiNR3td5LmM1rlRJr4Ff
YxUpXq8rItL7o9w5eA0DFMOgtdOGtrHwi93bMPaVnY4tJIvnngUG8wbKzXJHeTtT5lXcqB2Ma++U
aSqdt5wCqk8lg9zI0emjyNh6+hnuF26pVADlZ27pcQQ00bfhYYkPOZf+BLbPl+8gGKSGd0yy1wdT
H5dqtXENIBIOkSKgSC5Ep7XF/tQck9+Gp3dFNxNUZl4lpk5gC+D5nWmv1K4xNF6T4KH0LMuL/b4A
IGZ1eJ3hnW4Uw2XrcsCsL5SZzpscSfil6bvzi1m37zmHxjjXOn4u+I8mJ/ceeZH9a8dRIcq7nIbG
K8jl+WzW12Z5STnuscC5OmB4BDn+dySjH32VNvCgxI/kA6VQ634gBxDYY4ka/AHDFJgIhciz1rRp
l6uz4AOZgDf31088YDr2VsVdIqxUONYMP4pNNztt15pCwfXtmIfkfnpJ7zzbG7zkzf7EKIh7FWwr
mukUCg+KK27PqcEpKb+6eLiHk10gHPnDFBYzQ/JtA/BDqkdD7/WfSGp2gZrZsPJcckZ/HSHj5pZb
pK+WdmWwHPUtIC7VZIIGuQ/co0xwuW/gmrxUiKmNzuymGoJE7eUBS8s9h1PDVvvl/3lUyDgNou/k
ewnzwxfpPMTVB5BNyfdKsm2S0QOAAXF6ykd+CFr0MipUnIHkmj8NcR3+eZx+8KXn1IKJDYEWNGc/
2Pj64lJpfm+kBYV4Dfyjs3DqjQTTIqIuWBlC3KDlYWP5I8lv/sZfkrxpaMa1g3dG50jOUGqMC+mq
GAIB9IOwqDf+DA3jQvCLyoovfzjmAd/nSJt5tDPbQY8khD8FNKd1vXbngOKqaANJ4g77KNVj6nWU
u2gDcTfGX05IkmbsF8sDxYQCWbWEJt84eVQKdGd+Y3EaJLMA71FRKKYNpxpTPW+KwDKkwx1cKpaZ
yb3AtipJqXQFhVFLMZ8+E4x4b0TmTlQgPfMh7LJH62vfWEj6TNlcoqT+M9HqgP9GdG44cJiEAjRx
xTdVHlb2WnN2UohKXFWK9SGiiBDHPvZLW4qmHMtJv6Z+VT9A+8syrR20neGqQGPrS03Pq/w/V9kv
xWlByEDBAZQU42ndgKRwmvZBdTFAT9Q5seQ0khadN6/5eGOb0yrrBvv6XuEZxjjzwmg76P/D7HAT
mu5Zb79jEjwdCLtyGh4CfGUlndBnurxOsHsKFOxsd/3pj5zDyuCxrcWhVas38hrkfHLq9/st33/F
ls/xC7fXbq1hTeDQ/ZN6ehx/eKdbGcvy7FoFkYzwVY6UigP2BxxpdgoyiiP9lq5Xba45s0joOOja
x9UAYfMn1HeoA4H94PjQIaV4Uu4OYSk+N0W5nGE5tcrO0kl2Hbg2ZMDbU4eFG843CRAcWC9BhrxL
/HmZO6nSyoGLZ4qAXIr22Ijv07ZyNPiCrvMchajXzaUUSyEqgv5c3uHywLWl4FJbammmoZwx5YJ2
3KXoq37sXl5vGi/n4FBqT/X6hPpV1Ywhk4TZjxzz1Sn4WnFo/fhlOwLpy0P0knoj5HGr0LEyyS5s
GDPcsqK2x+euC/UOqgGc9vB++zdm0vK+xF3bWRuqzE/cUNgcedkyu60tlaOdqVALn/I3jK+m5ZaG
5Hl9CzSsZR0MR3mj88FO/6LzKttdqS2ZwfEFQo7MhKLvY8+Doov0gezsDfjIIu80bJLYbXw8FRvI
0QfHGdrmv9tbyFWwH/VIM+VQSdlwKU/8+5QRlvhGkARVrgaxihJe2dwakXifnGCQwJg+tYJaxYi9
vCW35ONLHkL9yR7VTrFbdlf4tG44J8nN09gJnSco22UCf+itqyWS2ytMOT1x9pox2aUnSESD5QIo
+iw3SeeRiVhRivLYAAg1c7o5KwDGifXxIaDnIpgAeVRiD7SaYOjxBI2Q1myAEyQgXk6rRqIBHK+8
hqKGwZWh4LYbGTJjuo9E8pwsmBjYgTJNMopFW068mkPUDqJy7EMsVDjTFPt7P1K3A67ItpTCvjzs
huwX6qq61w1hGEyXMfWY0e5GDDnJ8ZxDGBZ7cqQkmW6sVgLPXdcU2M5W1Tk+7vw8xJKfo8pftIRR
62WJgGF8B/m7PmZIJMVmxvBebs76rLZQ1V4t0PebXvYabD+7quTPiej99itacNTvjJ33QcG1XEzX
9Hyh9pZ/5LHMrAeifsJ7gM3nzuxMHPdiGXBBpdXGbdiuGkuldNBteGA+i3UWyELG9HyX8D/bmCW6
hbQmRY0PX50IPPtIOC8/sSE2cb7iGuhThdMLex0RuqX62LsAJmw7IQrjFvRUP1bxDeCi49weinlE
KZXxbgm9kWNSnQvF+59IZj61QWhu2WXjyAj0eJh32j3777ToHaqIMPN4Zf2N7ctXg5BsTaYZfMrw
ybmKDNf5DKeBFIm3GKSgRczHw+IUn1r083aEqomCXCWX1DVU0SYdn06N3t2H6+nx2jEmo3JowrC0
rF/3K6a4zPxgBMLOqw95oiOiF5AF9f7mmHsuCBuk3tzTJd1FI9lJhzf4H5s6dZS4lFcWW5DYilwd
3Af7dS26M7dhYuZ9rXp4iFaVWr5xJgQ666eS8Ekp5QZSeYQa0vgGYqFA7M+6tzk6HH45VxNvXJGy
uqzshNK2rjKgtftL9QW+VYUO+7rXvkPjjU3Sg+a4DBM4G76TXuj7QeIwwpnSlyGBLb80vc49l6nr
kpBrgi/Ln0GoAfZL+cDL7KXmn8CJmjQcWz1/ZVj0amhhFklpDkq2izPOR0xqd3gS31AKj8N3yPXa
EKe0pCIHT3pGXBfqHwklQAkoyuXGOs4amVnTk0u1EUyuN9S/ZngaFCwp0ycwdeIZ2dseb4lnKfEt
Ajsc2RuW/o3eQYIrtRkXVyaTuDARz5I1x324NTiBWtLtUoGc/1RPwWRqjDgIjKJ4gLvgvUpdeZlr
DH3SmmyHH4Lyz6h1SpfRPoVvafFAlUa3i23YF63lEshmUEVBDLn7ZBb8RqwniHXdBoerIyJ21Mhm
Rtd29CKXzbsZJVCx6zeyuJWIESAsEbKdVkWdu2rUqp9zcwp4XliOzvU7dAlLj4m7wKpy5K94MzCS
/2wdrG+5Krv+GvwS+3ue5SVbiZzy9BXXQREIFOaTSJ638Zm911tjL2rGwtRAA1Dk8bQxozfiQb2c
DjH1vMAWzci3T3ofoF2Umkf1j5N9qKwS4HEfq0Q5aXuXAqe3kDZZisGTbCWvN6XcIMWnJzdxD124
kGIG0n4aCIVidhM/hTn6ck/9D1uGIb9trWkFyq+bxUH+cHXoYrl/aziWWMZRauWYZ/YDmBbmGXHl
ZTqmR77e2QeyBzgEL4o8a9IuIP3Y2Q1d1a6U86mFjIxZ6vL52z1hedr7MnJj8bHo/vrBODGwMgIz
icJTAJN1m0HO3QAfqjYC+AKWzmXRSz3dx2qhRFQ75VeR8yHkgQbL2egvAp3uPE8wqktMtbyo1vL9
PTMImV5X0G/hDUoMFzBi9eQSI6tbNnvHTYXZOtmV4vd8dM+W+wxmWAbNZKJk/HYKoHm50zrGTdXX
PhLF2iU/HtDQ02Tc4Z/aN3zctzZP/cjthKgH5n3esY1+0TC0uckKhRlCOq3ad6wvp0kUIEeNE1CH
ji58nJ/aVYbna2m5J9NknPR/5bdQFtLbEP9v8tWGUY1fFnNqAg/QBrtaXK+b8E8YEH41pPuIRNHz
iypGV7sgTMVngCTWCrk0qkCrHI3+RBXVcJBgJlszUJZJOlyuWZyoWrLeYLQNfEtBJ8t4vcGq8VBI
dGEX5nYd4JVBfuYCViChrrx+ckRxul//mr1ibC+rPLRR6PGQiKBc5r8MwENkzhnci5f7+Iyi/FRe
nAFGqG4gat0Hg6sMKHUKxrzD+MGfEhXoasim21YwhMQejD1tb5Uix+HiTzaHzxZGUUfZTI3I1OV7
FGx2OFsmG5UDO11Ki5Q0Qh8pDUBwGBDIijCWCp5Ch7ZR0dQOqTPUL7t/upXm2FvPTAZqIiCI61Bx
+/OKO58ds2C/b25AMglgfnsHcjno7KuRBFI402/LySX2TIwLC7jKdEaUnWW/8uY7fx5/wVGkbmRL
5nUMMTzHbOlHba/MeRBypLHv//jiuSEhiCT6JuSelaxxZJ82nZYDXiaDoTP1pMxcQxuue8wCh0sq
VzWWN90kGpuHqluIOOMKJBlJQr2FmuMTT5Aij+s4w3JajgMu0iMZ7XtsVK1sUdmGkvSX8l0fMuHm
ZNQR5m8tK4JZSp1V/cB5aWe5ynGgtBem8badZnLvyX/p9DSglprzqEtIKjipG7R5GIfazRv9AKRu
bVJlPq+DsV1BkCFSoA3LvrGGkN2o5AcDGNZffR4fe10iIAtLYF2u9pvJndVJvZu4kDvy0Z1Q+Or0
2X2odX3st15w4+H6x05MJ3eSVmG1/vfhtfkY2k6AHXp41Zyif+p/NpeAmUogcSPKN1p3JdGdvoGL
3yhNHV5Sds0dD2/oY6EXgvSyDML1JMTvhumBj9Daef4lEeE1ofk39tUI0238YexuXM+0G12oSBNm
+zuh8aUKUVvEYqnf89GOqfkHD/ot7LNeVyZ66FL/EYZCxI83bFrMgxt+q2dhnKHk5Zmc9im47ddG
/28fW+L7aNarUgQ30KJ5Okl2EjQqaICVqrzy3OmfQO/8+w2PWs/8n84we8C6ZWWZRbwa1RLvXp2J
jqMXK+7/DN0k17T7cnw+tEhbWWvqiGnGOw8YDflDHsBE4ZI3PIypX8XaIlmK2tlk0V+x24H37X7p
pyhuFkOX/RczgtX4c5LjAK903meZwqCs0a+8BANYiqEzwUYBC4frzr/V8fUSVJVNqfIi/O2IGxP1
I+X2jDJ+UqjR6SEUlL/gSvJZMP6EVPMmZ+zLUmvz1g2yEjpVtvI8LqG/SBxZV/vgE00+BIOBxXuZ
wCZyn2S3ceFdH+I32eaepcxiEk+MTsAIK/Sr+BeIFV0YDWb4ndmoavJrM154GYJXdmzJG3jszZua
v2K3zrv9jp5ePeb8fhsIPtFYH2OELL7HTA16ln5NQDh1Mxk20maiM2MnA+drxaGm3s0mMps0AHE8
Lums1samr8dbdZpkpLnclHbYtylTvqc/PD+HaRUuvKwvMBHymv0juEnJ0FT71oki4CO/zTIsGXd2
MuKvMksHrAW9yb54y1iA5TB8BiwodyQctOX45kjoKsXB85RfNyZrKqTjxmkyQaOW3ElLJJOqEPiK
YrJzRrMrxg0GivNPEv/gUG6tNELi8f80qIhMBDdrgaQvD6N4R9xiGWy7fOBnUUXKzpcWB4kPhbMa
KrGiATu+TK4THT0G1SFt1MXFP3ycV5ehey/x0sjTVbw0fyhvh+wL9i0b6hhG8X6lyvQVeKo1a3ah
imt3gRO2CambaNPbox0oM27IZwXxdh4Sus1Gs48jm1UK6N5bEpI9GL++QJw+u+7LavORfr5ZyP30
BO1PW/1F+rBBx4sbOpy3kGiPY1brNSlm19fUdJVtxuRJdS9+Tuba9PbOyZZbH+C2HL1I741E+1kK
J7wWn+keAS9ZraI9RhlUXncPwXHtPSoGTDkUH/ZQzm2Wbp6RrQa/mb9ImwrskOXvzDMgJOC+DIDw
dTiimtRwBkzpIKGbNQU3y2tfhb9tWncU23WRoEnVjV8LbHUYjxUCxryyJ77DjQHJOMuIIlAL5ABm
wrUySgdc6iFoSCLn81JZQVyACHgFyYJ5K+6z+6Pud8mLzooJaV08+H6WKgUQW3tiQN2vMEJGZL7r
SbW8Xubsi3itjM9nVoMv5/0vnglluTykJDn29LBIewamuNXWntqcEUXf3CkOX0N4Kho/nQYFuxee
OA7DEzqiHabsmpBliEZvlngmaCN4/nSi/cuEWdVUsSrI0eGtq+7BxbUWwd1DK4N2rHZP0sZdgZQ3
5G7LVjRSh/fyO1p+3Btqq+FFt9cK71QL3QuGeo8DZTbgbE1GOS41yJvcYzdGFBM78pteswQC6LAy
0GZ1A6/goSdvkkWQyLkS5gHJY1SVqgWCcUr45BhCK5GB3r2AfBktawqdy/K2LwDP+I7YBqABm9Nq
hfQX4h+a5+DQPkknp0wPvvabuE39nFpssABNPfzrWHSboW8PS7xkfQhjd15STWc1J8eutLykCvtu
T/oxIJ1RHshSmQTWxcj3LiOn8NElckDTksGWrCVKDKggA+zbUuyCIjqEXyOiYO6lJDsQJktYoajX
n3wlfs4wa2NClalQ3qD71AA/ZLDWGB87G+H7FpAxJ7TjKURTAPzrkOweELdz/gSHgYiUuZSHoKT3
MlaSIdd2Rez8FIyprZ610WkoHizJuIVzsiVuMO7K57DnhnnAm/JO9HVKg1ZH5DenJgsuM3niTGG+
wxZVIT87nGr6xubg5TKzxnDVXZdZqqo9SVXp3lEvjEfH+luLaLFJfiEwkZq9113V06WZkDxelTb7
PSDNWt5yeLS7aG/v95ChBxNMQ5Vzl5+i01eshcOXLghWVbgdqbFocJ23sQT7Tk/0JDQrc8sXeisn
GMOB2Xe/k6FgkdLvelcFQ4I7vrVKA25EDYBw7WTdpqJpEdmt0kQCu85XhN4yuodFYfBirXMkjE5C
IQbGvnWivSZaO9svZaOIMyT4fBv6DH2Gdqm4KAMmM9AeChcPiIYq/5VE3NditjocoMcj6+o/C4g8
GZrmVXZAURqiGT6RW52ThJT/OxMq9+Xo0gzXhR5kT86s4Uffje6P0XwRAxZ+GbfmrW45p6QH5SD6
h/c00lGqYGXkpLOe36cp5j/cdYofBXF/5K1zwENzKHRaiO0+7xD8U96cM/e7DznxfURTEZJGHl5Z
KWZqEh89wMbAnXtTUenDgyhOhYAqhFumdBUgeTXrbcMH2wVg/nQoLPfJ9gljwvdYQGdAp8swSHaV
k9BFRR0H6997OP9DHduNXGRoeqj/YIKp4zjRcUNQuHoRaCjXBc25sQAtNmv9eRYFO0fb0bb0KtWg
biUxR3hZfXgsWHb2BN4JMar7CAaE6EYEl5x1UEWnc26OVCB24jKeZhtorJgLtE4ZhOFwkOvgC6v/
7ZOfxe80mAVab0xFyV9YCOOBAG64/dWz+IDhl8SQl3dln3BzFgdVxrpeS7PTi48J1maHcnvJ/Jf4
VZ0MTmdaelndmc2VcbgCOPM5oDivm23WHmGtuVDV/C96DCcLGZY9LPPUmDdvQA6gEb2iYxLBeCyO
hI9f4g838HbZCQYi+wyMfsB2aLMI/igUd2SGt1y16D0MTrBS1z2deahutCCDJzk7k/upKBXhvMLJ
PWM0s78XHjDI9mlEPtDNH2WV9FE8d45E5UVzmpcLMPUY9XE5UmikmshcvU/LNRrdZc0wa3VdtqUP
gaZZRUDnQQv93zDybYvzMK6+QO6LepN7jbHZV6+HVjAbvOknn+w6vKgX/fpFInDyUvNpcrXVf68O
2h/PYaTQ+G/5d26oDKGSCp1xdBISG7al/zAeetqu+485t4fHGxSzkYFY42r/kh0R802JsL0ud5kM
KKge20Hs0xaU7nWUoYrqC72Fe1to/QCzn4c4rcMyvzxC2Xg5CJ+DheopndPgv7dNxdZjIuIiRhcZ
UtklxK7qak/yOGuhwvSfwlQCfB4LvOixAiAC0S+Zcx2NQCrzje6P+X6UWQpNh7EiGMz12fTi8wxp
gZsaI5//EvA7kTN4GYTPK5BT6xyotigbaf7ZLIzcu5KEhyK3cGBT6UHNWg2PohfkTprr5wwdDrik
gSX2OxcLISCTqFoEUGDa9mzud+am9XrtG29QTVhhrDuxGitRtOM4lNY3dM19yS9MRmyuyyxqyYBk
DmOlzBU4+Wu1yqowkLECfWycVRAwRSUIp5hDcgBDuf/l9Gqrx4aAs8FFMTaqNznRKjRvwm/pO5/R
H4Q1qJHgWykicE/pcBoldZsBpnWgh+5aLpYQ2lzDpqwNuFBxYo8FG4VDj31TK7k/zZ0+WLmxXsnA
/Hy05+gJW9Fg6P0yjVnk8v1oL7Wk1FS16LKGad3XaZ2cVpoESOxVf1bZm8rFyP7ExzarlY4TIJcd
lUl5Nfblpx3E73gXe6JFxSYMfUlYpDhdtv9qh2CfAB0/cndhU6HV1gzDVh/lzS/rAjpYFojnk1cY
zt3I1itGJQuyYELhE/12EVNHMkMKbi4FkJW2HRw7lh/TtRrQutBciLY0WYnL+MzpzN6M4TV9sim4
PqAxX0twMD5frtgZhXgR4GqtmZIS4pic/I/dpzqTu19X8SLRF6FZFRJbZTmviU3REmu+BPC+Zmwv
MrdRgr87R/MvzVOWTnfqxkiyJoXftvN+V161SUhUGnXBmsb/59PNZWf5fqVwFTR8U0AWfapkWHQJ
dJms9u2vpkFrps2p9hNEjQOKL1BbEX2aW/p+1DqQMd7aqLhCMOeTNoMrpruVPd4hgyJmiyrQkgca
HxoVwDL7cM1yNNmsZb90Es+d2nkSVwK68D3kjLQ67JJFYsdVYO1DuEV/FY3ClqT30NMvPXSeyxPI
255lD0XW4S1CBZlm+U0t0/nPiTn2Jax6uiumK+uC4u2ml/cR/FbnT+3A5H0SYhILia3Uq7qRpbCc
vlLzx3DGP5wu6rraUNogRc4nRJb7YOFYd0ZFdPgViOGxPOfLfqGol2CGlL76GJq6WbMPnxWyMBrL
OwiA//etxx415+oqsfC5ninCRcAvSgSIUZ+NjZOf35RtZH9B8dVdNTXuidkmh0ehmpsQNbpITE7j
LNlAH7pCxOMEay5R/qH+sAE9eqt0h/jgomLI4klQL7tK5UL7xgKZ2f5IMHPbxXn3mPa+eEWZOXNQ
cG1BnF6bpYSVlb6TtBbwPACjQkWOvKGzuIs4/mK+4axyFRPo8/giAR29EFIdSFFwGE+qGva3Y3IG
3HFhSnKFCV8nyvKbCK0hLzEjiHsbvOy+gOoceNDwKjQLX+LIHPu5Gy8705bp8CWQFxVYEICG1gky
nkfACMD0x/EX2TNqJMmbp8FmhATStkYw33QbnbFCGRaxSX2M2SEwTVO6muDbs5JTJeHqwzRoW3UQ
b0maWz2nXk6/AyvHNc5HLdFOLHT6FnM7j5KsJLzOD73sGGYp2F9At73XzSWHqGW7lby8abYpiAXE
g2W0CVy6spsX26ULjprIEhIYquPTtM+Y7iPplehiRlK5Xvb/GDwhNZsnBs0Rud1BOuBsJQNni/4R
0vjBhOK5sR8Vl/uJHB4UOJbgEQ3hjzot7Zw8xJ6D52MbKveNh+DFCpF5gzlqKsmeniA+xx8Dpf4p
Vfroul4k7V9fQvGARtNclop0SiquzEWizKTfuEf/1UHcBbY3/YvJsfQ9xZi8RLsLK73qpps4BWpP
8ZywooC7uNZxZMx0Ca1MNStQVCF9WkM2EuR9jNyJvP4DS2enH2Ft4A18iSY9Q3NEJzg08Aayl1Ho
R+za22hQLMlcfDO0YxOrC7W2ZLs9MojX4Hd5g8Y2J0QKv/S52OusuEa3UIlQrdbBO+30ZHs8BUXr
NZ2Ap1aw4crq1WeG8WXGtDph1K3icJnnvjcr3supDIYIGKP01Try3d63CkfjtJg72XX3LnyAiDu1
ddQA0B+NxSm5eHtzYlMID6TzzcLrQZzJEs3GiFg7Ogea1PDFRtUYX0IBmaG2WF6jemEgbHMfFTcm
5CJ5B5BdVLL8+LdXKNNZDm/vAlvCdlZkj+3ZG0NPrmoig380MTrXa5TfmiYRnPeaIdPfCAydNwCp
3Wpx9XbV3McTpa+q6YGPErthdgmQHQLXLRqvyKS+++ngn3WvT6rV1PwZ3COkwDQtYdLPPmhTm/jw
J079UfimgE5nTNkTAQN32jnqcvJaE+5LGd1n57UFrvYhT3WOg4MFguROB+6edJ/FmTfQGHuREvpe
lH4z0c1H6DGpH+m9GdmmF/FT9iLOPJ+RhiDdOLjtooVsYmWOUHNj8ddbDry/DRNXP7wMMImev14T
d1QvOtwdSR4UdSw2Qrs3le7tfFwlbtTyJ0+zPNG6CIakFaZSrBtSc0k3HrgXRixW8OEYtMqwANib
L3eY5rmyvn9QQQJMy5kIiuSYX+mr6jY7ekgLhroND26GzRRVmWM4Mu8/ePwNN1YD/0kBNWjBzM1s
eDlKqwkOkJ3Lklmk6bfny4pYrb1ru5PIySmMDLZpMhVQn/UGzUuSkQgJMC9T5rVWfk5j1Grdpfva
w2Lpd/Kz+dycMAnHu9dbHWQFl9LV3XzmprKfUIaltzIn/geglCnkPBE74KQp4K/OyqdLed5+6Wx2
zezi7Iiz3Nhx2C8NYyC9J/Jotk1EIh44qaaJzuzt6/z8VwaITTmioK0yC9FmuZfDoIcWfkGbPyTr
1WMSGcwbV0NDxCWwz2PF9DUy6ydbpPlEd9tB8ipSv+jw4qhDRvTd+P8tJkacfH6P8qio8ikSfR+E
64tpBlu5H/+74YW64K24WGzcLnc4iLTHC/nZ2DHZRxxF2UNw0ncvBPwjzZPgkWg/kUl5gCAnngQH
3wVHFs8RSOUS56C4HslmgKloth6rCcxCUkjkwLdEzBxy6h4MAB0XczHXCeUN5iqKbejhUESFo3T8
YieqE2jHqC9miRK97bXkQNtAaKaqpY592EWU4OXmEqVrexO6j1VcwKHcKYVDfg2aQTM/sjHwhMNu
XXRkX6JaGaFs42TMRBhAqi9F+OR+7Y1BU/zpJpNugwzL5fRUMEd/G94PQSFZ63jsEH9zsqBapTNC
b6lOErU7P6IZvPmrNBdsbb8Ad2ZhpXYbl++iDYxa9KJNEpNQhGFgln8Zlo0iaslvBFbtJGEHBpKa
h3vSx70Gf/MxgRNTHlgJaJq0on5g42knjSm713WxP584YtiDE5ZidGJKJ9VM66/uFrtoedpaaabZ
5vfZURmsiXJJ6roKJOAMoEoVWA/UGbEEvPLGAE5eEIVVZoXrZWJHyKiS9yYjpkcQRE8NePLEbj5I
ONfMnf4kbWOrSklChTLRbJXPfsifnFK3HI/oTj9hIOskwXVQoZaIkbWLdtt8a6yvH6pIdhE+Jn5Z
UkSgj5g/q5sRM3VjJiMQQRG+AzOmZWhvW036aPRmB1q+Q/dCfXGA02tbt/IZkMOOkYF6tgkMhVsk
1JLULKdo/HvXbcAE3YLCqjFQDdwxw+fsSUd8bA2uoFHV0vMRd02ECVk1yyu7hZ6D6V7BXI/j8Ut/
Ehm/vKfWAzNeliGHnzvJfPeLEQjFM1M93UKQ55rnyw80XM+nUJUKDfSs85N4DP3BGCOr9wc6bGWu
cK9q7T2v7FwN/p0A0/Ifj09WtkNSoX9ggHUTx3jOta8KXtYULbXzI0pYMX+plrUFdm2QoclICT1I
q6sxauoNjxadmug1sNPPas6/egO4Af+ax4uMk9XZ5ut0Ac6SbceIwUIj5c759nzNoY2xw3B+ej6m
D0+ngE1XzvMoM6nnLdDpe8HrsfuYIgmptMIcQBBow/rmyEqdivHkpPkQuLx9YKI1AFYWDw7wv9lN
GzhQ1csNOvnVofJtucbyWaA7DnPGozp8GaViJHyR6i3I+oGiLvO1BeIVXq5KojywrGNJMNco7fv+
ydTV+z13+Z8q/4SCt+52tn0aZBp0NIwlFhb2F8GM+5NvQ9ZagBUABsxcEcKZP25Gu5uWE4YEIBwv
FRksgzOB2KU4cCbrcgS9TyRx5R143cLA0FWLtb8O9CbjML5t0syZeUIIbRmCGSktq3Z+4Tj8n9kL
Q33ZPePoz1lf4eexXw4jwntdcWX1qOQhPjIdOvhdjv4KylqshAlaHi+LHv9UMD1drRsTfhaQuwxs
dweM8TqEPTk6fW1l0NiibUz/WuPZrahHgEy8Xlz5tdKzn4JUsaoCn9ARdR0ukXAHuo/xKoMlEdYb
jMw14ylbQSgGDofClfFHNMt5C7xy9/ikJgVjtER1hSAvoSwgOLrC3zBWB37egUJ2aFqQNtqsoK+k
piKb+xiAFcXK8PiiXo6ID4uHEoA7RyUcFXuZJOO+b3/xFIIPGOkvgdSHGXjpj6AQoZspzQAoo6FI
Cz/8iioqn+e4ZFX4TTOk/HA+RCMf81znV2fTQhojD5vZX4CletZYk9tJQHow2rG2fL5IQ43my6EA
tq+40O3g9ThvKXMoyd9RAYUx2EnpOMbmZrZKDiMRMjO79SM5vCGjCYUEVPHLcRxjHvnPuImSfjJk
EkABFX08CxAvpqcB1HPBrMIl3A8Sc0+wFQY5BeXmHSy1HpHfkJoLi8n17kwYuPVCguGbO2If+Wz8
sYYwKc7fETAt+C+LMaWrXoXiMGX1wzHYvwOABL+VbMRjq9u3QhKdU4FqRRcYQSIN0JzanI9k9Scn
sBHcdzOzPuntUXTouQVR5JZKUa8gUua/StBOC0oOW7aNv/LKM8sJzyTsuYDrpeTuSe05Oe3ItyQp
j2Qj4KRT00L13CgC0eW0YN15uH8fil8XCuVMeCD8rN/Ee+P8b9ltRtF1LEr6pl2qWp2OQxogdbjI
/q4hoYzhvzlvyN06Tshh4NwlvVxLdE96/JV34mws4v65WANGH6PCfAWh8tjJrWWZWVRR9NX+YsNz
vSEgr/1851+/Pi5MMvkkwcS5agiTYgOE/NY4+02pKy0wiFCGjBek82VE+gPdAYzhr4pd9qXPrjRk
GxIRuY1IEKqN8sJdVU1GghLcPLdD9Pyzi/K5FsTqy8DCt4sIDRynrn7eGZbZAs2UYvaMoIruv2xY
jlBK2DTMQj3sNLAPlulARhMQ7LjYSkYueJxDgdWimWQJ4GQdfjXH0PPV/R7wi+dBREreXWXev6AP
5v1NT0aFXNOAk5eOsiFNMA1rSdwD1zY7k7i0DZXdXl7ir90hNHYabHjphDjtsP7sGr92bgWgqKaj
adNbwDBkZ6o/4dCv90/EONo0sgPnCEJMG+D5MXjEgsI5GEkARnZ8V7zcSG4Fmab3CcvKspSnUv+c
Hsp2Y5YwJByvhjNK/xKAH8na4T2IuMuto+HXNeS13AvheD4CkunD42PaskKhg5F1jQnN/KIG2YHC
c88FsKkXyT9zdoI7t3OqHpgBB53bY0rUZ8it2mCsZGQpFdBw7LtnF02HTw2zeX7p9an1on2CQFZO
NHRs0ItYF/ghFTZO0Jy9SNPv95f1w42GohNPe7SSpPQj4KkXSNHpuIgGZO64Rz2uq2AHKcAoPOIs
rKr36Wb2GtIzSlf9NFE6WyBEtqMbygn2BB8c+MiHQYrmX297CWeRMfkTv/EwnszTXON+7grWplSf
Xy9rSn05UuolCn71tzjvMg7A6VGafJOBrsf9ThPXG9wDbc4CBa4q4WmtC9YgsJER49Xg/dWWNDVZ
jtQyj8nxBnGVuJBSd+i+kxj4r3Zwi/3y91Kk+S1qKBY+zRp7mGXZIEnrULnkifRz+8DPUaIwNtrO
mMikRqvGBIPVkImRaqGpTzFck08TrUlQ3STrDRthlsHyzF1E7gMsC19N7FFGYHBDXh/utNUOk7R3
AJT9ZUYjsGLF0xy1bNP3GswVJqbZfFSuzPSuWTdLQXqCXLZ/YWGrcqZRiUORCmOQbcDMtIhGEURd
1IemT2uX2pbZRAQl/DdgipAWyTdGdVhA0IL5FRi75Quva2PdbkRvHIYReXf7l98kOf9XwS+t8IHA
OfL7FlzMTZ8RNlQBFrZXlj46Pxl5RhmTaTkKGTVqwTbKrpCCT+4NQFsgvUL3UXv3K7DgxW1prwMP
NQjMMM2zCnsiv1h1OJxtu9o9EKo7SnLmrSOXi26M1RFQ67nIA2aEd/OXLyimjrXCitAYGGyJ/ALb
U/3JmCsq8v2lJhJgg5JOAT1fiJGJTUoQMirPGDeV+3OcZLfFN5nDok2/HGCDMK1db3RLorSLoGuq
+q+HTxy/riI1d++j7BPfWNP03JXvXDK9VzBbGTGoQNzvMNEWEr3RirufxU4Ff96G3cZEjeNzcbhN
0ITplZoTECLvxDXaNrpp/KWvEOmt2qpVZlSFcmnU517u1yrZevkju3nXneBONWomYFOUIROUVf6/
iCp51uojWLHxeswHADw7D3gFLke8w3BAJg+wQMsqBKLzjKJGemBghdLN15Pqq6HBr0zu5hure0IG
Mp+YljmkvDgHhPDgRc1vdLS5zO8ZLqYPcSzzwDKniiHEZ8HcOzi73gm9orAzyunaOs/lnLehv6Zf
nNqhGUx1JTOoGJvekzZpmuJ7cslhG+UShmU6kqsCGQboLZygZmVb/drSuwFM/3ezUHFJxNvPjyWD
F4EeSjL2stFypO5p6f8omi4+Gd7/ycAHxPHDllR/wEaMnAj7kbGQ88AbZoeuUmXHeerBgFXI0Lqq
g33UsNgLePzGRYQWTAPQDd6p5r1a2mLml0Kx2VjCf6/B8drySfmYeDNL6m6XK5YXKmMHgZw89yQq
rfcNbQmvHEA7fRfyAJ0OQTUNOMtYeY7Ij8+x6J+uJDZS9XMtQByaovM/WD7wSz91pb5tux/wIp0G
U0UvmhxDP7k45/39HH5Yy7NEIPz79vuNuh6iqOKuEkbJGUp8zpAo1rH56jkQjA+44G+aHuNcNssg
ZTvtafCjfHLoeUBI8QDACPGNvGxLCA0I6tAq8sCWlEr9T2OzlJ/jSo2/7mVlG6GaWdCQmcRR8Qc6
8LCtMwMlLnIhnjxFFKBEcWbcWf5EDmTm90npGBPAJRNNTcbhVPoIlbXcDKQHcJQJ961VhJ8GbO7v
HnfciztjcBAm09h4q3kop/bFWfmyODM1oFfLtIvjs8ueSYog8bYKLS2DP443bDHh0RSkJUUILdJq
se2wUtC7dfzQ0vkp7a7g6VVIHIfdlEhplG/IvpCAN87MdUrSR5MqY7mgxMBG4ejR0CSp21echwrz
hCgdmUSO8BlB8Lt19D1ipw8h3qNKXBEficVOweKOta8IlHPSxFz1P350IciJ/gCVLDNoeG9qv+Bk
oXpIN3n6mNJzdimljBb3rug11UWKGYPEw68rKtL0gDHvd4TMVB6+8daHCfbDbRVid6K0WDlo1lm3
pHQIyeX7SdUPqjkXkxUbKM4BK4VpascF1btr7ssTGHA4aKi9WagjaWfSxSMxL/qLhTqYyoI+TKak
tlkWYXCuBhuMSUPv3EWt5/dxKA2v+0dl+scttM8i7fqveeA52mNU7aX8u022kQUBXdpjHWioT2gD
wmDMreacXaDdszV0vGcSJAQFYh3f3fwbII7q4MKc+y9Mg21L/ScQBxzGadof0YM7cyawrh/63Hbk
sfMHoU4TjlZ9XS6hVR2HdPX4z0b/e3GI9k8bz5B7a4LajXLhA/2sEL88fOyNEolCeaM1rHcz8PQC
pyhMfwtV3KqYQMK9Q0BLbnvJOqgm/03EuPe2f279TKsSaXwMY7ueVeMgWategQcLPnhu0n5uN5On
Xcu9OKjkhld+SU15u3868vPtjVP+oUaiqR8pnk4spL1a6SyNgSk1F3AOc1QPlUy8uZyvr66I+gWG
GgUWzspUNk4BBb3pKfDKwwrscrPlz5RQ+05TbWeG7YkvAGvpgFYXORJenceBIPH0aY8xLqrqQmT4
LCdfTUD2nurgE2j83P9atODdTXLeDSokkY5W0fhoZMYm3mxJrPEaGYfusKM31bm9WwWqrCqDy3XE
wZIdpsGJcEV5OU5855u5Hql+D6s5vm8IijXJjSzcY0dzeqt9NL7a5qH6TED2kEL1/SqukAwxCyGX
th+KrHSSFMUYr6VBGPYM83g8s2OY1pQ/WCWDPRfaeFnAZKLmIItHQPmzwSXoaEyZOd/IpZt77DLF
9zZgh9AdVDcjP/gDD6sUwNynOSvFHM6cvoCEhG3wK7Tjrr8ihAXKcsXAySc/y54d4cqSB5hmXBfm
3DsDpi6tlKGGhwTJQtQIgqgCmGyD3cisxouiMbG91BJgU9FMMM6YVL8feInurBMMbTkd0AT4bL/2
6uFJKkPHn6haUeO7E1gZidD6xaKGwrTTI5ZKVaU94ji8nh+eXHPBUYhzR23KILNM92I06dWx0H7S
2oyIHPxhsRl+RexYuVnMWUT6pK/uKqiDO8iIeUzDQT4H1OnynhLfGf8UgwSBbxYlY1P+i2Sxyfyn
atDnqflVQ8zLWFlKgMAy1KSR9aVxNtdTmkbsK6N5YiVvFzdHYa6WsnftT8zdrMfHs72K2c03XULl
8s3THaZvJFOeaMyBxgfuZSywvDo6djaZILYSiMbKXc7pfIKfY/Buc3IdkI2ZF+WDDvQAya7amMdu
YPt0yPbaIaZv0OOfUZcG57woVyheJtG6JEeUYzViTEfYlyFE5K4NQxl/d39tpfAWm8rN7r+tabZT
FbpdGygzGpBHgd4jy6IjuUHO/FL45+ndQI3+epk6/rU6LsoHh506vO30UwMcrqYdYE2+tglbl+Cd
fBJVmOOrP2oEwIUDv1r0sfX/BccyGQgX6xL+F0iHvGeVnGCCLu5J885NfbH35XOuYE48p8LhiwWt
PzvmLSBvV9CSIFFpRyKkSW8r+MMaOnzT2bafnhkaWlaAe1ET+2+02kHWGHQWPP59Pv+j4hoZcYg2
+44FUnGEpfWInCrDvYLrRTVendZUU8vtrhxjPqWaFJUutS8GDHOkQCZs7TvxLTThIDIw70U880DU
MOFOzF322/uNZtjjGWFZOgXIF9N9buJyAamRh8vA4snt9ku0a3j/7QYGEY3i7402qCn0NbyZnnio
9mnUVU7GEFfFXPd58VZ+XY0aTod/BylPzt6qrmLadRfmU2wlaLQwQZ+LcJLyG7dYYh3MBcjIOwys
RhqNm398PelNa4dp8UuoSAUW3F0vZ9OWnuJ68chmZMDTTn0IvO0Xk81Hm2AUK2k7ZCQg/iQGRrXK
ETs9fKHHqChQnJ8NYankT8Fok8gy3jA4xyHCbMSl3xXuw4c5lpp13eJNLC9jWPn3eQtUms7rDOmP
cj2L+ukC/txMXiX2loLMcJ/4p1ezctGEQcz8+6Vk3daHGtJUQ3BJFQ2/T49IBOw4LyvCsIqstCPO
zFi+a4ppvR0VLekdOozFNNOHfEwfGY2NMARkf7YHoG9dqWgjbAixNdJbuKnmCBIplbmT9AdNkhfU
CWTfgsdzh1x30hDQRANPSmUpjoNWFM6YiSmc1gR/zUi3YO/Ox42B59kySPxol29R7DlUTtMDUTjL
uKdVree1GYuoCCkT9zut5uvVXVwiQ8qCeq14XTahst8LUnsy26HcRyPPwKfh6PVQqdqkJDuYOqQa
2Nq7npCq74UJ2dJijxTC8CG7M80C8VMIJoo0K8Rl4s1geOSvu+8nFvsAlCqaM8pkp3xp8GNvt6BL
3UHyDCvGOJ+V8MzKOs0FbTIbDjFfNTuM0QQ7lJt+khXuGFkCJVnVKxT4sv7ZO9PkzKjLVBlkha64
dM2BWIK7qje7VBztrsx7+ADz6Na22hbEUm++EzQafUd4AcdfnIZpP9PnK4ezO4q1GpyoqjLOVehR
HSBS63JLrX4PvlYc+17j8PnQRlNVsk6aSFLQPoPmvRewMOjR7pgvAyuGNRjiy2F7zJvgR12qgYpL
wPN2SZinZs+Vr7GibHDOhobyih37ololgUG8mo+686kr3sgcAEmg+vvo89WBMse8gB3PAt2rIG/r
xVmoto9MunE9d/2LY8dNcPIC/yzaCimDAWsrkn+3WfDqFKF0pR87dPa+UyhZYkRF4HWZo6yVENVW
iT95Q7P5C0IBlc9hNoLwNUZ8uxHHy2FSKnduX0iyOJfXJMfv82oJ4hGBJjiCHUBkpiCYbi63VkQp
IIwwzfVXCjmv5JWIbQ6nQGvmAZEOYcffwnpi7+dUQ8YjCv/GS1RBoXPlhj7wZ3Dyw21CmvYENHNd
bbHoJrZA8Yj+MmFW9lNxGcs9BM/RR2t98Tosiw/rNhvZQzfpH1GF6Qbv7TAQpjDVx0SrIRLhNjef
sz/VugM7K3n12EhEE8qO9Ghmmpx0xkrYzgNqSwRfQsANTOGJ/2licWvTfki2e4CDZgfOucyvQJ64
yA4spMI8C4GFm3Oi5d+m2KM+Ljoeo5Hk63DSB0oLSWMKjFbPDpAKucbq3Ot3f6OQPFSqOX9r8tZz
Jbn6beXsN3Yq0EIZLSn1fO13vd8FbA6Jkz0EsmgKWsRhy2Qb/UuBNoiyGk46Wwl4T1kfMj0S2Q0t
Tsym4wWNsVUWY4SOA8imlaCN7GTJ6ybpeAkILNZZas1DyWxS1LSibg3OflfxTAFewC2nMliRvsc9
fk1b/Wb9O7DYPbTGErUe9Y2wOnZUseXOzTyNKCFByihtQfRij5bc7mRrmNTSXctPdipNR2CnquNT
a2V+DoxbChtzerjkZvbsVArkr2iOPwJS3q+RZWuk4SSQtTz/bxnb5uItOzY8HyaFfKZX/rueiE1A
Njn8RdFJaIh5mzk4W6v8SDgdPSyVvM3T8yuAKjYVqAuJwT5OjtbXBeJanLM6B5kihbiCYm0znB50
qrTnkJ6BRRk4QnqyYyRCLhPsJ9rSlSB+JyiTrlL903/4KwT56p/KH7A9CzS6B3bJwWlx0eIs6qJq
RJ/udU/4WmFtqUrAH9q5W09Han/s8M5bn+Yl1Nc0lGuEJhOrJOdcpWa/RhC1YIZWIpYP/huMtFQt
ghF6kYU1Q6/RP+PdElL+HbWtCUYZ8zpO7VoSeAhINwpjEf/qei/SsKD/TdjljCHcbfTRCKLusEfB
n324wlW5psPR+wcajiJTBnNZFZogaMoSkdfO2WrrVqOzvaHLRm16Y/heyL4PzP8yUnWFVyzVgdeu
2qNIjLZtJvq6//qRwmR2v4mwPIYmRYYgjb5Ij2uAWtzKmQvneurwT8Hq/NQiX1AJgyYhbpH85CSo
iDiYwg5gsaFhcCzTLaYBh/pZakGJVqEKgwQj0HA1bxp99r9QvVu8yWfIAeEOuzsfR8nJYzhEyZ0W
GsZRaP1PGUFdetZpgCoamXK7I4XTqEYFU/lCkGlDO6vMS/DRp5aIfqBLBVJaQAif/Z87k8jDsx2j
A/VwjFskmc4BMVNKExQutFekpWQihNrdCzCL6jHjBMpYIc3P9p+8OWHmFVPZOkH5MhMi+dn/4IrO
DhCIgMCsSsd7KcyI64BLGfvRepQ95m8gBF/6DSDtySRjgXvH6f1EhmMkQdzA09nUxFsxL76YAN4z
IAj8rFk3m6Ty8TDpFpjmTvmfMQYGeY3d3vBfbK3fklzAFrULJyH882LRj+XsVkJGA9nt8jO2UrEi
qYfDV1pfgjRacR1YI1Wp3LTIGD2c0da+Ql52p8OfyyMffTyugj3uQrDRcrAl7XMhG5v9juL/o1AN
dQ1CbpoKC4HM3/kEm+zUeX4rVAJIHq4O7JighvKqqB5VBZS2yv14wAKsQ/84B1wZ5Il1pHQm9xjD
VS7tgeXt/5/nMU/qzaBkXkW0A9kT6d5BK9UDWcxk1R9gkWz/oAIqsZ4XgBBsHoWNMbrtPSb3hkLM
A9d6tmhcdjGICYBcPLs+j/WJBk+YNa/g4OvXX5PQxcEogjNo8Zq+9zs75fqGhDZDQWQfk95Dmmeh
1ejCVfMH3HWifp2M0vM5w3hCeWPrCzOsBEOzGXwJ/mz8VI9qHaay3sJxT0bli1zQif5NKCTtS3eG
VMGqXz8bjnN4H8xzPdwe0u520dCqx7cLTsUt0dtFTfARzZU2uVRPGy+AkAXkTCY3eoShWB98KHTs
zDSAyVK3qzd1TH0fU86oTAHBL2YS7IzaMrHZw2ONp1WHgsfMtqt6OxR3/MLWxzIBV9nXHPtWguFF
xzIOyW8Ix0m5mA5eiF8mrmTGY4/vfP0t9xE8fmwldzwISiZXCLK1QgflZrGfkCJu83XYcZQ+eWK1
iUUt1+B6+1/TvICLWhRu8RyT+SndYc3wJ9he52r3P6S2G/eq61+y6SWuuuxJ5kbBQqEgiT/LZnBl
t/YNJCjHqhjzUKPRTOqEA+Dyu9NejnHkBGL9waY/qTk7cuNbrRc+ASgptmT0dKLFfD7zMz9/DSfe
Rb8jyfOhDR0004XXXRDn++WqbbBIvsbb3m9R/BkkSOMkXJTshZZ+uATsBTDeIKixkpO4IQPMWR83
BcK+3BbeaJKvF15FBQXA2wG+qZbrHaxoM9SGeM2zWRYuzESmXTXyz8+0WDtrLHvf2ecDNYF6GHPF
TrDJMVwEwWM7jVvJp102coznmw/reM2eVSqL4aCQ8qhr02nVGpBY1bnhLwidgesCTd/7rNkgBIYW
fbyE+ZaXVNhxqQywEG0wNw6YGAnrdgagb2xNy0WqsJsKG87jkMUGNNk2FoX0cgVPj6v4KDxXBu5o
k/gt02lwu/M9mPsxnj+4Me216qM1ApjNCjO7CmTO/s1svTE9B8GYiTC3u1cPPXldA6LkqxnwpKWn
KO/IkQ7E4jg99lXZx5Nv3/qnxfCV5cPKzE3xvWPfG1VNNczdqXZm1Jw5nB2nTlNkRYOhM7I8j8dd
/Awc7vMpbdxkLfxxK1st6E1cXqWNcxHPXHLz+oK9G17xgrm91NAwYobkcGY6XUo9htgWXGIa1w0q
6cjAUYKaS87SOlqGVi1K7Ks4yZtGj9AncasBawfgyrfiXWdf7yaUCASSTxzQzD3u94PB9o+nTPeZ
2jTH6kpQ5bM2L9VodVqH2idS7bwcD9EOl4UZsuFr9juqWiEDlm37q/4NmGANzYxhlTS0g79bVhjE
rcsPaZWwnIPyWSP/SccJmLJspf8H25oQ3cPldPUWhNm8mUYr1e3D8WTWRaPH4OXgnUk0uehJM4G6
UAP/qQcXEa8s2sC/YBa/pmUdcErUSXV1KFqwZn1ftMeFrCSV6VKT/Ln68FvqSKdtSXO6wYoqxGWD
ZBrjmI6m+IGe9JrV0KiwOEMl/h7qGJsqPSsunPBlKnkQneLRgmsHqNnexIA1jjZd2Hk14VutfIng
25V0PPrUmaN8tMEENFVMzjQkN3TGbHoEl3z3TwaMQHbvej9b0nzQSYUniqXw5S/Bopjejce6CDHv
48wuPQzM7zwmAaWSx5ezopGTBlFFqOsBulpQf8OlPTuoYcpkgsG+V72tFXNWnUp+F9MXe3/ygsjo
2FfuQzmqMvaZGBp0M1gYBQpw9pxT1dQHbDfR9sUjlRGA5s4+32Ta73+bOGyoBLAZUKIgfhbT9z7y
oclFcXtMJL2ipDO8fU7FXxynH8HuNb5KkRKcAEyJB9SNmpq8ApVDzfOgsBJEq51OPUou5J8Crcqt
uPgBoGLxGorzkE0ViN4IoNAZMzbKVXOQbMPILRWmHigfIajqXxzfAFgqPskslQ8lWWZ2FzVf6RIz
BhFqxT+PvxjelrQCcQraV/WVHfg8H7mT39mE6xqjirc6IMitr3FWmEp9ZQcC2QeQ/RgI9IX/eu7t
3eDyhnY4UlRS8NhwHUQn4QgIse3RMhz2ca75cPum/3cJflNPGwrUytrGNBqqBajSP4EXSxO7FSlo
5p5Cd+mPTxOuMyngiKJvFCk+0zCFzjFwfSP0KQvO3hv/xRLMmfVlp1b8EHTX1p5btt1GjOJsJFVh
gawXmrZcltAx3qvyhOI0r+bABnUbevbKrtGGix4qyiDteXwwcsgbIe7IUSgOUO8mfsf3/WuVpmMC
GQBd4YXyu5jH16mCb758aiwr0nermBvrQhQv7ityHWM1bNzQ9NfNXrlQNe8SQx4vg7GVhRo6Vwbw
NmL+9Nn1RmtFV6BwRUVMs7tYQQoeXOB6MogGGlHFuqGd85z+3Uc0wH80ybDwMdS7IC2fcpIvf50W
ABUVU30Tor4NHwSeqWJ0IUu+ctvQ2pFH0ennShlZoAy2hkCcyNoQ7IAHQxDrG67kW9BJoGWb6q+g
aFvm9N6GtzK6WYESAsBzYxXXZHKFJk0CIHRzTnCa0njVEh2hv7gk1jRPM7t+JzcskGnymRNKQ3OU
Z4jI1fsKtRDrBi+YbSdAou48IWmM9Mn26w7RkAFf1du0jz4U1WJvgvUpFVVid3MPZi5HnrJA0P0n
EG0TJJ5mXKwGxWBsx4e5Ed16yIrhEKtCibGK84wdfMKC/oS0VUUPUPUz8s4e/fhPpyPO33XFpMht
QQjKakj8+K8qHdVFwAW8Tx9alS5Qt1Pk85QMSlrTymnPkKiO8r2hqiBvvDHtSBO8GgFxnVRQuNEv
+qVCIp2noqeYEiLq/5d2HZ2K02J/5OTAXTd72TQdhBr/4rmKipKUSXEjzmfdfLLj7MmSAghKJSsR
tH7IIdH/KlYK0/Qty/vZc1qgAcaF0zJg0X22ujPKeMeluwCMXtmAGPvIKyoCgyvBQdV4vT9mdt8c
eN30unJdzWeCTcrTGKYRFAbBdaMdgQ2esnNJabtioXo2c1CC7AY4nuljdU/T+xZTHp+0JB1ynQQ9
zxEhsji1AhuXx9A/zBM6hDz+FJ+Zfzqsi6Ry9Xuw61470JvF/9gcRYE2/OuQvpGGAQJvxrdM4l1E
BGVUiPDOAJkOAMhMjMerq2LD+il84Hks09G9y+lpW1r1/R8Qn5twpZeFmyM4BxwTQjcEq0tp14KK
/HYYTg9xXsYb0BMHySMTqdXNyly806Fx/O90S0vHm6I9cQSsfzljG7otUWZghLrbjsQw5e5dvUf8
20VurAndO8ernaFfu0/nYznUOHf8ncgEn8DvDQqc1BgidGYfYuALHNlTwQGJMJ/ulFTrH7aSj/bo
d4maeShhct5n9AZveangNnU6LcICFcFngxhKec8/3vyRsC2X5R/45yzbFt6QqgfnqsRlrh8uYXKo
np/KIAtJm56DbBSRxqtvam1/z9gAUE9Acrf26Yb7aXxW1Ih70mHZX91rU6wQmNvOGB93MIscHN4W
9Ah1TIYf21A6DX8IFeuWnt1lbPug3X9KJYdEgmpZSyB4Gh8jt5gn6GQc6jxOJZEchkwHqj9E7/DU
REvOwodt1E1pGtPEsSwt2joc83eGhHCtFKSzZQ04EBuNCYnP++qBj9V9ZWvqgnuzcUfX/eN+WGQX
0OZ7hxt2ytL6L2DuHJtdVGpJCyec/x5n2Raq7QouBcLvUhsrEgn6JTnvKC8YC1QYM+w5NiC7hsA7
8bntLOypXHYj1RS6uxmlpqpt4sZDPfB20BGiiHPBVTN1bn2CvwOs6JXHtDVFHonUJ8UpugsGQvRm
m48LsUzmb0E0r/nq+B57A+PhfSSLkcExB1joP7XCnuCIepr8Twe+tGPL2uB6WdUMAJGjwN0XdBcL
uHzR36dXV/V0/ki6c4PCI5h2YE4lH9ivjBB918n8nvKGiVkoVS2XVuCgOibU38opaLkUZq6P4JM/
Gxtlzs9Vo8zh1t2wzU8DEwh+PCDh0OBvlKGhdjKy6tp9QgMDTf0n3kgJ/+DhgUo7//7UrwUFVkrq
ZtDNdrHtXuHfA3ttO8uqvuuViSMefCKmdngy1RfaigG20XyPkrY1YQ2HkVk2Z+hpSDg+NAEO1DKv
4uojyZNu+0kN5FGFyCZZ4Teb5VKA5NnwrV9QkqdStPrc0lIb4CNTqhW0yi6uvATcdPGE1Cs+1BSf
yQmtVMAcB/POtPSLCkx8zYXPjA3PywkM9Z46h+a9EuTNdPnkC8dHSuksqc3pz8B/R+4hK/utP1c2
4i7e32qDFD9mEX0X0ocyleEVH0UtNFVuogwiXoFQ/e3q0OIKICp2hsEU7/iAhjZainCgXipTigQn
29jaSE5QKvITSRJQjnVXvzsw+Z79qg8uZyiK2bBVxeFI9AuvUaR9YJs5NOsCDTnztdd6BUtRjOdB
pwX/e/tzXq0JJX1K+ZvBnCHJsmX5WHIsaefo7u6mj1GNHmGEg1bvTVF2gjBIWH0bHK42RL2PhLy7
3sV9pCBqzt2HSivmfhwWNuxs8Qz5T4npKk5Gv9oaBP4qBwLc9OvjwstncaMQbuLUXo5yOfcLEytM
6nJqXDAEw0NITLgI7gesgbDXQALx726EJ63dxeUFft/M+86Jt4glpgtK/G49q8EcRNI597ZSlp1k
RLwJEyyT/paeXGlLvZIn/3tyr275TxZ2Db9H5hMyJkq2Zb6QBqLgD2yW/9g6eGywNOiGsfPPITHC
GmLRAUFdAOQygLFlGB0x2xSgjD6ZK+RJHHxJhrvkMok2Drp08CRa3b0js7yIiJ73wrOfARN83wUX
6wHTl+H/3O0D5381BstSLFhQ8p8d19b0YNJU7/XzIkh69qbVjtjKqltF8HTU2XNFv58C0J9bMHxy
xIKj31pCUuiY+yFtPOEMwXf43IJ0VWLXO0TydvIwXCmoWw3D/uMHwaogR1Wu1mA7gfJoyt509cWu
7IIclJd+mZI2aUf4A6hs/IGa5XsS7jsiW/1aPVcDSDrgj0d6qDN0zGHXsf6HiTre5Diw1lN52U4Q
wLvLvrm3fupr7iifQHYBMGy2b0r9TRNq6HzZLV3wowwE91xXuo/nYsMqoLhja9mUKOUGp+VbE4R6
yw+q1RKSEqW8HSTaopXRQycjGhCk2tLmRvVDLuUs7lGigUfs/p7G3JJchAjYSyO2w0zmxWCbnU7k
ue0QiVDMjYV6V+efOr9K/sE9tNhpHNdag9svjOd49brkYJ8I99+WhD+39FjammNl/L3uVeTQtcS3
oskWXOsGRWMV2C/qy/8EbIXH/JqE244lNoMOEeUAoqhW7Ckxmd34OGLdTM7ir9SPSo/hAxQMIOZf
BBNq1blqi1DXVqJCUj018zW6cCdKszwQjiHiZn8Xq63LJJMCscw/FmFc6pV310Oh8f21Pg4xTklx
NmhYkE9BAGf1DoI9AolTLU5CdHV0BC7mLiriEsYHT/fT56CUQES3o/vyW3Fycbpr04b6vpdrw0kW
Z2h8syNOrTtpa3JIWhBsqs/GISsKh9eN0EqxZWVmWo8mesMITqCd0T4sT8AaRpl1tVbAr1SkjobA
Z3iBkTC/FE8sWOTagseHY3lgyTn1Ho/YSnwzmQOLnvxD1Sq57OU3VnKN8H2jYOBwxDGq3kW+B1r5
jgnTFBZXNEP68szyS5/WdtbuG2cTOAF2kgxobjE62CyNzagZM04jeI0Ci0j/Ap/j1y8kkaLmVzta
AvrH5rLMLWWEO0BOOo8n24VbFpzwn+NWWVUWzIYfq9551ybFioVhkcB/m/oN6fsBLWCENd1qUR4k
dHGkLlIn72ak6p/j02QRiiqmgyEjUXmRYygcHkSRqzrlv91OWlhpQC7gXHhXClcBLlUnExJZHdfZ
EthYUaTs3A2pK2eBFygebMHy9Y5lLV7Ai79VwTtBUzgFZyZvvH9U4YMiPaoB9WIQRMoYLtI0qEvD
VQC5FYp6gW6ZMTHHX92jUGoPsQ6OUEuzbgHx6MyI47Ruw/ESFZCu20I9KAaiZKOjQ+60svsuqckt
eXa6WqLBaD+mWPzUAuomm3KLG2WZ/iwbKOmg03ZRVraI5ECeNbMEH5dhMjoZmjm041lImBGfpOmC
SKdlbitiDNginoWMRsRJJCsK9SzhjFE393uGG+yz2iPq3HByr0GzeUef5sYkLtsuHhN+z1dVPxjL
WZD98PuTz05KEFd3/WLJSK4nQrU0buNzhcJ/iQu8E5VKPtxvIeDLUx+2pgskn5jIgb/xb5LlWXyZ
KlAkJAAbssabKLxuy1KfRyv64mzHMIdQdfbuMIdLQTh1wsKMHmZM0j9M31cXMDJzhnGGQn0mzmAu
R+NnON/iof/WGaSfqi7ITxXiH0jDTe5+zNVMr3PFhEnKHDKGqyu0cO0csg8dZIhBERFb/7Ff4GBc
cxZoMPsZPt0C+LQqRpWWkhfe+rENBZ5U7nF/WrENMZe17b2lg0rPu2szBtJOJBZgKIHM8XhDQIpN
VrA+RB9e4vz4dNiBoPOX+vVPgv4GBcSssxNEqHrOyz3qLxFybLk6c+tWskYgz3w6ol3tLApjQydh
yMSBHTViqX5InKFQmBsleJsEOFnD/EzDC5lA8jlNHdde1vbNh0/QtyOWu6mfzngK+fiKEWjMLHuv
w/vcxrRkHS3ujBEky9BKwx2vPBr+8AOh/R6LjVqe9/KxpQ5y2YVv7AMGldYZgkpjcCd5gLSdw6w+
FUwHpL7eJnB3RnUWI2C2WXBC3IywBQQ6ujCb9i6buhSOe5lw5lvrrwqWnCHVIOg0//ZhGh/Cf53Q
elkTRiBFn4vuYRkkALN1K7RLyswygF+lE20egnnP9YM4pomy5aiefIs9JUP0GtePLDiRvMtSBMKf
n/LARbFjz/m6vfnFDnVaZZF5A/PB5A9EpB1MxKb3SmkTqtSHRHDmdJzhdr+HxqA6mW5VmqTXYcT/
E1cePkiiH8fBEfLKw4/p+LtBk0Y4uI0ucIFbMJSzP2fImTC7sg4DnR0MgFADRZGRfaP8Wy6o9ins
ZjDSfRaTnZRIJOjmn0JGMGe34R/0cj9VzSh/KPYfXlljJBJWZF25nkJAeqdGiUzDn3W2mYQ7vz6o
1bgBzXMP5EsukYYPwG3W9vGxND6N9d7LBuBbuxb0+YTZnYmtyl/KAg3Yvx7mTJPIsy26FRURhYZG
8iTns03U5WVtBaAHAaMPy5gbVz1k4eqGh7ng08ed7rHZ0rc6nHwdp9/nfmw/A6s6uRHQ3BFo/Txl
3VKqCDWcZPkmvAIoIy/DFmDIizvmyK40Z6sZR2E1k1bEqcPYRnWMHiSASXZchamLhZfaiMW3VuiS
HBVya6iYBfidic4GwIPfyPj/PYTQfjXF8PvRHredV4hlLfQozDkWyQxtnssz086Uqg8a+9ruLsNj
k8BJlrYem9/ZmQ0WzqJGe48rH09mMLOy8UOGT0Vo0cCfc1DlqsV0pSxGimEGrGhip1RCjO9QiARA
aTC3qHCXl9mFRiQWo3gDTdjLA+nGhbpJXRJRsmMb7t20F4o2S4Hm8InLOzF0dbMJS1FvMA3DSK/d
0q9ph5ElIoCErqxxjMwP0T1NHlluS9j5i+Z/8JiDcB26n/26MI7+tug+kfN2F/nM7f0s45BlXxZ2
mJQKfRrHn8ekrmgvXFjcP2iFzNiY9//AhjxcnjKXjf32DRRnZkFO5ceQ1Afee8T0WS/Vnje0dpyE
8buTnW54/bBwsgTtIrvgZiFQP0lptGC3yN2Y2+quIdqTQtUQON87rpPpVd5j9bq+6zxiPUXgSMOv
XrRZ0Gh/6++gtwNlu4oFicrBVYy6jenJg70lg14jujZotJgkFzSv2uqJSGZl5s8iPx2Qrk4acOCt
ss0hftXYNGWnKJOgAt3DKGx0aIFwkJlLo0wVi8LY8Np63lCdDRbPhxL1LbZYpKzI1qH5Om34QCSR
X/aVXe+p+JnM3vIv/gBQkA4NXteq09THlZOYxc/+fCmds9iRb1XjgTQQPRCcbgO/9oomr/r1JFIa
GEsLSZzorx4yDPMLryzpVs3bCh/m7tSK5+fJXEFGhsIHoykOmQxkFnadKm1TqZpg6XRMbKC/PAOK
9mtUo2km8PrgaTh7JNGOashvMQYzVuFDW0NZFjDzT+a/stqd0AiZbXhrzuCUdjV83Lf0nNOtguNz
E0CR4ZgeXwcPj8IJJvpof7No9vZss6p0gKFCDsd4XwIkASAkU2trN3UkkuFFH6AiVedrbXeAdOSd
jSvRsEdxU1OUalKyznjjzl9TSavQUmY12FwbaOSbpqVRpe2ilkKAdHceEIZJjV7F7u4w2/nO3JUg
MSaDbj9GZRXBnq78RgiA9Mf7qYdR3kr56uu1frawVufnEcheapjyZFCSl70ITwaXjYGSAXZvSwO/
jIqCsYAXiGfLakktg5FnUdM5NBtiIoY31S2U7y3dQRIcA0EiePhHwYezrTlJDftRv4DQzNJrIhmm
mjSYsHcJ0NVh5Xi7GGBrVDARdL+XCL3/Nc8aP29LggGKk1ZbaSJHWKRmQaj0a0lCRt0EMUqTSPtK
UxBMmN0DVNxbewRfR0tI+yQ2+iyCh4+DOlQv79V9xVD1BuJwF1JFKGUAR3VDlHfR6/EY13wYRE6l
BJFf6ZWjgOGFDJMZg0UqDm+DZSXZJp14nSAFd4GnbJzjBKkt+IbkbP+UeZPc5lxWlgZKD4uujU1J
gY01kpJK4G97qg/Azv+4yU75cv/tTS1OPHEgsr+uLaqlDc6ZeYekb0In+7chO9rOLNZEkOjB5dWr
ApAfzDe4zYAqPM/zCgL7KBVupkrOsfF7hrDluSZBrLm4HLu2sZ/7Berm0PU3PS/QZo37BQm7drU/
lvDdhUJ/rSzMxKBdxyb8qjlffdGqpOZzYWhto7kgHnxxqYCy+nbsIungf8/ll3kOoMYc+mJHEO0b
Jrb7U53a4cQylDgTTDzy5zeN1gsuOs+4tHsps0XF6YND7XW87ANLpn8EPeRtvPq+lSloRFHk55D9
+Zvg1HitQWa6mOIBVfJY1EGJEP2SgZgUUMxXW046uZX6axs7qjA5t29tizKpP+ubF6FZGrbk2hNa
sp772cf5YNseu+mTEEi5qxSeOX74H0HPr8tL0Z4uS5vLlSzHgz8hyaStVqJtP+FuIVkpuWbY8oI9
0YRKjTCxldL6hauRYbUNSkqjiiEMiz5xu1iypS2E7u7kb7ha0xzfAYpFkCa5XA5Q9IfzmrsqvR+G
+DmJnNi28kZKK6/Sofp5CEH3Y6a9GPgDTwhhbw/yXw2S8yIgcL0HGBni5hRBAPzseMtsVzqwMQub
ShMrHDcFnc3e0uymdCjoP0l/DsKbHmLGKG+8cM8XSvlAL5rTKXnkVDOnT6P0pYwW66bz4S/TbJhk
PY7T8cUPgIZ1ygp91apCHFu29HTT1v4GovQ2gGv6r8iDcUiMl/vsBKq80/MlJw2Lg7qtGGpy65wI
j8otts8kPteJJ8s12ZbE1AzXitT8Zzlb9jkudEp//4uUy1LkedadwYohXFKeFsljuY1OaE6f0oyL
6fqPV3mZwssEhqQWT0FcvqGE+j3EmruBKUih3JzmiLDSrazbwBBd6g+FHlY55TGh0EpXg3ablDtq
0TqrCkUeqJR0SAqbfS0+QDQ9t0B9ri/wTYchTFOYAsON5hvr99j9kp2ukJDeDx2qQSlBUk0Rczxh
+k7w1rhrAJojk2UQt2TRag7x+v1xVaxuBHkEs8RtR2AJxO3PkMlObOpeKzz24rvgaQCxQ/+my3YL
RpiJN1yw7jXYbA6722kKt+g8tLwFuZ3st/hVCxqbAEA6UzYdeaFzNB1uJWCLOPuK0Nx8FxeId7UF
hdY+jr0CyaNCddtlCjNCafmLZf/SXRnzwVDLZPatzKGm8A+vKIKSk6aQERZyVkyN+85+SS1jAqMN
teQ8FwXxqvOmkbs219YduYRZIUIcKt/5cBVrhzSSo56BYyq/Vh+Rkoc/T5BEHXARUemCryIoK/t8
ZXEuDke0YG5DoPlpcK5wk2bQhyJCCrRCU1nhWtiIOJRU2DchSHXTWW8CoDMDB3VpnZ3/tgzF8zur
k/XFH9K7oiXMXHbRTwNsvfcJD/8I+GWyDt8dqOcEOCII99WRTPBLu3GBHyHssfWYCDRrVbRG6YNd
eEp2NkRHIODqn+A7WV1KHSwLJVXoVcCsX9WEloNywyEvw1fwONYTO+DB9putQGkPbBjF3UWOo1R0
aHnpHU7UhfQ78zmhBOx5HYhQr15U2yIkp/7DvYV2UTGihAYSrf2eVkGRuVkuPFmGVt+3DqY9RQ4N
nFivpL7hTSbcygjajWX0Ht/pHEFCOX7WIe9pJNziHMS5d1kBuhPJ55rytvMwZL1Kq6HROoX80hUt
+nXL8UTULfyTxIxW+sxqul1pZFewWSy1/VXH7as7e7ULU+7QqyieyCV0iggOhwM97sZNM0Tl+u21
Iirup+g2YQ+kBhcBlDV2bPRhbGOCREpN7eJDOM6IPxzsQIblhNc5erZMrC378v37mT/wBhjAWsv8
xuiZk8Eogkmp+OEI/opVTaNpE+EtKN/ormJjyg6tEE/xnbLSD/5T5nEvhShclwJG+2e+Scg9u1ke
gzzma61MhYy9z9CaZBso68olGkKBA/pFBWvfXNV1gWdkJ2Ywyoj9mR7AnLu+uhlinqxcj0k0s/DY
UmaL44WVECS5p6B0DDpJ52tFTTW5tc2ElQS9y5cn0VwtHtvI5o/VNLTdLmuYM6k/nWwrRcvYaUj0
n/vSQR/Tc+qUmZKqviPWxhCIs4zzSDXeWTUzymX4TIhdA+6I1Ehv1WIKWjJQ/vO9mqpFD367+l71
ONg2IMqCuVOnLzODUZwDbWXCJF10+4+tSPP8Jh3tFEjRJ2/rFxlv+vQCbfhNEfqRSvkDnytyA9Gk
+27SVD11uvzICNEhzwRIa42RVwuvIoLPjX6z+6G4Nf3XVH2xLy7OYW+aWSJZUlDo+TD3mG0422Sy
IYUv5XXRpha2oiqfFA+Q3Soz7djcU6DmLb8v9W6OlIqSj9dIJc1l67icsW1NsHvkY4VRIWywXwvo
3HhugHW7LiBqwvixhx1F45bCM76uGZ6uzeX0bNtXshD2ixbkpHLMVoDZbWaImYrt18NRBNyrkx+2
MqT5ho/d8rC+Yhh/DLxp+HPboRgiKFvtBYd2APArHYWCmck7/KrIxQe1nsPpQ8TLnKrQSQfodvRd
DzCOq4UL5avewJh7/6DbCm7GC38PQjxbPBlyLkm0dMs6jIo/T36x6UMFoDPejUK8RUI97bV8a/GQ
OBxYEi4a9y6YRT2a7RIk96tpBFqRfLCeKWwht5tYkmsoSrdzssZzARlKkeemacACmjh64Q4V1Gt1
PNOir2x/LDIW6cS3dWwemhKY0W0x0EWSDBKAyZcHBCBc6+8a0dBFKrshEFceL2D3SOXuTBTO8k1k
uxzgoWoXzjEGhOIaJTMD5tw+BGW+77n825qogr7/QeTMy5lWdmSK+aZ/mORVBdYvJsIOz2rcVMsV
TsxCnlPCPyIOFCDqutjUCDkNOuF7bexL0MjjLTdrkqGaYCmo11KKatKLImv+i1qErNkpEjH+Nqbr
qsi3eYmXxpsoK78n/s/nH56k4meAnBYpvAMvP9oaZ9SkTaQYG31e5DcnDFidFUTYpt0Q9HzVMIgx
cyPT2dqQFDQuj1lEYICCrk0IPtICfOPPFw9+HJyxuwXnCJRyoniK3nxprmAVsjsjRiZNE5pQdQY4
Cxt3hK0547xIMCOqv/T34t9uG02wHOx1sCJ+2cjn1qeeqX3FH3gEcb4QcX8d2RXdanBVeKQfsD1I
oGZw4aSowGwYs1AhosCDVDIV/BJa1cXhbj0no7/D/u6td96Aqjz9Q24tkdTaOmi/4WLqXpctcduw
AT5av0DIyI3IoY1Fa+OcwEmHs465MLutwCTabLbfPWAJhjvu8WujGDaW+F72d6+xs/yR/3aQ6VUP
pxBLGo9lRG7s9SkzYc5YOumI8D5qaZ2DgMxvdmSzNJW5rUsV2S8qDymdjjonB/xJ+fzoqrZxCQbC
vaGZvd8BtGi8msVHoJW/kwIjStTbt0C/d23gtuhv5VbkSqx/SXNEDfeT5mpR4Y4YfDg9M9pvmq6Y
Vb/B8pRMrIgzwGsA3hURxwIm7Ghh9ryZ63Xq/7fom7ay4JLu2QWDoqSco1SmwKX5FHMXwQ4lCgT7
RGsMFUHTpuazSjfXZOulUL7F1i2Y7PHfnDtczqwDJ6a/dXc2Vx9nZcSROUtRuDdV2sFteAXlkpcS
v0diuFv0jSz6FTPvhMdvJFS7uNPyWWsbyGNwHmzH2AW5Bp1Xp1vuuwe9LoYj9a/LndNJE4robVvi
4wZm1C8O/aWnsXoryJ9uTAuv+YZANG0cd3PV1GJKGjTylXbK0r7uo6Lx7elODaBVO1v1B9GCbrDf
ZDx0f4UZ9zp3yQ7U7WDmQe5IDXbiUsEvQsguagszquLVlmoAllAJ3tt2GdbhnbFJeBogeuMRiFX+
rLuTfWID26P8ux7ew8+O7Mxq4wSRpf0+6eBWoARrfZ7lY3nfcWNO1BofZ1na9MRShF2ud8BMc3Ex
D7X0r75v2HXwEMagGYKle9bdcU++G1U4XIBEdDGVNHSPcTpSgvuRjixcVBmQpXU0ZwVfb+kxpTTo
2yjV8yVVFESo6rXY4BENcU1ZaONAfEUeMX19x7Fwxv7rZ7oo20xICXJRwwyiC8OFGuOjdP7n5H4A
kSpIiMDXq4Bng43B357seOr/Qd61vcv6Jgocwh7yCSoIne9KPVJbxZhqVmV2ylV0Pk8/yozeF2qH
mKWlwrLIr+tf39BbPHLqOkbvJkFVE29gUYs4+wGjJKWAghpd/ImCyyU3txvQ8A6q0WRfN9c/iN0V
T/cnis24ZLludHCmr+ncuuOreQ5mwE4LhUAlimjLWiikx27ufnImdq0PfW7BDTO/v5bHq7erXy7i
DAK7tkyxTsWZD8MvW+OVty/gV3f9VTr5BXxsrAdZO3lST58pCKy4NxLTbn3cNEABhGr7Qo+6YBtY
6Fzsyzt53kyBRX9zPN5VWlL49WB5qUEuSbYQdlTK+bFwGyjWH1hBuJhe6KU36n6/pxWc8DfWOeG3
o5rp27AZ8Fjzy8wuFuR+DnHKvp3vnxQd12D4iax05++gHmKc/6quFeTUOug42oqNmwKF1L9ahkGc
fqjx4xUF/XLlBmPCAxY0XaXF3MY0QodGfnmp4woHEZWet/JcPWTDeXSLCUsddBft0xU5EpKbzTiQ
LHeQyQ+uJYX57onvA9srYaXG+mxkSx+ol13sF5vpeLSrG+96ctP3eTf8/UZVcLCMJ0KGkHiWjidV
ZaOWmWH0YmqJukUsEc8vNJEXYpsH9avJ/wvrcP09wQ38sSv64AoCcG83k7VB+G5fTBDp2dMSKI/X
b4e2qBEgZ/dymOAZQ0AU6NOPK+ItLm/R5q2ISy3OChLsT+npRN83eCqyQmQt/kepoC2FRxFzpViX
6mUDLg2/eV37Z4GaOPWI1RlpLzPQTygqAanVrTRR7Pg1+TUI7MnyeY0eBKnLbnezjsLRwvp0nuN9
0rEza+QnIAauYdVAY4D/lkeEFrr3yEQeWz8l1FrBsR7q9bzjDkll146dOaBed8e8LY/huGK6KyHg
lToimxktXSP6avzMUOcmtFp3coQeazQMVo+9m+3AviMON09kH0rVvY7zsU75E7CKMo8p0ns8LVJJ
416F+YTln8YK4qXIMdj1TLtGxdSsjMPM4dFWa2dBWe3MSZ6Up3ejaow3inWR2t8xmy3OPfqdsEXj
2xe2en/0PLHzc4229AonSTzbmJKImWcCn8KPlivO4RIWfMaRfVtKb6tokOSsQ2R3+KRDJTpqJvkK
XcCXF5+5tiZ8p79WrQQmQXZYKgv9g6pWYI5mMnQO8KHlEbpvjltGVb7JiiooMSOy99/1OAMK/390
OZKmJDFHeJ8bfDvVK4T01wRABx7/P7++P+5DTH92UfiY4dI6qFwprBizA5Lg1hDZj+Iw3k64Q/Uo
czfKsnN0iccA9e/44H5U+qsBz6D2fviR0XQAKhXz01bp2RtOBiFUzX7jOS/lTtG0Iqg/9xKdggTM
vnuH1KMkfS4+llvEC+kXhVOxYg9G6h3epx2xJKtKajpe2DZKzJAVETznPM3tDPH5Jjn8tTlzeZ1F
HCuyS/lIafuBkZqwjMQ84QV2sTbw5+lO93Pclr1DA4LixpRs7WUQsPXL6KkxQEbg8vttoXI7Xt2t
WjOToIJUHVWWrzOUU64E0ZwDdGAKVQfRDAO1aTL39pxHJIGEiB2dRE8zcXQh3ejgisHCXbDPLXJ8
CyND/lrZyWVdpgYKyD7QPszplRCV4vBq7o/t9BwPCrH57eXqbd5CMiSZmUxRurXECuLly3Jkz6C4
0m2tn30jy4/eVbAubUCZN9kfs94Vrfhz+4IdsovZbC0BUCqDmiuHtuLnuoXSVZQSETO/f+Rr+Bw8
lIhm3jVdQ2spUnwXyipgpKXa/lbrqB0XYTxPai9725HO3hvIAsJvXo703bwKbPVdtTirnrCFnTlt
JP6sZHf6CmT12E6CZJuMkMNBovmA/RzvvU04QV3um+coREtrIzi7UjQnj4l8VIYfDxluoA3In38g
GJ9uWRiho92X0DC5Q0l5lPZO7Ua25BVnJB4UcuxwlFd/MV9gojQOXMA+5tivbAuLwlPK925MISaG
zvBQPJNJ1X3FFWhJ8ZDXY1H8uGDA4LFJh066GW6FhSnLRrL0pX4E5L9wBmAMmQAq3jN8UOOuNujD
djsVFuqVSXrlDf8jPK9y7bj06IF70jwKph4MoGLlwTSRGVKFZvBOvTluBy169z9ssZageRKFV4k9
wQYf/C3EtQsKMKYzknVdtzFdLNdbNf43g9SDSJfR/VsQXel8dcUNbCEoMakVizaBmFzS6fXHB4+3
EtpG5TXOLeB1hL8gUhM7mOtyjuRwohsQT7iBRBtPJ/TING93XxOxL9Y9zTO/d1bQftIfI2FTsU7n
P+O3yXsXu3tkW6e8TICPNOhjbP2aHq949VQ1bKXBSA0Sy0R0/lDg4eimqCoSKrJIQUzpyd4L8LSG
2TNQmfbDVd8AdC7PyjrNCoV294cj6bXOVuyaEL+U48D57H1nnq/8uJ46ZK7NolNLq8Qxqn1G3pfa
TTLHKaDbmf71H4gmL7t+7EtwZS4cc/gkMYQtoHSMnAWBDpPhNhQapnDtMsCiF0+/dBC7Fd8ydHMn
bXXvxr6WgTy0yRQso3p5yTnVUHAEorIsNNuzZHLpAO9aM85UDHuM+JysdlJNHGXDrrTIm6OepzA6
FWIcDJzxGaCvovLH6FmA9tuFK8IXuggh6G6SpfOjypAE6/PlFvAJXpuOpbfRRTTvtaTyI2C9sbjq
y64xKGBziyd+t3MoHm0PiE3ID29jrhz/5ZDB1u2QFxLxiwLZYoVMBWTpC2bpPC4e85PjF3TH8h17
KGFlqPXPXGGqeXAX2r0NAsMY64RpQshRqADfaW0sKh90avPPsy7UjKiyo3Hx+YCXq8BLZgsPRPeP
O4a2C/ScK3Jm/wCntmNsEEaytcix9XNQc9DXXQ7dZewv451B5kPQBKUW5yfbi/NrARmCaEzhKI6y
1hDukEjaL2HZJnLGkVoxjWXV5BPI0z/6pVp18ER0C36VEGoddmUFHO3QuGet3ylwey5PYDzCUNfV
4ZYp1eMohO3QutHcy/0btejLIJ11Gp/ohBJUpEYyMDa81iAzsEw1knawdKeNvpSL+g0qKy1iPJa8
iNgOIYPazdcjB2gGT3b30riDZ7RAFYmJqio/Km5ZmOWaJ6NIqkXYbK2JKut4k1PB0CBj0IFBbM/C
irN18eqsSNreUD/SkeYTTgdHNJbmmdKQZDMa4fMJ3dxAfBL9kGztexGTQ5HqEDLy4uWNM5nkHSuU
E462kFXyvZ8oelFsZ1OmFNt182u0RNr/z/5VX7vm14t1UBWF1iFgfNm+PdXq590qpIiXMW+1+go8
iDpY1iDgAABDnzoN1NOWs45UuSjffUoKcWiXlBANoxc42Qwk6dMYmGdKOxnUEPLBnM/LBsuxV3Lm
cfGlBZKnpIAh3KY8oMjm4ANO/6peJvJUAKwDiZU9RM4C0FhZU+AJ27YeZkF6ErlqMtatKC90I1k5
PJJUYFFXu74PWVKLYRB6Tj+5OEN1kRsUCcWR8tiLbblzNwH56k1gpLc2BdkZPKqSCnl8//OBsPzw
rRoGOOXvcQ+V6lc/bbnHwH57gtNxlRqtv1DDJ0tuTYMTVusacYM+uUEvy+UH4+lH0KMqiVHSz+U+
7CB3IISBoHcIOoBZa6tbrpuTiwcurfeMcUHdoMbuzlYiMlI5U+wGo6yFmdMvo5GUiKMMcVgCTkWq
Jcb9p1MVUG4ity/mFD3p9kOtiFBgotkGyxdLLzEuK+IJOElMFAEKxVENQCaUCk8TfxAs1UR3cdWk
EQ3XObf6MqyPwp92OOdi3Hl3txQItlEuoCIfTGTOskPZU7nb+CSnMmWcBvNgQzvLKpiQBm3u+9v/
HZq/38o8UfabQw621k0tjpe9mMBaEt/YJ6JX/XYAYSvp5zmZk8pQfCA/uyXrPSW6JKs0cCq/gsG6
UWEJOkDdSiREYxIa4iANgBfRBD/y7wZ2nCRAH9RvcYu9Y+n0ij9kgrNFKnMqi570i/j96IuRMCuM
Ew2P+eb7sDnBG0b01tILIZAieCesmalpV8TxiMiAYA5WldDgHuhG8Tm/Pag7D89MmOdWbR2NcQ+o
364NPVK6yDIQpZcLElMNqvWDXT7GUW098OLfJcX7pF7J5x9bvYIyEyQUKqFTMIGtqKE3W9Sq88ad
Qozaxu9bg1uEMwLhrQ86r0/yOO1yJB7NnkKseSQ0ZEkKSnoMONvijzxLtW5PcN7xyAltuEhmv5QT
pIfMPVUCbNUoDUkhqkMMNQuqM4UH0ILsmmxw89/NRzLjBJZxKZUIl40Su6sr+47vli+e9B4msTq6
r2yaiBrkkXnUuKFOj7axj4JOJiwIsSOk0o3Q6BE1+RDK9DMzGJZN0TaSEbhK1ITIIAstMtV8WXK9
czRuKqAJ07AcPwrYxtv2YDWhLadBPe8QuGjOxk9sS8kRINBAivEP3Shz5i0uQnOfYC2blgr0RvNs
8ZeL73udop45574yDqkYdbX9jGapKxwt60zjHwl0Tmrzgx3hSavyoyV/X122DCFYKYsaPLmeFOxx
Zw0jynT4KXyZNOgDABDA2vJEFxftWkZ6cGbotnp4fq3au/JTNngm3F1OKVznOluweQIX3Ca6/xMu
AG0bf1ammOVEuQhIbEdrqjyHx5aA6wjeeIxA7nD3iAFh2Oy8x7cTq2tml7tNbiKpIaXVB1fSLmR/
vl9+gn/cGmbI3iWQLG/FF38rTJ7TpFMZBAsQfIUoNS/7fX8WK5MlahfPgDqRf5AVQ7omrvQAuZE6
r4kHELqPa5SaYfm9sZrIGC0uVoq09XDUINS5+a34Se5yyJTerBevM+egejlgHRJcNtjRXemRZOxF
tVu4qGhRXbtSkEzEJICTxi3EFyqsBy1wJCfzhf68rjo9pgOVhPFhCpuLg0LJzdmQFCjZex4zpWVv
NQ48MXnxwE4ja/AmE9nIu73jmH/F9AeiwsZNUz4SPVcKvpzC/AenWpqFWxpstNr6mPXk1iYdA5sF
V7+2DRLjg1BW/AiUbzsTUkIzW+07X93RDdkFwT/AzXfeKAR8sCZadCiVahomw86xcLKsvlIrcdGj
hflxRrbzPd8W3MHgMyHPT615rHuTldGYcHqMLqn5BS/IEcJbMMORonmWPo7CrXWXZiamyH9W0NUM
MPL34t58AwvskDQmjYiusXS2LY0aj7r1AiRzJXuM4Tz5FxyGUlFJYy4BT2/7lx4ugy43e+3Ua3eI
ch09Cs97DEiUfEXlNeP9xgzmy7Jkz1Nzo+lrk4hdOHjW7Cx+BJsUsQrG8nt1xUSS9f3jRsuBXed9
BfjSTmSjCro48qUpweYL2bAOnQL0CTVMEwe6w487DS9aLvgbhSg+UCfphgPOB+y8auluO/19hMIV
qblZ+zPxQbaUXoBlIYVYUFmzN7Gk6rcB4T8WJ1ciswmd/1GPb5D/NF3q6XLMEVuMm8wegY1TqlVI
JsfBDTwQo0yO7GM2ZdkyEB4fbfJpNu/+i7LRwKQfQeIjMPgxPLQVtdU0bub7j4j8AWxgfeMyOnlv
YQ2xQ7+w4zgUxAInF043ngUzYZIMpuD45Hop5vMjm+BCPa1eEEBjXP3A1tW2xgzMFQJ/o9smsOsB
YcCcuDIkcKou3h+dRXfBnmJHwGJQritzHuI2bVWgByKo3VyRrV5Fg1qSESV9cTNFUQGETFGnjpgB
npxIPwlP9cnKu6cU2Fx2o/VJ3HJ7c20bE6DYwGuLL9Ps5xHBmf9Cy5q16spw4GwfaVPGj4wW+hUm
4JtoP0fFv00S5JhP/7/VuKWR2Bsf5QJRXHYxfhiMEAVQauie/cWz+VEjwH0gE3GmlVGpbmpJjhAM
tXLqZY0wIU1W1hH7nyIwvyhtXtm538s95OFhdbuBY4q3X0sUhlzlCghqZ5Ac9mO59v4naBPucYh4
JbJ4h5TKHYl92jDMQbYKoecn9nEffDEESLgvtDXZVfW9l3MxcypjwduBPP6ubi2m7QFipOG1TNC8
ICAu1tCm1A9X/BgSha4zXThbi+HQxhFYEMc2Mjl8cCEQSeuP9taEwxq7mUP3ZtCDxcUvHbMO53t9
J2jNyKv5q8hFSeKwRKVVP189zN+8vOLxIPWwxj1E6jQlswSAckNjioM6M+gCMNs5HlEAve0xS/hk
NI1UXZrjFUv8j8jeS1mlq4vjeM7a5mXkVPnKZiWmUNpwQf4kYqTZBFiXnHopu9FOgLzE6Ol4FUMA
GPNBwtT3YjCMnqy65HrhRIt2kWw2JpYnvm2aUoOwxXfLa55afgHeleEk1pOwM9yUGvkmemHbOld1
lTd+iLMiSSgVab9+yQiQFaWvAJElJHSCEnbz/ipuTwPeKNdfiqMT6h+VayD7IX1I+gYPO/m/m9tX
sAhoC0jruGj/yY1ze4YLaXAJKp8oVoCHr7UctiyOdA+Hw+tHFDdWssHa+3Wynk/xIjirAP/Owlwr
XPZF2b+LxRgd7Mzku6MRL91pmFfizD7eEy+kecOL6JDPkc6KLBGS8nxwxV7Rg++QItzu9CC7O+EY
/Dlu3KUnUPa8DVLzVm3m0mN5qxbEHd5hcikRqonpI5VLkzlO17OXovhPU7Ar7ql/kdfHULcI6qAq
qlUJ51PuDi53TM/oWivHkiAVsY/MA+8shN+IGXr5+jYyH+4dcjpD/1dnLZFiwxWQB9+onwMn4uuY
z7h2p1VFZF3V+YcVxMCOXezZXh9Gwuw7D+EWHsuo2SWiuD3NPlpxNJStJMD/fPqBE84MBGT/2dCJ
45Qpq2E04c0R2OtVdxjw24DhDwTO7wRuk99/PkZfQj+2TKXlWUSi4R7TdlewtztSJZICcNr6JgNT
Y247vVJeoYgLmY1dVRQeiLEXu1/iB+bvM5sbDYzikvMfIxFzFTENh+LV238kd810ssiTc8lfF9MG
XnB4zaAa5zW5P5qDkgBODCMrI1kvYmZo75FubHjSI7wgjH0fSRj4dkeCLue50Cht2Q2qpDByxxkt
VVCuJX4JiIfzKkoGBPOWlwhX9/hbp9MqF9r3GOaANx0hS69LWvt5thxC8zJA7ZxkLs80kZlTgppl
guFk0cjlrhQG2iI+KzgUlI3H3PjVE/SWPGcF6BwTWU0gXECH8+d1vzAwBc3nmp8swpgYr6GtIrAw
poCmVh7eIx1G4wpiXs+LhbXzues1gfTiO10Og44KWZDyjwTXwp5aF2KWBHamcNAK4LDisG4i8gdW
gegld54dbWJujhk/QHMwbPVLqA5tM4dtstJrm2WGEqSmFVFoOGHNlY4EvRlcTmNOtXUUYnL9nxxT
r2651ezalidJY4eQa6UHmr1ql/CSGuvo1kkQA37+yH0+bxwuf5zv/ZtrlXzg8KrRFbewO301Xk8L
APLqpeTMBUgWn2mPwY7zwE5y0rywwdOkwzS+iY0M8z9qGiBXLIVCXYz+9jHRrq64Go8pMsiljuD2
/3e8MlANmg7+dC7ENTzbBFPTPDgiZFMle0PiHEJNI9fro3TGx7DYo7BC8+9grReNEJIGpbx1BSIo
aou+c0Rt9U2C+Rf5t9qclmoTLnJUCwu5Ff6HUDqbTWnfOeYUrrO86IHe183h1sCY1fKuJEAwKXN8
q08toJTwqZPBd13vqNO/ZRHFLvxfN4WJNSjSHzd9t3PkG4v9ROdQeeePiRMYTusjmmHZyg0rYLid
d5EbQyLEujB0BZNi+zUGK8l6iCoRMmyGwazwQ1hE2cSj3AU+g9sj4KV6MQZ80hAYgEzb6ggln4BZ
X/CydpjvAb6y4IyEvj0VS9g9SXceP/5GHpUEDf+SzZW/8pxwGaKxzsTOWyTeYuv23w5qn/hUYl6y
thE3A6SCCsRZUWFLKIT3LwSUjjkubhaajL8gLByZg67ysmWXLLOyaqUSMLgEu6o37xFdqCmyWc6f
+Nmw6+Tny4+JFFcvBKzQNagAejCA5gDen0rwIOWbBSjTvvYag2+hvKLvR0Hj+32G+kOp1Osw8r6k
fMH+v8DDz6gSVXlxV46cUZgdjVPl+7ozJ6HDwqsT/Dc6LR7cN5sZuDEF2kawknAqv8aTEsQ7k+qB
aKhqaroSElep55KhuocF2SHXtM2qSdQcm0R1nowQim/7B47oCwR4p/Qa6pGTOoARxSzj7z/SjrzH
gW9Zt5bp5tcg3MjfUemq2yn02cIO6GiHMEt68eE1CiqTWD/+TpgKyLsh2YevwOfDk79RQALQCQUv
WekdSTMCjS57IcxbLNR6Lk2ikgLotYk6LEQi4ZS+8DPqRd+wv4e2NLT2h8mNT4x64sJo3fWiMnqj
GLPburZppcn6UTu0r8uVq3DxN+X3Qd8z49Xx6Hru/bKTLCX+pv3/ik2bgB6P7Rrdy03xJLRBVK28
gl4MDZJlIaOLlNXyg4l7xlxCsWX5TV0lG0/16UVleStMaq4hbhrzjCTpisrbjplW3NG90Zc655GA
rfnmBuKAWYd97Gsz8fAwfmOFQRshakPLkfkkLjACgrOeftna5xNViQsCEZ39XG2ixqF1DYZzXGz1
DM+8P1jbhbTgJEwbNPWGVivMAcMr8YvNd37+UilIl4WzhKsKxiZDu9hhngDNoEMvYCgJVykPa53P
05HZk9ltcLwcmJWT1NzGBx5d3meSsTCHpySZk/XlPYcdBbWLoiiVWKN+6uaQPEiip9l5e7SmGoJO
/oTjwfKKaZloujiTOgvjUeWbFBmHRN9VHsJX/nCVOKtrRSP6MbsM+aDXYELP7z9WGbDXXR9cZQ/H
9ucqAxrFNumeeDlDU090yUWnHFFfX5xzyhYhyB4JhdoHFtNkDlEXhhtH1qg6K9islv+YfTBlT0AG
FjFS7lULlOkkBZElmcAv8xunsOYTTNC6B4C5giVFmiuRug4XASlEanpOiHxGJgqRUKpgdPt+2gLE
9L2MtdPhAg6yBgIinMS+gHNy/O9HzzJ2z/4zH6W3r61FGaUDwEFYE45z6yVf8sK6+BT8XgbJdwNs
sSi0ZcRDZuQFgO3k/GnUSx254KkLmifCagxiEJtgx5g5AXwilvfjB5ZceRx6U+BLa+/8RwYVJj+r
jSqIHRVKCMBfURXukV5Gbh0f2AFNBvlQ5UefBVYtG0sgxy/J8PUeffkOyc4dXNy6lhXiRmCJtwVK
QEjqbzlKxUcUlQZLDiybONNkXa4Z/QiPPAodtQUcIO+yyDTlhWbqFUHF1E8yzgkI0MnOHOIF6i3Q
G6CKO3qyF5anP4+3c0saP5WoKGPB4TFwI5qtaP/BnyhZLawrqyVOO5FR6rI8B1doD/VvNGtcS9Tg
HUlFs2/etfwpillfzcEHI+4OWBWqOFmIqZO7oNUf3RQ6nKHptCUgGpweIU9ufs5HLqCmLwmQrGLC
b3X5NV1iJqAEpmv3juFwfLaZ7EUqA6Uxqa9WZTLskz0f+r1SopcuTqLJq3DghDzzYC5ohkR3/1Vp
3MM3DxD453JeUocDXn4/GO8sv68VhYH9l3NBSfriDNxhjlIbP3C7wvXb4v3uy3rcLKIQrUXUNFF5
Es/rDNWbQLo044ptuyqk5D1elcxAEwvDL8jN/fO6dgQjuVmXZJbwbTmJ+gPj7mD4rVnOw4OVmB5S
x9uMZhdUgLbkrnpJmxAdgo8TvOa6uR5VXhcCo5SjvXZ77esbhVoSaT03x42EfZNDW6LmbtYcPb0e
ySHoyGHVegBZlc46Zofhc9JAXQ3EYsXVPlmH9d7SPn4oIhJVBZ15EjCebQUfAaDbgbwQY1NPwGNE
TJiMPs8V5xsGy8IcSYw5iwi6FyaJueuxgEZlr/EKeGVnT/UoYB+/cHOvTKfikg2dehzcHR/b0grP
IyEGLNJ6f2AQQrhvSF38rtg3EEtZX7FUTZu8RdYhcvWouSWgsJMMhtnW1GwYReiYCAxq8YzyQxjS
DlOl93iAO9OHY/vCrRGBckfdzAPKDoKsFG6CHZPddqETvBCS6u1BRYaXnluvVkZGwBk9sUtD5pTG
d2Glr7zduL8gb3kTbYGatiOYIr6TXTfizT6JM7OgwPlqDy6AR09tbhB6riLB3618jLuQxYGn1HOt
aLHxo536UeUpReXn+FwNLrjjafdpdoBL7hX37da+fqOkPhcFNpW6TD9L72vwd0QWYtvWBR5RCqWe
Xb6H9G97lP2TbmaUvqzzbdQIVOi0vAnJeMWxENoFRBDFPC62js+Am4abRH4NWiQ028QqpJhJLqVR
/9Uc6i2QK/zGG5bmdrFTq2XpT0QMsXeLRtGWIUkAdMipMYELgFgPqVd/IHGWLF8WJknCBvfZMO8a
T0ZTCUcBbWCGuWG0bq3+hYZ+bzgAjeUTkAdLj7ZF/vPl/4W8peo2W8md3iEYklTy6D8ECHQNcE9H
39e4QvlzLsAS6Oj+tiY2Fb/CDNKYQywuHMkygbOqvZu19ZPKbYSnKRcfvSAocr3ippi2lqtn6roM
dsJ/RAiLgKZwbVP2K32s3W7vhJMIvJaWBnozc9+eCd0wwJJMeh6Asx/WLOOCTP4lK995DolF9o8X
sKc4ACS43rNWU2fCrh6+infhYErze6bhVuz1IPYTKN7KrjKMl9r9mboEJzkWC39FZ5OxTup9HYzz
wTsC+NwZCxNdHVg51TBaTQphJ+dxTFP+3HIBR8tuw8yh41DL+KOg2Ukz+8tRgRE0Gq3cYtgqjulF
gW2lcn2yNPEQqh693Y0row7ERURv9dycGY1ZgG57np79N/ZYy9tQgOBqZPyNPUYn3FiTkELQKKkt
sTa87o6ACTyUw92s2Zz0vvE2otVsmCUZvU168kDnIqlSqWein1I60Yle+ZDkjFKJJV8XiUNCz+ZQ
ubJo1our09rkRL8Xx8Lrt0AEJaRhsEX9qBlUJxhUmdSm0BIwzTfvdLqvIx5wUUiSD+feY3t0SWdy
KtyI8jwaXCS/AySsuLQG7q5QT7XpQvuqoj38mHCKlEBwHcd347DgL+M6v9FugdWAx/rXD85FD8Kh
5DJouM18ayIpMeyYTOntdpoDJzOSJcpOSuTmaf86Mu0WdblLi4QCJDa+IzhCIhy380MM5vKM2Ggp
scJpiua4V4N/hlhJOF/yAK1dJr0VAhKL3Iibjep1UPODgQKX3yI/BSsaE0M1u5lKYibDNh9GCU8V
6j/ioV9PUCcMrEkw0S5nvlcAUKQWPK6pJscs4YtHIQ2H0deKtguEUZvywFO5xkrIR6WjH5sCBLT3
08XgWbEjs9MIqYajhWFmpGHDiyj2Xa3rS8DNqYWZ5vbZEuLl4+fD/OtKN6thRxundbpXtG3xv/4H
oUJVFKaT0hDrfdEldSU9WcJlvjt87K/SQ3DUQPrRrVlYPJXp99hsrLYtv92kB8yfqu5M5xgOOguT
AExHynXWLAPA12bRrSqYwQC/5+RAOJY6Vud3zvWaZ6CVhShbWDVr9FqvqqIOeFB96GmfZrwH3eXT
9pjyp4VD/LPaAAUz1dBwWlkY4VX23+5lDoPK+RKxTyZzKxUCj33/IOEWR8KTPjJwLtQ6Mesen8mU
8DXO4FPJWDJWeblczhnC9P+T3GTsGD68pFh/J9QUQSkVoFVw3FQc0thQ4XKIxafXJ6Nw22HuQasn
oTMnLv787l/5ow8FOvxR3lABnCFG7imjUVHPOtRYLwq5sq8uMG2vxZqubAJDOgm0qIWKNpXFDkVl
UlpmERH1OYRFdu66QusQGLacxvTbUgt3x95rCQ/DyaqvR6OdzloOabvjzJPl6YVA7w+fwZioRoZd
nf7dEOJnpHrm7HXBCNLZHUUPsLbnkdQiRbUNlW4JYCXOf200VtL4H/osT9R0fveyJuyuqZj8jFYK
AVuOuOn04asK20dQt/DPvBpHd7FHfrmodbtbhI+JXbBCEHq9qJjepOtrtWcwpxBsvi+8FRw0jRqG
8y/W+SlmH22qwN+UEhn2GkmRh1/Y4gPu3nVINpcDWae4wuoJFeq3nUHyzJd1i4FAui1BF/tXC9Bi
QSaGEaDvUBaCVfMKpJSDB2fkAz13xlGsIILgy3nKdSzvA2d4DBlMXrcC/t10HY9yAXELG2jPCvDz
tVRyT/3H6Zh5AwMgZ6BShbzrM8hoTTH+Ojc+YuAJ8OQr2O6mzQAzw6BXUIDspuMKj8dzb6lH/xuh
m7g12m+IXGv7DvacNEiAx2HdDeH47NJjuMiQcjUCS14rSkqCMTQ2j91tqXdIu8oIwHEajMVW6D7d
tquqvaMAH8ePmclTYnSJ2EYLf/RElqESxjUCfuJaUpzLjwuphepWk/W7Ybeonw84XD5afV1Bq/Af
Z3gXmOAOOfCcp2W+1xqfIsLE1dyeDHAqiWLI1oc8+Za4nm/2LxeJQUbKuxQoXQ/bX6aL3BlohJbK
7WxbTdw2dnp60hm0DXlyF3Vddo/fvLb5NsNZyrGQW/CI6Yeyovp7Zqf+JTyopvu/RgEqrQvkOlqP
o/PHyXHb/Xj/VfOzxZgz52QvodqM5E5+0MSeiB+ctQMoucSf6peUULa5pW6u2sVwQCk6Y/WkVZVy
bId+PHzj1ITAcYch6yRIgEw1lUPhMl6cXFMH89ZNpsLFMbvWJaj5LiBifSCXXgzJPownkgPdDto1
TxCaCAT5vLSepXxPmEOACTZByCJNrM3A1k5+AVAfjY3y+DKrQIVjs9lx+bR6GXN1CPqsMhs8rJhY
TaM3fW5nAwrcZVexfJblD/aELHDCQhb1vgmISR7EhnrjCiMeqNgw6+2Po6UtQ0OxaTblIJfCNMos
Nw3TOh7Xn+HyZL0b1LmjDUpr1K594S4M6bHBrfpU2MfShVHZWSXPMoFBRG3wA/eQrnzYD4jtEXMh
UV8pz+VT+ClEaxN658ppjiEGL8/5iNSsP95aQFWwVOYq5t79TRdwOqJUnFwYsiVY2DQY9diWAFb8
now5RabFluh4gRnOH0zJhXAB/P0W4HSIdFBE6swAioUKe0d2PjC0fzyUDG6Kp7UPebbc5wNOjeEz
P/Pe54uUwHXcJKL8QQBm8bAUylRgqGycMtJFGD6rTadigVz3hOB9wtGZZHBaSerocjQshOw3Ejiq
T6ZyNwjWWRgT8FjzsCicc+lLqUw4VefddzZcmXKtMbnKDsDwH+dbyzE34LEtyBy5773IkLM4i5Sv
EhzLSde2my6F/RqLnShCm9BcMqvzBH/woI8VhLhQTwFuxmxNJ82v2y1CGsZJ4vx+psN7rH4LLYBS
R4Q7I0TbriOcm0oB+FGN6zJPtaFEtItZrontNdAwrBEOEFRlCSov3osJQiTgHNtTQgN+04bPQ/Cw
Jiv2ECwV5pnn32Ah+yxoWkW27juBickrBs4V0/sWoDwWUEXeNfViDEdHV25R1JpdOqctwJmxrpVK
l2xP6pnFQOLy8izlLORRdtM6Zpiny2SWqd/aj0aWxfpE+ZrUAr4SUhYD0s5xEkO1Vhr2Xs4WUtDk
QU8NnYIBZ63sk5BsVYo67Gvi3PJuirWERo/bwBt0cBN0YksRF0avr7qb7zWfxHMSrSIqwWqBD0Gh
wZzGNt3+DlyqTdCSmaT0cuEcpZXkFMjkqRtaHP75F1pcGhs9/e9bh50oRMyDCx9bvbq6FXqHYdwf
vcLqJX/vkU9jkC2VVXLdlSb3SnRDb/XkCXumxXAGw95bHg7M2KEY2KSzayECCZ5YsYhBkDGi+hHb
FdxfvyHLVKEJm1YPkCMoY2ju5MeHfNpLCuMvbECl+h1LE7X0MX4nMTrR7Kmh/T+ij62oomSDTYFA
UjLnSj6gPsw7U7elROHJnAtwo5Prue/OBwi05SCb+qra0XeYSS+LR4ZZLCSP/65MqK7otvL2pouX
dIXHCFDi3T1S32IjdCtzrQGdypUrPSf558DngRiONRIjQcyxJNe81mrWS4wmoEyqApx1AujEm9Yf
DG2f3rPL9u6RrJtrWu6+8OGseYAUHerztojioR6YUhHKtLPLsUlu05GKtlG4L/KVbc+XPNwitDXH
wekwPS+txkREcX7wQLLsP56uerwis+wfAzd99Ai1Hz2IgWw/bhd0RHGiEBHLpevyr3F1CAmQXcSk
8JBw+hE/k9K6X6DZ3ZegsWHeHF8J9bLCFAMkrN1SonB3uFawhfuSRjb2NbE4K5ghDCFZx1ZYiTHG
th/ytH3BchJ3ChL6h/Cj7TJ6K3mSomtYtGZRmceoI7m26x5eyPHlBmCiL1K5LN/2C8e7W1XCcbQI
uC2nxVrKJpr0n5Qg4GvSR4AwDJD4DlfX2FhcMVjmLQHvSTERDLmSer+uvASnkfnIy+XsOv98yKBF
yISIEGVvMLNxkPJw3PuV5wV2q3gLeO6njqjU49DLA/8JvC3bkMB9ioHykw92epACghqWmlGqQtil
QtEm299hNi6NQZiVLs/Rh2FB6YSeDXdzGG5N92gWqNMQe6qVNkIrDzBZmP/A3EkGRm8Ab3NCPTp8
oXwVMkyBawQ3IlpY0lPjaAyQFKJ57/kBxPPcpBetymQFU+FIXN466ZSUt+Ob+HProkYIJNiBlCvE
njdbSyisEObXul6tEEq9xFpjCtxa+ep5nWuzmbYOAXJ5lVucPzWspRKZ0CwAVOQK0kk4fyovHKjI
GJNLJ+vN9SLLzRcgl1j13foIDWXiV7ZHQy47+OtH3EDRI3swxiSeSBQZFagrTTgiDaUHHTUgAELr
6j0E1Fw4ScicrWR4SYkJ1jJ681UF1gb5iFgYi8kQNghVFxz6hH/4CX1A+YPE4+J5mSdmmYJie7xQ
6xfrIHvyYlhxd6AWH+wuCWXi66G7k01e1oi6UCk5yQiKSviysKbiJxDbbCYnElHMnYJ3iT2GCa0I
6kHRHupZUKG17vvSD+DfP5bVZHRsnXHHnB0nD1B/qEkqN5DDoU7NaCaoBntFB5+gH/EYjVx1VmGZ
cEqmOA2lc8/C0zbdMgakYaBQqo0eZKVCWfbR0cU3e1lU6m0S+n3Y9rJCmKN7v7AUQD9ubJ7wWP2m
1pRJDKhZAJZai15+u+pXsqb6OZso7lhz2xGU1JlGhTM0hwHVWpyWaV2h34dlEOgLYe7QRMwlaJoa
MPycgPyRdqe1ZhG7f16pEOo270aGovAV7Ogf6ZXexPeXdy3QAe1lxzMgH1GN2EQOGX9maBNEaNbr
yzgrPpwMOb1RE/M+nu4RrQzRKR6IUn4N9otz6NIOOrboQBZu7m8HXPW4/aE7MqN8XO3/KcA58fTw
f1aPPLFvjOL7fHZaaRuSfF0rT/0LEs8AEK9qDCzjbcKa59WRWyqo2pmKjyLwIm/NqJ8PKWMeZW2v
VDeQTHk2vFZxNipkyPCoZNUYk32otn4hskry6ptaTCFM/fNWqOlez8ufb2Y55x1m7ucNbS1wwsfD
/ATuXoqTm5F/e5zCiTfWp8A6cVRZJgUdD7el22O9ElWUWbvLFq/UhuomaqHFb1Jt0rG3Co49qyc0
5oInSuXbjcQCZlS0FfQTvySRgh4+cu7RTOahDrM+sStuH/+hGQnUA5RN5n8dgyDsqc1rL18K9I5b
Ree/Yqgxy9Y425vEarneWp+QnDs/qxt5XOxss9+qGLht46m0DrnuTTRZglz8i8KqjYuyZ8alXWrT
iH9Sf3oV8cY5Y2SHvcXadD6FrxjGchYz3HeSQyVs+NRedvlH1yhSHa6BesBBVewifrPoXVsHuPur
5BHzmM5cuzZa6bZs8gy3OGs6eFVLfFUlCaqCO8ITOmG8WvJfHMjv239Jv14t7MIicJc1ulFqOdNC
cF1a6MtEcM059VDowZbs/vSVTJAcQZZwREJT/7J4xjXxJO/UqoBWI8QSBxdQrOm7CxaWJmsvlbCU
Az4C4k/gJZRrCn1I9uMrGwGnISxoZGn7fk+28bqOgPH4clhYu7gv5DtWTtnVEZ2zvqPuAKZMvNFZ
Gq7PLRPxxQuD/Id/XohXMRjjJMFdJtpy/HnF+wDVBflpPFsu38SWqh4pBaiD+p3nQ1CH/lH2GYlD
rPD9ZJ+mRRVH84x+mL0Vxfy3oWi4WqDojDUoQiutQCkDK+FfFTwqVAiNOIxHCC2Z4JY2gt5VxTKB
bGkRyUrQMe5A7J56GbyKZ3vRFqg3E2MYqw9ZFYBte29Y0/mq2ltB8ggash2/BgExSBAKY6vNW4mA
Hez8Oc4sbcdyf/Z7EHXyXHDYwQzFDGelr7UpWJrieU/hmZzY8p6C7BAW9yd2I58XEF/VWjzDWZr5
/vgc33DpzQcKtNPYta+FFBzT8Fcw9Jo0A3lojbyMC4OdenNEQb6bp6WMx6CxciLNu5S4oEl9dCIE
bcy7XvUJQLKgOwqzHlS2fjQIIBhuWIV7hCu/FS1qapRCy4UG1BraTUMUVS53gHutngn6ZhJjRWxg
pSyDW3rkWzG7m/NN4gL2bzDqiCAGwuAs6hVPj59tveX5I0ZrGbn9XQbnE51/wntc3tVWrLyCKa6B
/sgzsv+AFDu4lIX98U8DT1rTkSsGIbf4XYw9AcqRdWIoRqnSDg3Bsj7buHUdS7hWTSEuxAVxOf2d
Yu2gPYNF8mInENb58ATqrRvrXH724r75lU9Ym7x43X3OXkUHJZ0QJpIdASg3JILmOuIalBaSPG46
qer7IvPn0QRwpu1dcnPbHUlFfQwxO9j1e48Zu2BTTIunLbIHU1BonF4qYvJh/VqkJmHLAfMTEwcm
QcKf1rWymJZLkijvR5voYtR1oIJ/qEa6cBGLxuLO/R2biWV+aLm4yHvdiC5nVrTG7CJ97111mXYM
+nQSj11j1+tJ+NuP2rSPSMiQD/3CxN7ujUxXBiZRhtEFdE7GJDqJAXDp1FbZT3NXc9k5MRSvvupU
uKz/QIB1DXgkJC7Y0fevxXY6NjfosGIlVzzaOWa8WX6Dlq3HvcttBBiiciy8hFocyKbdVaIlmHQ1
UGmqRKSc73UEFtptS3QDMCsO35+h5HTMqpHwU9fLkkWIhqHqmMkHUkpE4z43hgYzJ4MjFsmitckO
LtUmMy2EaDZSaddl8vvuogzX+P1pstOS3RX91V6zOdl2xBnLj6oc1U7SRPqf3udEgcMqfUIUhdje
hZpJj9obRmbI5dj0Mk3DnHzo3aWoy6Jo4wi4R/KJVfEKz2BjWo44VFOsBT7uhSh8ZZzf5F8y/Xd4
aSyOecZVcBIqVrnyQ7LXqR9IUGpF7CWU/XFYhzJqRgZYdYP8UlldGrkyLgZvOX45S3Ub7bS6Mhkz
bM9JU1mlbCGH35I4YJOQ1YHA+nbArA70ullsTtudEGdO4CH6LnNbuCcourcPMvlL1UpPjP5vLPjj
ZP+QCoop82X8SBeYrGVVgAOkasMcRn84Q1QtHKQAPnpl32OQwAQjKyXadRoXfjjqB5yFNC+a0DiY
WgNpnak3BCXu1aB/WT+cMsxsPWoS7BDbCjqmADYwRtMHVgYj1Z1cQsgxL5q3VXJEYC0d4qLjf441
dXurNnp7hQremZ7+cCd4zhTf/zI6drqwF1geP6IgRsumIa2GO7vEU4cqQUCTf+E+efiQ/4pLOBXi
PScK++fcQF9V/omd0YTQ5nQLZQtF3kn6X4pNYNLCrbbpB2VpQOg6cGeuTe411wfVL8T3ubPC+pz5
W2Uaqn1pO1qsD/+lWcEv0B8l2YgxmCGM3CO1clbzBtYLVXsTZXJ+TfUgzlfs+QQ69rwIDnpZQe0u
50AHqhYOr6jeyrfRP+Mq9qk8S9SOCziPQs+/D+Ru6ia862Zft1qfT5bptmxQv9m6Eu9osUvY7XuI
J5zcTWwDtV/8pG5MLvnHoudowkGF4Rp7CPhE3RbEhcuHu/cPH+yKbbvndfFczdkmLiqqla/va1WF
kH8DAfUQQBGf5JnJOU24JDHbkQbvT0o3G46IWiwI4meJry1EMt7uv3/mz4SanHbU9GCQUZrrJ005
9DmcSweKyT4oTDsbCAoNSXAddR3/N3r7f72hVVnIv+4BMZJCNnKBcxwdCsDo2B5Bipvl2C+AHDwF
xT9L0BUkXY+wlHR0reKgnWvYqKpl1Az32kW4s5ipuC7QKXgyc4xn77plD/4lO8Jh5Dzzb05gTxlk
nLIJPipGpaq3mpoO0hGbh8kkPMBKnZYMEJvf2c6/l98hgr9A7SqYb6jckR5lDI3VOcaV+hSlgZAR
751w1V19FRwLQdAYxDEh/Z+ey0XENvjnwKDb3l9YSbvcU6pQcyF0rjxFZtmIClsCPmNWGX/q2Sdn
uyUostUOo8b2nivH7kunIHVRmOqLIIfIv17wHwzj+/qgMDdJH1K8LhVxFgWgIfWN9ndFLPK7dk8t
Q1tQdmqKrGWSROap0LkEijg1bfmPO2XTkNGBJw9ssT82gMmvDmSkfqdMIppllHp92COgjn3L2acG
xy6pewzopGUp7krOymKq6VN4M3xGqp43kSKg/oxTCKuMV2JCAsi7u7YHTXFy18SOP353pVFTRXbh
OZUahzk5zA0lh2hIbB+izs8zJf1o5gVmLRf5DRtHPY83OrJScIqqGsgmyZkt4t2buvWG+/8VNENP
C4tKmHdMkWj9F2sGxyQg6tKXnMkhbby76HX3sGYiRKP52tMNe1di/cT7vvOpu0dxIQmbZm3b6bIm
RdArYJVgHLvdUZaAf1WDYj4ZfCXykv/QUb8BB9gWSbbFYCK1ygtyUT3gB15rbacGjqQ3bOPWR3Eg
n+SR3Ve3iLzIR8lO/a5IVDeav4hwzeGrOB+6LAFPmtC6jqXIxPj5424PBG9/Pj7QAcs4G1EDq26M
KVi4386iS/WliOvT+VaJ1vaWxmB58TA9gGpJh+F0pSheXH445QNBcqIh22Qby+R7/prMhbhdqjhK
eQv9Za4mCV55t1CPFSJj9kDP1c9jIfrLNomWTEVHUH386G+5vJOLi75FQOosrcWTGSTgg8IdAKwl
hfUbU4anw+FHDC3be8ymhXrkkb54wBIUX4XmGO+om1Y534SKZU3pJQpzFAIeSyGEKVSyadD1M5Pc
Z5dwvHQpfwx6Qcfn0BpdfZwdr1q6lIvd79Osx1IzMAB+eEtkXfg+SLl/Xg1W2I40Il+o8adCj8rC
ntjdlO7BWxB08e6TPJo3/MpN5s/SrIUz3iE4RChVxw3vnZe6vQq9ZQ4xyKpEWlSSo/Z3SM36kiYB
aIHj3tTTWP+jDoqgE6BMB1YalCamSLFDSaMk/iLuyYWTEtUB/y2g6dmiwRnS1LkVQluIeCntn0Z+
6N/P1cvCA/GDPLx7WBU+uRUUVhzW4HDTsdH16mHA9WkDE0nKM9KJ7Q0qmsCgo0a+QeVXFego7io2
oF5h8fiib4yCClg5diXP90Idb5UuP4EWTSCMbTgA4TllnByuWZMX4wT/PY1H4+YvpM4WPJ/pRhLF
mszh4tQVhY859ck20xvxmoMD9hFgcFxZMDViXiqyUw0SIAQMAzyJlnvgT9kAHpvhCrVxZGZ+f6Ei
uDdf0E3cOOZTHHzzTgBcZOD9lNc1boSmWDkp2Y+C4BJkTstKzjQ46be3RqzDAw/TSQAGZf2pmYEm
b9FqYI7GUtWnA5K7iTiUMkAnFHqFb9sxuK1BEhnhobkc/l8fdJ0LHN3hp8PMyGUScGmIJPYhP9t5
GjTxqgnbKgGSdwNhyR2Z3PCyv3HbageL3Yq0zarDoiMonqMBDnPv6qmt1HpNZdCr4X75KW8PHypz
2wEPPv0I2naP5NCXD6FRFGOK5RhGTlbjFclMpsq52g5LurkDlD/GvHQzXvk3oD8MUYSlroM7Bs7d
DXQeO9xzkhexzYX0xZTAImJC+WxhUCt9bcOTVg/Y0D9kcK4/GiPtzqYt2zMUjz5lSeSxJtkOt04Z
RR+0IO83qT2/oY5MhvcxFDb5yVvw0cQDYjPFMpb/cmGEGyPVAzPW4/d/KPyXVC8V3Ebv+X4wSTR3
9XTBS4tsDPDzUWfPNa2ry9H1L64lacJ8R2qN5iCAgKuW1l6sNW1I2Lv+tTqcVUddswOzAsSdCguy
CoiAP/7XIU/lfA+bYefZ3FZCPFbiqmPjGxdfff2SOPTG0JKUkFUsJ1Owkab5q5HpRzxwS9Fig6tI
bZga+AAG3Kkk+uB5dyQsz0bFZ/wyhZ1oJqDMllBqXXd0kzOPLuLgFPKY/EuT+O6weRQy0sEiQs43
WIIOTjsym02uDK5saEfmzibdaRAlsaN5HGymIDoAAjd//jfLzcvWhnC2ZiAk1onA52qUYJlsS5YG
Qgx1mc43/NYHdRT4YuC/YvSmS/cHhjKalIjxMDmyRtmdck+ZNQOhYOCx85wR8jzzmeIxypJQDLZx
B8EP1yWk78oadO1Gv2INbrqlbavs28zvn9kndMT7kGLXVFxZVoFQ15wLRtBctosZeo90jTclSB8Z
guuGokodoFtJ/s5qk8/50+IkitBWhDc6MEKuxFXa7U86cIdxormWsq8qd2fB0WGI80mszhDL7MYt
gGQ82dj4Pi4fbrL0rSzckNlZP/dNWPfjd/eKNwrfm66abfhr1DXBUMyPaxhpxlOB8J7u3v8kH6ih
kNTHBIaI8OMvR4g/AW9M9QuvNLdxko73N/jhfjx86X9B8rNcKp0uGmVh50rYNUQFPQ+83bMnBpRa
rRNy/8ZR6Yt9znB9B7Ik/fgVmfZeTYnMEyEw5nUuTH2ORoAEDwX9Nz8Qd53drvtKIXWT4kaWDr/y
aX74XqwIZS25xSBF1A46YQBGmwlt1HSLjW+cC+TF9Y9or3ksDcyeiPs1p8ZZ3W4WW2XHlZhozBwH
ZlAO08CpXiPLyzxrre2ZsOlwk6Q6UP1Q+ExDXd8ADgaUfLUbVaPB5M5YEdRAEM+3mNsCztK+mnAM
wwa+FSsj0qOaf43K1DNGud/mKos4J2QGKjqc4FCVOAOfqYZ0xEHNuo9ph47U824uNuJvexSYqCMG
imGd8xbxHpwJq2zMxwJPVYTq9ukKp7Mmq9bQOovsnvQzMFReAnPW68HfH47xfIJzBNBX/w9h+R5W
oSMHNYoNkrQvfSogGSTEYDPhNVe16xQ7pHIFNLjFER1SRB1pfAO75IWSE6ghivm/P3uCctnYZhG7
J+W9Dc685rSXY1RcDTHgFZ4W/8T1IsTMBX4NJDXv5Yzmi+LYGtogsxx9Mnha9vKAZ585WTI9zEnY
K6kJQrLHXl+cWeqzHX5r6ar9pO2K9mtKOmCyHV85tEwI6ULGd5FBGiHrI6E6Kfw4snJ3R0Y66CK4
Vp8z6wVmZTZ2NS58alWVNe/E7G81hR1kYm8iDjT32fypyPWUkCXwtjYuY7HG8/tUy8S97kxEdvQ7
52tuqh+d1VP/ik+hNRGT2oySqGfWhI1MGRynGT8IGklLah4zKR4/Bab91j9/pWdbgbm1GaLdJVHz
vvyOpecqs1HJtmxaWfjxuTEHpqg5+fUbpcYmLmK8dc33vaBrDzfuHRjgBiCSYMS8xyPKSUP44LZS
03nVil6MBGSFcK9x0bNb1xBkUMqbnZvlWgdgCL6+FXeuLbfVClimAiLkN84RE2txYIHRns2Jmf8X
puGoBMKJ4bZ3ji1+mtaFLrDJYkzhCExfgG2R3HlPl49AOlzrhRMupXcP5//oR0glQ3Uy+XYBRQrt
xqebRIcsSWN5izW6pIWQI1b0HSG734ZieNtOzAagfiqsKkt7CCPfKbm/YrH9crslAKux1gAfwzEg
B1/AUbB+sy4Xjm2bs8ja/Iow6weqAG5iVaiAiDqt9as9MwBzjOyP9B2G/hjxjwxZOGCwDosh9vmo
2VAxQ4zIpxJE/GsreOCeDdZFQZKOhgffY13iqOp0WGC/aFOQAvqM0CTZ1jLy8GzvT6nRU6WKRwz5
SeuvXyUuyIs75nsSPJxHctqDcpRYRJcy78ac94neJAigmX8RoDPhPC9HmE8T3Nu22oXLbmCdcjuZ
5WSW8XPvjff+q4baY0jRHfq/vg3uoj7wGjEdPtD+e1afuFWRsSMbTzVNGI2J514OdGV42NGi1Qa4
jgaJjA4nuxPTrJWR/fpoXsdIVCjqNmW7vu0H3rtSi4SQ8N/SXiSZXtp12TWkUOYkfdx/8OAQctXY
6XcYXpA6694G5K1E3xovhdzhqLOV6SbQ7wEr+QiCK0/E3MCbxUoJteHCVSI3jKHML85CUUR7IgfF
FRnZ1vZV+4miuibx+QVvY+CZFgzLIOe4yuv4DBtGNnAf9VGQODtlsRGwva8xYqrJKnH9x0hc8Ibm
KMOGnAF8EeiJPPZVqjmkXlB5NvJ+wf3QcSkcxbgqseWBB/EIjRi6fknjFmPeRIsaLWGVo97/QDpf
ztM39BXv4wXD/6rVzaZEz2+eg62/nvU7/a9fKbw4WcaG//AmhW9fRLg6wvtOYx2Z4HS7e7y5zQ/w
zCvcbQgygDDqVop8nMc1kpZCefy69xMwIK+3v1bd9tRhwZPXWUuymF+1sSbAvNGmheZCH/n/R4fN
m8tIZdAd/aehTforr22FqPYOcK758c2C3ffX6CWnMKMdbGvYYZAz0ode505/ACv2k/jDMaETHlq7
Cpy+91hYt87y6KCIrUzX4xJ6zWtZC/qxsdIIV2i14/jiC7f+tdW7N1p8elaBBO126JzuhNuPvbHH
tm5r+cG2TooHSH5ek/87WbxldclterNodwyOpLx/5ZUVE5sxRJW7sZAw04pHQanixsiel9mSOBWQ
JT1hlOKuhoJ2UIkGCY/fW1VlGX8XrV2vbQvA7JK1ENmbTghmXwR/1wK7LW9wETaHTIAIC3k9m4mM
qLAr65yWkrTYTb8yM16vH9TH8HzdEe+RECpvPU3NCWOwOv5E8evwGIkOSnMnr0h8xVa+KSuObPD5
JkfHSVMWUJIwvGShTwgRqMPexqT+u9St6i0P+Ts+NUoTdeWDOvJsNfAbkkNxHaV5JmhhSb5kaZAM
qPbL+EesSLDBEDEDxDTPl8KArhmk9ioEmoMnre9M92x/mnWOrXcKjAdtFBMi03aGfm0j79tLFwDA
Y+KQ/PSScuGMdyg1DOcByX+N2IjmDLfEMUgoejt6YG8HA9ITUVTh2OhueW1g9RLGpZ2Mnk2gPgMb
2fgxUIrMii0lmEiNR/Y5h72o2WbpMgd0mV+N84hw9wER9yYjSzGmH7RTqGbJY32+F2upFE4bmNX2
voeBrDxu8fdvjZNtPkTuX0VBYCY89LJKRBkbNy0gU7pghESjflC0k9xYk+2TYcLnT10Jq4Y4ve8B
i9gqXeygSmzhlU3gqd6NMSCteJJQ4Dud8OnHx4cULpNI5WP0u13YQkp4d9GxSRj3ViJowF6R/mJq
8iqY3pBfxB3slGKbi83fMSAipqAG0PkQVmn5EZcS0or1YF2gCSbJW2Bbkj0F1/FYViI49mk2wG9T
QEzwahDAnUJ+BqyrWf96EP+GbBPKU7w6N9pN0Bv/SZX++v1TpJUZcdTU07p0Pfg61LN0Krg6OEkj
ASn5PKpqE/8w7TURb2O5xQjU7FPNObVzkOBxETtVwT7Xb8DBl6KoGrD2qc1PfYx/8FsTyVXTlQUM
cG2HxIMHVfCC8LufghBEuwK2WUbw/k1PAO/dmVHPJWD/Ee8PZNEagAyAm1JsAy3P4zfkDdGLRRZH
xvKAfRV9i4Ay0vDK8N7Ji0b/BbjvdxnuPZuneWoag+AO5A0f9UjA9I89lmCbrYJEF0wdrs1oQH0S
5BndNoNICqAlN/bCYtq9QAWTWfgygbkNgzjO2Dhk+CNt3cqU/VOtymI7jOF7KqwgaxIoAQJLgk4w
k7NEemab8D2l8+xEwA3wvEFiHTOAfzgUf15sHNDZccm4uWsuW1iSMFR3XDLBTPWzHVES8kn9HwXD
IoNqNP9FqSg4TscXkdtyBLjG4rbj1wl5ID3+WCwOmCUA2KsU4wdvmIE3mSlDStFkyuYTnLx3AbjJ
53ORiiZSjVNk1jUuAM8KEESQsy7JTt3kqYGMyT2bCeT9zb6z49sq7o4poBWUJqs2vLFj88BtVt1W
QLIw9Lt8dKmI2Z8LoEqXSK/FDMxlNYdteeBRVFf8zreGZBXUvOhh3ntL0MX1PI/rKgHqZVJXMlKq
bER4bsIiXIUxvIz40gPmcom4ENr9vYV99n4LYAEgFOB5drvCfUnlC5CIfyXhj68PrnvoYLdZGX6+
+yA8sKN1wODkbYIbch6p+UTfs/pT22wLqr5aat1sxyLc2gZ08JCDoaRme91WC7ONyXE3olo7BoqM
vHjtvRUzcG/aGPRFJ76bcPQG9NoqIeaxd5q4KBI3kDuKKMHYb4SNpOfv+Lo+J+Ub9wqEhfLnCJQq
htVVjFKkBgiRxxED9ZurK6GOVpILYGMvDIFHO7x9+xSMyieME2sM0TrIiNCitz1BeKeu8GSy7lgh
UJWcs7+2Iw3cvBMUku/QEksdyjHCwzsCsmKKJYfQXc3Ila60C8Oy82wxVDpwQFSUirD35/1Tehah
Uz0Z+FYZ+swnh0q4wKdDHi30ZUZ31VYs+Mr+12Ckac6t+NlynvKvpj1V2YP17gmww1WPUILPoLm6
UFkbsd1gfGgbKYQiNUZK7j2N0aPC0qfRyoYApXGBYhuhmw7/BDdyIbfpmXeOi9sN4QmbOz3malmS
xqJt/AB7MAmmAZ01CgOgumwaBIPQf4ROlx0w50pkWh+7Ah7ajfOzJ6EnK0JyHLgND7/9JPs4DGSE
YzcxpbJzylnKoEl68H00Qh/KbmHlphrHNM9Ec+/tJtqvTwU9pMJS3uGA6gyeZ8DyG8gPRcjGCM7r
xr9Ri2wSHK1r0FYcfCjOZZAlZ/Mb2d1QVCK5CtMG32Bq7bnbqmjf8KPZmEK8SqQVrd4E95dwATIy
3TDxpoRQNroQ7/WBi1tthBpft4bYJ3/Yadh0qFhnhcCJewEge2cjJWR8atuFKrWbg355Tt1lhAXi
Oh5vsh+H49vU3nnYoxsphaftjTtIT85+B4Vogr+wu7KNeFMeeM70F6zuaS6LJPnj7Gkg1LhsUsU4
gydMNpAQc5VE8CLQBnG7PX2bVA/Me8Se276p278MbznwWKyLdmmsequH0wNizP5qHQ5UhHeJKLPo
DE0+wB7nizMtOmpX/ED4BagJVK13bYE5SK3xt73pf7a9tqeI+Z5o7xXymD2/Q5X2T/fvbA5KuKEs
MnZCzc07Q19EdZaNWy7WXlowuE6zT67EbmUKX49yC4zs+JTvC8Y4jFG398tYThRYypNAGH77qv2F
d4TW+2E+pwAF33tzmSWM808yS7y1UfN/EfV0YI28Vhbdm8gzr5vwfmBHuQ+3pHcXbCFKYoCuU0Ps
QwmWHSd2hRlZsDKLstWQvbsGLLJp7IXTjW+2o8UhGLcBkIRWDxqnnVGZGYHT4quJQubw40bR1M0O
NFI2AZk95w4CiYWgRJJcq03EBM5xyWSQZKUnwls9NCCpW0zPxQIqT/pvIkME+RLH1E0VRnWAEnhR
HSvwDexJ7RVVmz2gtu2GwtBgnhh0dC9xtwdMO7SKBtDilsYzbN0kU0vh6ODGabWx/zfyAxoQfL9o
tRupbYg4XeT2+qSLNWjFX3/TavplzYyJQkzaKNJf+Y1KePcHCRUKCkvhMvS5cjONF5AYPycLg+73
lrZtBg22wnIwreYzLAfAeyf2DzFbwyinIhjmw3iPS9NHl6TsVuoMou2KCtz+VB/MwZmt7Rr9dROI
y7oWpB04yPhtX7m1lmqu2s3rgqB/2WCTSESBkBzCJ++zq6e7DE0KmjGLhO5ncTZBbqKDpgxeH4nY
S8HV7e6OBoshKYazFDHJouKEX6DztzOvN1lSiJxA7jbdop4JuVniXHkjVEw9IUGhjiJ4Y3gPMRRP
AehNTBvh1suxoHdjsxKsbnuLToNS20UaY/bEBYOmOm/A1sTDVtagAhAzgfCRMVBpmWxSW6OwOGMV
j4jT5l+nMK2SOPe+UX4pppN9xlbvQGtMLkulLd7Xd+YTQ2I7sdocmB9jBUAB7roDfd/CIFXWQus3
Xn7CL7GbDlWMn2FeV9WkQQc+4FvWX64+CcQCVpvXVkaOMaWVzT3BXlEccDVogHBIm9wH0QoKz07l
eMEENQhmpAOXvBTr2yT4nT8zPhJqW9SjSPplpmT7f3xnzlMsFZracaEY/ZDzUs99LlPDsPFh56iw
1GI2SRNv+2k/NCKscspD6Q53lnak9I3lpd69G3xKOkI9pKVYi56H1iuEGVlyxuqR6q6h2m4SfJs6
lItuQd2XE9TyyBTMdO0pGBI8zHn6mp20MNOKt+CH9ShvTrdNzmUfcJjJM8BkDlwzBSPUafvSJ4B1
0a9Up1TgbjBp2QIV6/M3vuRRWK/add5WyOXqtlnmhrvmwevzdoMki6An0eQSAiuTb+GfP807S4PV
vNnjIptt+TlOZsvSmGdXPWZWiyQEDBMWmJinlM8KegZqG1TxMU49YdOd/uIpIUOuBzjwHdzEYmuD
Fszq3pFumQBocsIgH/Svj+TbZ5+xYoJz0wf1SbvBuvlYZqo5VlzR8DzcFay0jjogNBzecheyQFkJ
R+29ZxcZJwIMsTSJ4X9NZaqQQuu1hbcZZwTjhCnMa3K3+RmElXxeFDE6/uxfW1+z/4l556mfqAJX
81AhzUuk6upezz/jUHCOaz2bEdNTIO95ZJT6nEGvKL+besS96+/i4Jawr+PaGPtF2155UDoYvDh+
wnGx1/xgfn1aANmTHpia6BZV/Pa2cA0LM4dbGcgfW9yzpRbPZtJf0Na0ziCeKhgMQS4H8JbN5BOp
rPCAXCzSaomr4upVDCPQ5Aw9bFlHa5Um86iA/fjl8dWwmLELdDpqfP+CTsYh5sBsQjcLeNfsBOtP
KyaCuvKp3E9NAXglbCYJFH7vgkfcMPm0Rr5z49LHj/AmckCN2GktQNurGlGSXLCZeDwlPVBdq1Gl
FFvHjdJDLKTXMkzH/CIQAeqxXfS2A+mXFX5WFfj3yT/va+cOVQ4B7nExSMvDC5jXowUo1eFZbC7k
vsAtsvya+QLCMFGFh91mGgVYfjANIc66tH2NkiEwhMDCpDP6qyi2rxc6vuCj1zpTl/Zkn9bk2e/D
cCpQMIicnUpStc2RhptCmfqPuQpzDzHJ1RTRFDawxgSMQXj4uT4yQHm6z96B9DMcYghPRFATNF1Y
XZs/DqTqx2CQyL+Bu2JZEhOmhov1+F4pU8zbIVYaQUWgRy4z95+kVMdTCPD29HmYUICNtPQ+QoNn
JU6wLcygZs8/Ab/IIWPE0e4+reBeq27au4pabnqaimuliOpsO/7jIwZKAIkOYhvPidfd/EqioYTR
8aXTjTbDZ+Mtecl5GvxZlaSo9QQZwDW+pUuGzNFv+jIh8eSLEm7Fls4O3Lbr5L090edTzCr6WQa6
1aSXDRU9uETp6Tjoic/CCnrD3qCJijC3sGliJnWIvWuxZBwf/T4qQJaXJJ5Tc05JS0x/rHk5D2ba
yB5SpPjvNgDkrYl46ul+PUzHbLgHBcKftYQD2P0ldNJnUm7v48CY+EG9EY//DKc7himK0XZnbt6c
qG+NPEEIhRz6+tKXndXdZwwgVnBRSpml6BI5jckwEIRnNbOUb44AfES07u763D+jzoBX6AK4YOM4
efQHyrqClx+/A9hAAAPvX8/SVSOxqane91cFWGYdbXqaLpxe09pudsASHMgXfLxqSXECHzKosGIn
X+sSsKubZBJc88K3/TBZAcDLAzOAHBbSjxVowKvbzwEEjFR/u7PuSwLAsRdQ9BdKj9bVQgq7Ghyi
P7tGb4iv6SFyFEUTmJvDatgzG3gPrsg8Rtu5lITQXimCkYaBtGfv6uOU/0iCaFnwtMDBkOuJUAim
Zgz3EY7aNJzFbdXt0glNyCpUWDqEn54caSd3ijgqxIwxEvHAlLbgxAdbUCEwaf7RAa7aw6hON2pF
74zCj5qZcCwolN4fr151Ca2pgHiKb32iDqA1YTSmE/Yxr8h27twy2fulXZzN2lFh3wFLK7kIMl31
IaynDhvv2VHmgtRfOrY2PVBIF2L+zwZp8d0qdFfnV4AZ9/4YNyFp24p3uwTy82Kz3u8c36EF02jt
PCc6Cnt85oSU/tqOpMUXWSDZ0I0fhLhyihLNXV6Uvds8TtKKmmfF6ioiDPbpwv3v61eUHC1H/5oO
A/0J98zvY6g3Awwq2mdmCxUJBGMkeiinpLRdBUJ4muUBP86+STUnuwFLAI/aiaXEuqN4wKpeg3Sh
VqJY+kQiilscinE/RA8oIImsFIFNN+RsUfSVjVD6ZZlKd4uinc47Gpm4bfMQ6N6VB+t61g4jgwUO
p31Ed/NzC5YZA70x9VUqqssax3NRvnSq7+yV7l4cq9mzkBOQ3MFyGry3qITqZR0VamCnSos+fx+N
mXyDqiG33wtFMZ4iYDclkLOkrjP8JChwGL0YYygCkmJCtMtcZ1NJIz+UGBnVWljupbxLHpywRxma
alI/j9DsDBlp/mIURn+u2m66II+K4K2Xo7zpTfqXVKMK3cGPk+UI90H4XPeeZZ2ESbhyWB9e5MQZ
7xRPM60QEQuPr8I0NT6hr0AIM7ZfkYv/7k9XTnYMj0rIg9rpMfWg5snJxDHNG0sjmLuFXdVN4mtd
IIuaoer8PLd+iAwaXmKBWUYoeTSH+yVV1XghZKulUWiexYAnXjbo/UAvDk0PNwmwPJwcj6aibR8p
iIz/stkxPiVOP9WLv6+lqQ7jDhms4LY/EcHMU9BQy15YKIjjQgsRvWgAflhakQQBqOeQfa6rkBMB
3vnMVIW6lQ8VBQv/dDa4AEXo8h7IuDtSmRYmZQHu3jUFgtllxfLtIBA2PrVcWivv9cO4N2kn6bd2
Y7PXhdaNdQPTbwqy8kb3mOVOthb2T3I7zpurNYQeZHhs1dB6CF8zzdH4Jw4lzaNBOJmPx2TdYNTg
3i4FJAJxI3TYAmhRmlQciAT+O3UQIQHUEJAa85O64TXt8CvQS6fO39EeXgnrL6m7u2U25DQlx/NN
lXjaXPvPWdmr7SkALiHy8W5lPd0tGB7ZEEl1uYnpnRlRZ/7H8283BOyap4wEgHdK+4f+L2nCpQBP
LqIr5sw23ToPmLh8JENVIqoAnlnd5t9PAIyy+BCT9k32Tr/O5yL7ayAasBELvv8+2AZngX48JQ7n
JZt6pVTDTqU7hqKvOmj1bsJ7R9sPcjU77BmwIqI5TtoxkL4BI56lUBJHETIGTNTHYrOZlnam0oHj
tv9j3KGVF5yWFYirq6TXH/8LSCbBREcDUMThrnYXq9/X2TKEBTN1oiLFdZabCftUnilrs2exs8p+
cFJBRtq5aZ3fcVzmd15I0TvL+p0F7YcKNGdolT+rwrBgFG3hOO5mRHOSaeDcU+8WqDAdxblY2M3O
I69duE/xnh5Kwq1zDQuGTH+ryLF+meALMLc8PjzB8Kz0Z2PJ4Mjv3grrpREgAU3XqiGzhQJ3BA9u
OQfE52yE/LUu8MVNWFvO3tX99Vw3JvK0++xMhYSuvcZldgvCjdnRTE/abCniRh3YVpdSuL2TTGtl
4wL99K8Z6OQJ8jZ/YlEMmLPtVZJbaiHV7k/0YUpHQ5VzFvBN0mRS4ae4jGdz4z+N7NI5eZKLsgYX
2V68Hieffo1zTZJNVWP39VguVGVKSIwCChUHnoSss/+7WT8NSp/R7U3gvN4GF2SiIfvaViFbbJm6
3HyVIJBHgumbI1luWUB+2Gz2TwZSqIHRyLbi8/hhFm8/s46GevZ3kpBBUCIR+tkzx/UcB+cd6L+e
b5g4ukiAGgbsfF/VRx3o8b+r8KARxDkPc3wfozvhjlWarl+59vVqm/0cUauwjaa0yDDMDshyaZu0
yEiDN4qDtXHRnC6tkz2csf7mE0lyoehGLrmz4dpK/2KMXFDhlXktq82PhLvEfcJSfxjLkSBgwq5K
zXahuJgK16EwX5IeN66RElV/hLqgT3VN57WjoUS73r3wMoPpaeqjAlosAjPFXZhnClbrMaTVoL+D
Y4WRO37uXwc3DR0SNQwcMQ6oeWq8P5z4q07aA6vENyfdwu2+U0pH/VfTqwLtheldhnRWe1R4yADg
CknepqZn1x0uc0XZt44vP7FdtJ24+yhswN4wuz3nZVUuO9A0hhr36oXiW3BfM9MjvrGPQdF7s0sL
Vw+0a+MUIiuPzksuDBdX8b8olhVCmDzFKfcqKD0LAaO3GoEMF84YDSOLh5FyIMh98fD+/7ipV1QQ
jRrmjpiGk3FKhuI3HSTMik89e0GSV+0rDqAxYHBCiRGDalGDMrIUEIBOvMPcfONY08jRPnzsnlT6
gLH9aY6bZLL7Vrjm/QzcG32FSzC5oLEu0dh/Vv5YQtEmLcsMe7fXzTyjqzA17rBkMDKjGF3uF/bN
Rk160RC8Vi3RBCOPLptkQuPJEuRn5D7hOmVU+CibQQlHxB0r7H0BGGJ30EOLrUmLVT5xPvT+ZPeX
Jza4wb2xcSUjzm2UEsiDMSX+UInGSEtSkf7bcx925H/A+RaviwNPEAJ2br8Zo4XuK6PE0b4vmVOk
sHma9tlm3dIi0mfxtyExt/9EpPO9BMmrlMjFT774DXd/2wWduW0DTbAJnBQqrDUgzaxqjMEczC/G
yw7tI2oJQLz0d03DS0Pt+Yf/1XDHuQa5guuHx0ZHJRCne5rerbBWHsApQtvrmDSqR9LVmvCFFO7p
goaTr5IPXB5CjtfmQZov31Zjq29ldlD64AcSwV32f7gJQb4+3tARIsIpKfCX7HVWpy35db5jL9MQ
3+SKlAgmcyvCW+X7Hx/8HIQDUKlQJZOaVJjaynfERUYfsmQ31qUNqc8pmJUARJk7lm3eGxlw0rl2
aatS3FEgU0wgJM2Eb12REOXJ5/eVN/rptfLDd9tpQRh4jv5sArcuen69e0Kxap+WOq3/q/KpD/Vc
JnSbYyhTcrqRfefqbzmfr2Ct+q7m2Z5zwg4ax8+a/gmbf+GJbzXSZJHAbMkpUNy1ibVctND4ih7y
PxBj8NCKEdqQmJeXR/W4vhAnRoywRxGuYAIva4hbQINi8ho2WHLgBD2/o6izPpxmkkL4+rFG7XzA
X6O175fGNa7T/4YCb07Tg7ojbtAvorCxC+XClfzyUKqphCFfjnhM+i7Cb6SIhjlpMFyS3SK8OJ1R
+rOfvqpOMQrEpVtqw5hox0X4ojA8aI/t6BCVXeUXxhMBrHppXTasM8acpmt/q5hXLhdR5kc1xvXN
WAQNwY+ZbVS6M2+82Eg3P6qDvcSlNIlEfZnXJ0OfSlsv2vDsjQsPPK+D0OtPyNEqEsN+JZ2keL6n
sq+ggqezOJZ/hp8ZTfKLIPEIiAf8dvwwlgD6M2wsTlSrx2s/cQZBqh5GyMWiigwiLGM3mFQikQrB
iYF/RIX2vZW7dW1BwYU2lZEG50am8ngltwUbQIjfhWsFQQCe0XZW/mimww5Wpvgl8IUr1m07RVpw
qXUFf7FDQRHvM5/Q+R5+bNr8sPOsEYVfXiNC0rH2+xOeUBoyWzrwRqRjPaIhq+4McHPHOF7FPzaO
ssbMr1AKAtx8QlJNaKOpN+FpD986E8JFVOlhJ0juiiEngxRgqK+tOHekNIVZL9wHXU3bKc9zxt3F
qT9oOOej5fHBGG7kqwpY1degnf8XVROrakzCYIV5Ul3QsZlWmr6w0as5sNQlcJVUglT4JV5mQIFS
Ti7GXIjqcUo8lAt1kA5Xfx2yu74UGE6cIQBDvnB5BgMiyI7GWkPcZ5GuU0YoQj8Uv585QjxflYXi
yi7qdJzhjMgd+/kzWmqBEQeUuOy8MbRThexpCb4C8LKYC6tw9kaTPBIyAO4lC16rOxVxoyr2E292
8xhi+mHF/cR7AFW90xevc4TIVnR00DYXR30z7Wjv5aY/aBePumxIEjMBg+Ecl2xpAgDcs5ENSNwJ
TaCi9hxdnLhFi2ByUQeIHXwmrJndi0a7hXrASOqy+t7WUNSkSnzddm1PxCSQB+zf7Hocdg3as3lY
RA36HdS8ulGc194d4UL4NvLc23pzVaQneFIdDriPaeCPBUf7s7fDd/Rkl+zrglD0wWfN63BOZKu7
BqpvbKnAoPmTAWtk77w9DGcF9QTF/ITUg1M1yiVKl8pVaXtE+dMx9+2WtEQY+Fu2oRzJOV+hnv2b
17O6PipybOoIOIkQzIu2WLJJhU1i/jYkU1mOfP+Qt15xbCZx969JMSYlukClRWqoxDKmgFN3cuPZ
Y9ir7c3OwL4UovKVWHzENeZ80VK2YRMzPqwN4PHKfJszrSiCSGK8JVmzWfjiW4jeFiHEW06EZM/z
SjiyW37B5HNSrm5gqyINsujZssL7UgrmjZQtJTzF+m5DURa9KQSph18S+YinIKqAcHJKv4tn4Djs
5PQhfJxYvVXMYrZmLjjFSkAwq/xft9aWAVG0KvuQww4PDH+aR7MRjEBaJeQdwJoOq2T2Sv9Y5zZc
bH1QlbSPUOD/w8FmX1Znylf3x4KTTEeyC15gpq092L5cWC59saFZbkgPSnBTzDl3aC4bHw0tn4cz
lWMJaO4MWhUev7+zNbD8TBJmkYAnjWXoSsKTNFmm/9ai7VONO8FEyk0B3aDeEVOmRm7vOurxvd2G
wu5CHYor9E0rnkXtAVnMzfSB6AE1ARx90oe6EP7QR49EVmr8/UX3PATYroQq4q6RnQ0Dy3wxjwAA
kpWjWQwgWM4NFFfaJsVRs9eUMmAjLl8HE4/r/DQW9WYk3OsDo++idFj69U+F0fWozRcXDK6OBfOY
n0B0IRrsiqQ2HvYZnJwLZ16afsZB+tNL1UG2LlBAiY85F/NsX9h24El5/VSM0a/aPo+/+9fUVyei
vVPOQD21FEZ2chRH/Ga56eV/JBNuBFMRMhWk66wETd0L38rG26nEyBAGcPDvk36N6H+pmSnLfk1T
8N2fG47D0yj4b6Tb19500Qt1ly5FMuL/buZ9exutcVJl3ckthCcL92bc8x2ObKn3h278cZvR5i3f
stPPUkDI3X0PpK92Avu5bXjX4XXZCGvBR9T6S9pbwo8Ee8DwZ28Fg7yrS5SdFmfmWr2ewG/hdMS/
ngzEGpZBrmNS9P0LgIfzshUy+Jnrz64baKEHepPD6G+O/X7j7GW9PQMfGTBWlXpRqCHumHi1shN1
8eMC3+qJBrlNwq9J616tKrkroK218pbLkzAalEQjBeXD5XoN2qU/U/O1De2MWhnnWtLc9QuB1/bA
PQ5PZ48lHzwJgdoiB0wlpdfIAj5GN16LqIO9gJNYiat0x6cF0Zr9HSRKBX/8uTqFkYDxSsbWlrnw
4vUB/Akd2nMzRnNcdeLZPCaZ1XjBSwGyVt2p2v8Wo0S3wjbi6m+wzjh0V1RImLD0LpfckbakFE//
ZQbePGUsZcNKSuF+D4dpdiMCJxjumRZemQcRWPnhGyl9yawkW7/O6ixj6BCCTjMNno0TqjsSln3O
NaT4F/2+hTYVBGDg+M3Mr/Gbow029Rwv+nSyxl2oSk+kdUz6TVdKfGAFnBI/LqeWTUmQhi59jlFw
NszITQUGn0dGAqISjFR5gm3tj+JGUEnMPUfsHsiTSL0AYRyW7WGjgwD+ldqD3f91ZlL4P3/X34lX
L3T5LX+BnZcl84T/jEiam8o13Xkyqk/oT1Qgt9MJrxZJTj0KYutarAfsLnsn/7BO643q0SVZnn1R
2FBD4EANM4mkI8vtkLPTFLPKsgujqt+eNlMQ/O+Tt0kX+dAPrIQJSmE5Nt9G3KeKOn1WOtosGEKP
Rt2VXYGe11Zwvh/hkSbQmqrDb7E6Q0BU5O+8khlNc2eRdl8oOqGnGQFS7lyUqTd276JrqMPS3vbp
/3cIpWf30gwWe2Y6Bcc9V8QLc9zfzVMSdg3Jsy8AiY0wPDx7g8pFOQjS/AvGvehApmHGPfYI7ITV
zbNy6iZPqsBtvnXQCLT97h382BCmqvPQBTGhwgESPhoRP7MksyqIog/6jLvUlJMS/wzVPU7s6sgl
6BuH6l3pBKQdFJhaTsTZy9O0O4lk3MJq2vK9+uAKgFQzFOnWvxPQddCdAF1L1PHkwcsemkOgzh5H
3KV6AJcTs+UrdhIXJca3NFnG624eMe6F4a/t+hbGqcNfdojaGO+24ZcIBqBGgHwOoh+x/Ih60OYV
IxuOrvALzQzCjr91f3LQ7iuBMUGBYpy6RKVhapgMTcw6ZMmvgMSndA/bYmJ8RovCLSrfpZTWZ2Pc
RHsDCLI7Oemx5ggnrMhWhl6n8k1+17XYQx97kC1vKNYWYpUUZ14b2Rs5DQL1senEimmuv42weJID
pMFdhBnrEO3pwIfKdu+eizbMPtJONdGUKdnIarjyMDbTakJtp2gy4bmYz0tGPoZoj3PejkBbMSdV
qTasEPL8tJfJz8qRHSkHBCdPBxLwaH0kXuLE/99nOxiTm3rl4wa4mRoeYZI2/QrNqk9KG1cKI7bH
Sh2cUWz2LYxWehDWuBvwIC8It5izz7jbVf/9Ask3lLkh3Yh3RFYMfn8Z6Mdi96b9EH65Jvya893m
sSwJ9gVdkWtq9NO0AfLKqT/MTCkNkp1FglggZ5EFXa+meZHmNLCGKp8szoTldpCs07VVwIvfaxfT
hDothiVbxsEvdMl8JmzkcZBn5VZO4cTM9TboKPdoMnyy7LVe2czB/tQhuIl354lGfT1i/F4xac+F
CIZvusZIih2D5RTmh6HPs+K4aY0cw2xbWPmqVf0cyiTmbOWXcQoFJ+aFl32FcGJHcqfJrpUxFc5W
Dqv+s/V4Uj2lU056AkfNB/vETAjjtg7WlTV5nr2tHir3ziypnqHyGNFHh3BJNEavU7bvcRC9VzYJ
Uo1ZNnae7i/RgbFwhEL3ob5/p0PLoDsJ96XztdB2CTodv1OpFw5vMeFqjkrcqjbqTGFXZIhCZ40Z
7fJ3vuaf0/ZT40/i8OOiDHXJStXUn+3RmT4V0oVqUYsTp3OLcK++946CzTwf0q4emxE7XBYQNPhy
GhFwCr0qTn6vqRGIh8Y89cIE0veN/9MId64AKI2NrlA08zTfEJgkZRwiYiW8D1/R9Qd0OKgZOFuA
1I5dr1hjnhN1f+JR7mX9zjhxPF91UmyIaeAnqLcOjdiCmspm4c1xUGpQevWehBsN0GYGeISJ9FVw
P1YAqM+0tFdon2W7fXOMUWlM7xY7n1oM1B/CaQd0swTcbzngjKTlgImYXwU/o6lkcB7xkHiOgw/C
LxMQJVK1QFMmetvG1iKMwInYvRGivncWpgU6Kqbdf8Fc0kTxTZkPuzPVl11PSKH4WfqvuFJ0Wkn9
WjtpUL9R+mMcgNY4ZeyzzkawqDb1Iz4z781AlpakKwuYpKE3KPAO1XU9FUvpmQmJRVCSdkBNLfIo
I9nGtsjzHZjmvCvcdeJly0VmBnbFqvgG+ooI7eTnVPeaWcsYc/YLAFBRVsJz6uYSiZ85mL1jcq5b
idQL7f0lobSytRf9gaQCQVOUQhGj0590kTj4GNaKiHBQSKai3jWPROJGCTRUutnHMMv5ZaRd7YZR
4kFhhs3rnKzX3mkjAFgdrwDfGgPm5bruVf8YMrblhr6eQrGINUlDTQX0/8erJI3b41y/bOG5qIXE
OH2eDaXxOujyHhsnoDrVMNxG+7RVowuU2aLsa2Ktk7zVM0VO2ROsxowBsX9PkppD8BpQwQc0Y0oq
GllMx8efoipqkM8/0rwb5QKQm9/0+hvcMfd43iPg5RFmODwXtVs2zdz6sv7wlaVJ26eLzDNa3sCI
gVso4X/XuZUQW2izac15CnikIfFqn9lUkSxzQJ4YEc/nib+A1Y+JOjFJgK/o2wa38ZwUkLa3MH4o
E64OrDowafF2TfEDl02A6+V1RH3UuMbhMVV8ifeMLh1ppxxuHx7HLhGyJsDHFmvkZGJjQZanwvg1
hLADpsti8i9eeFvjyLlTzLId7t3uddsm6ZKG0gGPG66kcSjE0mfGZTwBN5akVJ7PU9v/rtR3In2b
LjFBeF8NFRYAfrZmYyapaiq2U7DQx4G8UNqKJtlaE+bLjA4zTUPk3NnBHeQmTYUJ/JkS71BrjJTw
4RLKC3RRoXj7mmd/BcNzOUAea+UsRgVWDopEf5wZXC7Yx4q+GB9Ih4804hUOJ0PNbD7+nBRXEG2c
dhgnMel1yHo/5aXYD7o3k7jl5eJvCheKLXg/7ajLrGwQ9ESfswkFmlO0VVqTuRLXGDjHypRzbbYN
wEDJy/1Qb1h5pDye6J4emP5diGXOv/t+yEDBUPu1wgRHCifE873rrwGZNr2SzRfVyc9lDZVlk4pJ
H+EDz2PUCNVKIi1npMaG3hhCGG99e5X6DNnDYWZNAyu1sZps9GDKcwPvJ+i6EM7k+wEbSU3/fCe1
pyRBHblx1pXjHENIWEGIHnP+4qcsklHc5zzXSBV6+/Fk01ZOfLkzBXuyhXtx5L9HpUvOhhm4EuZ9
N7aNF93t35U8GnsPwO+1eP9JTkNv7URoS/piQKkfnsX0lcMLZX/Dru3NVB0jkIsmaF8RDT/XkJCL
p9vO8ke4t2jaqTm7Hq931V88HyLf0WEOZSJELQZcz0kzb9ZdQt7qDPxPd55ICIS+sPEx2WcfOWm1
rCACGNgRn1Jrnww2pTwTH8vtQR4+PWCBZ+XoYVEbGC95Ya2beoGIlv02mT+e7gz26/bM+iRUUJRk
OyC8/fU5JUvpK3kE4bLAubvnwxEUntztKf7VcFwdj2TV86mXPiL/Ax/YDRVHULSK056R+UCQQeZF
GQLPW+Zk+0k3HJW8lrjLOtA74Omh7mGlT9cXaqsRECjT/CmNu9HwZ6XrbKwVPKnqrFnFukSCZiaq
scjqmv8Ik1sq6MAMiWKYjnha4a2uNY2zZZwkVP8j4zoHuYAfkjJke+/UwOoPoaO0rIEqoFgoXPOx
1KNQ93Sv1qnUf53E7PDBvtT5s85R+6zN/4wxP75Bh5ly2lWi45qooDtNMy6Wgkb36WZmpGzJBqNH
UKYpE/J4LdnSKrMRBWbtwILVHnB8GUmjYja16PYEHK+tgANoOqeLgHIn5jyzrdLMtaVC7EIpq6kT
086whbUSC1iBWaNldGFsgd4xM7EwLewuc2PbhwnfAgoAJkghdfUDzHfg9tDBCLGdp5IwO6BTminq
YQqHZ2b5pghZpk27a0H5FZEZtfOB8AqvLdFk2+fb+QfYCYwCEG1DBc0qkevIiWV6yGzdUiozkf8V
VzhSwC5bzWwvWfMAbLC6711b8MGhbwzdNl4sEg8rNc0lTKUerCD0MOmYcETS2emfUH/KFP5vdU+r
U6En3vIsJaPtpyzrKQas2l68R4FsjEGMwB+OGmiYTjbVfI4Rt2zuqDqMWfJhXi2dUkjRQsx0M/nS
aUlJ6Vl8HnI9qdJPPcGBBb3/kdSCfEg+T6LDftzBtaeXaTHuccwDtcudQjukWzK0hPXS0QEqQbdv
F4B8a+tyxM2snMYqtdS6PdooU4ODt7daH8kvVi8/7FzW85plC3dJ5JqIQZv7QWPQirJwd8J54GHm
QMf4hgBiwtZiF9WrgKQXOiCxE4S/739WT/NKL2KC/0HTWh4NnoG+Br5CHARX5hf2dp5qxAkXPMuA
ZasIInOXt379qrzXyFzdPmJbPpKMqv7vACyqhBY8ezymF7DgFgL/GFL4bbSYhP6OCNxz05MJNvOP
IXXbOiunkzoBltlBE52cx1RklfuFHrMPl2PrWyI5382UUbRzELxs7mzTJ5uQqSxVunfnC0YKxlm2
WEydPQxmKbEksuxwQjuRWHYjU+dk1xpC1JcVOYWVheBJEQe7+ashjAxxYlpXMEWR+VTGyHlTM4bi
9dtIVZ89rxiKMvE0Vy3ohVGGZV7Y+GBK5cuyM/D6eNYZdsy59radexwEG4WCezGjcuBy4g8Two2d
4l8xV6SG9BjMnkv9epc85oAWtMr5r7PdAuTaKWnLmlkmPUD+5ZA2AoFqaRsz+juN0QSwzOlHsO0i
Um9TAZiMtskaTgOH19s7lxjlK8/NGvV1URwtWke1mdp2qcZHAplJ3WAmNaudYzkX4uzWgb5R1QTn
0hY/Affed5Iz90sjaZXh2VA4kmgFrZ9OF6hqUXE7RhoDEIwyyWwq6yAzkLYdBTNzeBWSWoZT+J39
5tOGEOIzDNplF1Q6POH++dFqyLRteMhHgemVJp9aHdiqSO70I6qy9JoZN++ss9BgnG+Pop42Vwbd
k2TJaaAxkHSsKR2MP+I4+bpT/UfDX2TKeskaZoHOEQoEdwpDZI8I22tikyLYdaLqrSWlTzrwawBG
GKzDQptAI+26UZoJlFXKGhqAdxFP1uzvHrrt/S4lUhuSrjGsQbJji4bec2QLtCARVhnsVbqGJtI4
4p3hfzBYj4WqLIJo+/q9QDs0JX6QaxaCzkRIfeiuqokP+ETGNUyCknKEMK94oVg8gjwnalDVS0qU
vqqGvoekxvaAh8SFqSR6hLKN9Dz8dCGsjxEdWqlofNe4KxfjitzBTKYELvY4s6FFhuel3nEt+LeO
iDlKr1yVYIKPUOD8OA/1R1glpR3FSBGGVDwsBFqJ1VpsxxNzS5mPP8xAVjit4cen3H1pKmGCEgK0
fxCVpfUhGFs0m2CXF6W8mLMHZB6A7GmdhTfir3ZR9dxiiOeNV9noQNxLmssnyl9RjwjjhWMrbF0G
6SHZ7ndQiAgPTdQCW9yukWxQdJxfFlh7lw025se3XV+koBsY1fJ7Q6gyB33b+sXZtshN3ZLQALFO
zt7UaE4UbTfo/o8/0p9YowL37HT9GKRtrl5iX1bfSXua+Unahq/Uhxn600eaY9n47s5KI/Zh1O5q
SWuLC6pQ2f2yMs23aFCMy3pXBdnp07M8WBRtaQSCDrTI6H5r5LkYMuF6UOs6C+dD4jCwC5EeT/3d
EvStHeLgfKyvzd9HPd21wR/5ms116+gmUQWgLSeZ9qGoE7MlHZTOPEV0NytCr6XzyNV2NkKicvb4
WGKEBuoyA/Yw9U18zMEmBmIbvesYTtJuUmZdI+J5F7WwdMsAYnK5j92DSLfFpcMW7hrweKRunCRM
Vweb1UZZcqllcTKwPSVLRVtwLNJVJxTTUqEzdiiMzpF+lvLVqcJ9wkzxaafaGd2Q2qQxUEkfLn7s
XgKKzDBqAyFMTf8IGgu7CK05HtJbp7aViz3TFEzrv1TK27xEqMgBFt5im0vLX+VbQsK5afTSj/n+
qrMm0vXBgssmh8LFPqQMPe4SMulu5gwGLVQSixAIFVF9zeFm+bGsitrWklZl/XRcWkDjSgAaMcvt
5ze4llvKgy/IoqzbEf/XK7zKMcO/EXufhi75ZJtX+zhhVb56M/ksDk/yDuO9lnwhDlSgE5rkkz8d
lZwzufy7VE50Z8L1qlLVh3JI0yG4zXexa1AFe3hvxONnXGhIPVtcmI5HRA8hzQSo3etawwO8knHU
RYiqNPKAuKShigVqdmSz3uXEQw6G04OTfofupCJC1McS/dNHw3k8yPhGUtgrx6Zzu9U7U+mgqsTP
ukS+1Unwmg7RXMBFYcyN/ETtAIBwYZ3a1lwbRCHXIxzr4zJMlpV+zQhBWBOEiDaAV8xcMYefxDqu
zto0MTVp4NRmpbOpnaXf4+EKTwKvLkzkb4AEbFGNpmx4mGVOd/wNYPOySxIhaLcQ/KpipW1Afnph
CxeB31AJVmRsbMWzpt3S3tMcw+DrzsDrDF3TjJiHdyLFMNNfrEg0Qu/IJEsnaSg4wtnvlKq82nEr
pjoEjxZ4CVYszlUZHjt3296tsUj8EAniOWKWSgQGcBsJTcvcyJo2mnsw6cVFy3eW3ksino7iAGHn
ihQ5sJHFz23Lo31soVAelLVMG0HgKuy55lkXEt0HcDzLHXInT3jx/Ln05xNIANFUM6xKK5S9aoCI
5MPD5K35Zu3qnkDFPUzlllC45VGVuw7yP2RE8RhUJVkqxR8Z3AG5YZcrr3wTFSzp/7XTfABcM6r8
7/UB8Q2ZMnDHdISUgUI0TjXGLvtFGSY9ElIpMS0NBkLEsZZEoAmuQFH1Lq08p0Tf7jEFZyDSwiWp
ye3ZnvxEdPFaEcFyPETgjNPej//WWT1RRofGTUyS1jK83bBosjJP3aODfhbCgkirnmUiYovYIhhO
8/COj4GNyGf1ITIUUPcsaDIAfVlpjJl+EYcYaR5MpMJNQKk6zrHWhk/bIMFJtU8eC1QJle0uwjr0
nTMhOk3JyDs0UAaexcb8OYrgh3KXNjSIa37PdxLqJmSVJhaxDm1eTyryYaqOIAVZiC9FGmt41S1p
hqlqHPWOAHIoXds3ws9T/cixiwfvWArB5RY6wVTjgB+Ra8rzLGV9nkHojEzw0ok4NQXbezx3B554
wYVXI5e8i3IocLUBTn9QPK+gYRGIhFj/quRS6lQCMQEYu0OumwJIYoUVulvNNqbflr2Cb1GOXhks
c8uAnMGW/KX7I+vzKyAScPGuLDnHmPeqJ74nsAGR/orGiub1vKWFngJ5sJ2hqSTvske3SDhF6JfT
nZ2hVU7CMHOqbjBhyI5fNSRJRmhuzxEheXiqph8dhPcuS3hg5bhzUiEkXCZX8JiHusAwb3OO9tbw
HZ+PVZcQJbOyZspfDCZHW2LmBav3fWtgUhdswTXid5hfB5E67RCNbOjHtzXjGi+EUPTj5A+E3Qe8
UCDkvhiZp2KPGYXw5Dou94vn34Gca8SiDqeGpmeNqk8jNHWWEokdDtH0U6UrJYcTvv0dpeF+wTUn
pWc6CyVJeMZfv45b4ZYvQP/gmFGxKzGK3IZpqzd4vbPSIXEfcCcOCGq1rSSIuNAxMmTE+LfDHelP
21ffQ3wPV8QRu5Qp2R/eX28teDel9KnZ3wg3brS17BqvnuK2VmlykMGBQ1UgSy8SUZlh5MJ9/ZOE
AgHA2In+vWzgz53Aa3EOI1NBfn3gqQBNYQCwGEJZYEG3AX96t82+R0uKAKD2y+h7Rbl7/xsi8TbC
Ra9KqtVhZuuCb7jD8VksjFro+zHXrW9o+z9YQDG0rsJQoRxe93qBm3vC0BxYsQejPdc7YcOVj1B7
vICAUB4BZ2SKdo5Y9l6nU8D+fK2kudZaoJ1b5sd+e2qRMWOhkkQ5ih866E5k512hHXEZ+6WFxjjA
Ble1MhcheV/+j6gPBlr9C8oFogwCsBV2WVWQXfZtfI0TPxHX7GmONcZnA9KbTUnY7q4Gjmh9tFps
S2AVYM0WnQKU8JOm1AK+FGLJOJnUbzx1RxfZj0AfVrvJxRRB+LQYUZnJI+vBDgLDtNwC3jMtBPr0
D7OoKZKx5407esonl4xJwk5cdnlxu5QiNxx7mgIM1bKZtWs0zJ7/xTvMnnE6fJqdTgvTGpam0wEW
kfrTegcp+HWWQBp+N+qkfslbjVDDMs0QAg7Oa7Pi0BU66Jrv/ckYNmeUuOpXi+zKiafrOr9tY+aW
J+ZI0QWeBJKZ1NWpv5Kb2U3QdG/k9RsOPy8iegO05gf3kt6bD2tulU5zsM0mxvcaG3sz9nzAyDjb
zUcK73n+9bw8uuLfQmCkN0a+jcooOPA0lDNDdq/0mNy4j15nxDaRWwrEjrK5ebsJQG5XlNR+UEiN
up17zNIw0XGLiKFU7js9TZGHYr5+6EEju5BDmWx84cStRnrexftoiHRtYm6JLl5hqcjXqCIq6lIz
7Hboxb4pOk1Buwo6UUwe8R2UlbXoFtGg9IMR5w84FG96kigxjmiY3db5KnVf+HuWN7rVbTOsWFAF
6eA10bCy3H3Vz4/5ZsO+pz6/EcnXx+Vc+od0eZ24V7OYDOzIERuFCEtP8CyAsE+NVEj6XacPmgZW
o7bUK7InzYax0stUFvQ6sgGe11cLS4wEjLW5fM+F3OsD2Sxaeov0aJmuJIqr1EHWvtbHzzyMDxwf
ULTS9bEm5KU3HlGNqh7dZsaucMRE/yJhSBmYoa3THpAtc2rhHqvs2eFNCToUU7n/bV35A9vyPvot
5hwM0KoBO3Hg816uCVezyMZAOoXOO1Bn49mMVIpJ3Rw8ytVlCHPIaRPRwopIEuvznT4niiNWJpGA
xqDzqQrFmxIUB0MHitm5rsTMUqdWVjgaheuDKEBTdX2xycDAb8tukBZ/ReH+Df4/EhwlLyjISMUy
TGNuDHMEC19BP2gPMj49Ev+AmcVeacmkKQG1iQlcXiCxEgSCVg5ykOXdZIU66rVlXL0MCyyEtTbx
u0GTRfp57mM4dBajyEgJKClH061S/iHwlgn2da+otXa0egXb5GwfwJvMVoxFaI4XixE/OKlf2PvE
m4/VTkTj0WDrIbDDGe030y8zWnTRwscjU9Og8P/P7F9/zWYYJXVZIo/hmQOGToWqirFTQKJH4qt5
WgvDjHu7/1i8NDP7ZS4IIVRqg+j/8iR4Bh4n3Vfi6xdlABXlahIaEbxF8HXboMCw1LgLDehFEy62
ZlDeZwJMeZfY8PBn/0XzU8NWY0+cW9yYAl8LT4O3qBupOXOUOSMiFKrfT6fMlfK7WY4X8zUOy6r3
JkSHo4fGmzcbMwmVYPrqNZo3599EnzDvMldl4FKBbz4s7l2GFqg3lTZcppYncfzbMkQ3Xz3w8bjr
2TNePod+qR992tyX6rujlWOu71/FhIOs2L0EhEwVm3B41Mwj16S+g8RRyhsgKZadW/8UvAMD+vWn
LrKOe2ddVVDSPWchjABD2tntWuTuV2kKnlX8a4vrD1E2Gp545R8AJY6WZZQzhUhE1EXTDypsXXvb
ZslfwXaFET73IN/JppZcuRRv023I4wD0/C3iSwOdc7dobt4oOOCgNbbGqCtF8/VMWF+b+AKgm3yY
9UZHacvoKULH8QgIcJI/Oswx70Unkwr8+C9/iJ1e3bm1ypNEwxpWqU4IzKeGzLCervjiDVNCI+Ps
RqJbYKqdtpM+Gyw+rjiZZrmtgRFH4nstiqqPa5ZCvADUtoJ00igzrqoPB/VcD0TKLKcXHFGovQC+
+9fUST5F3I3PE5s3T8jprbhIjXHCdyjT7WZiTeJg8XlJulPa7ZNhZ1W9T02Oy71oRvyBdDAW+dwD
VB8ZHoR8NNmwTVruCcj4K32it+LkZWUjdEnbAieWbCu0eWXbvGJ/Y30QXB2Ga11wLxRnf4YxsioE
i7ocynPwpYUan0eIMKVmmwnU5LwP/hroR8PnUhvUdnL22yTAjqEK8unv4i/KZSKw4EPoYV4Kb8PA
17D+2xb2DfetWvyexFqmrcX4uEAQ8aCrcEQTFrdT67hBZvaNmYQZthtW6H5q8hFbvtQ34Qw50IPH
deAkdovnmeMv8Q1/uZ7Bh9alFefsXa6KUpkdoVzYD3a680Hu3EW2G4x0GuVL58/hDs9/Yr2kX02N
ubl2dWz9bsZr2y9dyT5zNguoN+YYrRXjWdLSqn8VQoGaB4RRCBlHqOWlDYGP/+Uh2ArW2LSx+7sj
cG403kAAAZ1vuiOPXCsIdjS4HgzuAbYVo4MonyH8+gDJ7vyP77Ad032GFk+CpCJdtFkgFU/W+n/3
obwAJB1tug2Xh8NGli5KcfsEfx76fAI832Z0umrlJBgma9nSmGUxc3ye12FTFUU74oC2+6NGIXHc
jGsp84AGk/1nyZ0m/xlqcOYim2xXur61au6lVzg2f67TL49E05PEBCgmmx2nQRuP39IStm1K7ZCb
TMjmanJ3sFm2D1V/KDwyH5/yV3jICEBFpVoiPwwtqszKf/ioFS0aYkVWVkPNmT1zpAARfV7aTCDm
Kz9Xtxc7fkO9IsMrWp0sQRXl8tEEAf1ppQ2L6LstfxOxvZaGo6/FHbRn8CUafCsU/W0H6gmXB/Ow
ij3miWFFO+erg/cyN1x8YHhHvEaAe/2lNFto3xRg6iJLVXQWnCH0LrHcHHTLdDyJqxOam4DS3+Ib
qgHpMV5XdLZLn8oLJWjYHdj6y7E/5RvZ/Vg2i6O0LhRqY3aZl1Zrc6Rqp+x4R1hl2kLKvdNexzoo
sMpYdveqR7K16HM9WIJrbhyiU3k5P+R++SnfNCYqM4b2Jmy/bvsSpTsToyKnIBTMuiy9URN/RTeP
teby36thVzK1yNHv8J2xUkaxR46rbBXzH/ImG578d2X4sahFdx0V4F92lDqQGaSfJyiOi8wRxlsZ
Bsb7mOTd2zjqcmcGYClqddxO3/ffbaGek9uu7wKoGAIGhCfNOpEgRmnIyykqOSE1SWc4go1WlH+F
YhM/nkdO4579tkCVWduNmmQQkvOjBnH6SpSFY0rgcL++DrfCsKX809A8S8005DbXKahXbGoQ6u5C
p0Tr+TRgxQaY0BEEP1lRnohZbfbiT22ykgm17PPoX0RJkHlvK2pHZxImc4yGg4GQFVgClvZcLJJO
N062Amcdj/ZvzhDdgJwv0jq/LKTtN28PzxvCM3A9Zm88gPUTg7KIishbNiG/rgZxAemXvAAKo7MR
CsZNiyaDnbWwDyM1J1gEttr2S0dO0T+imqS1w0LolS0Wk3IOn+RIYho7MV6DgNDQ0fHtnSLbx8WZ
e/MToFihwc/14P40tR8KAdRKpo3pfxepY4EU/I6dfGJKfBLkhntWMVE4eQmJmhxFB8Dk37nZ5lSW
ouHDq4JKdlG3HPAW6iKBtirzR98Do60Rg5DG7EFfG2mehatFUUAsZis8jsgTS/zvlGB6nIzeejdq
MbDVeqEdAwc0Z+cMcP1UA83TCwPi3HDW6dda9txEQNU07KDme62ZnHtdntal/7HfAZxyzk0rLipi
BQdbh8HPIzTC9/r7MHbrDJ1ZptGRgrpe8fSKHHDnE7ObFA96g56624XkCPpr8pXGyaz9entT/eTz
bDJsV5YoiaPvI7Y5mbkVeppkfYLO6C15YA136kCGMpTgdQ09yMKHrNiQqX4I5jFsIzeeGPS7SXsu
FcuQsv+OfKUSFp9QzRI0u4ATJQWeAuKxqck2WWlcXa5pm2LINSmfxofs6wOrLd4ePHCImbssuN/1
BvXEceWr4Tp+PrhRZoaaWIn7Sgr3VjEeKPpbEhX1GDx2SbOuoiR8FYhY5iEYepYWdKkeIHlvPFR8
r36R/3Zd1NuIsdP4bqu4VXyE486/1bUsPlSutnBEftOizAWwfS8dCXst1vTQwnVtnno5fC1wmxu0
BVSf0+eW74FgKQzOlRUiUDZVBuQKpHVpUcy5doHmkyuqIkRxoLhro8VomXV7E2le0L8mmBjWE3z1
3Q2qRteDk2Q+PYGMFF9Px4aOqJ0TvVoeWA7x5sUwXE5za3XBqxQBN+My01Yq/tZSDgOSQxMDdCGD
oiv0v76HChuZ6SLu22ct0GpgajBZ4Uu/R2J8FSlI3/PooXGxSaWnSz0+bdcoWlnuN807FjIysiJr
erc8MFpzAfwv5ljTJ6hb7ReJvVzJExV43P8csWc8Q7Y+cD/Sv68UIFwd74EsFjTog2mzJMAOXrhE
YpvtXYXpLccMkgRnH+GRax53kYoWhtJ5OGXdTOi8JcqfZNBsL5JeEOi9GpBa9pjk6gH9GYlJqTtI
TdvIjgkedCr/UlV8rYqvIS8QgB8PUIsaI/am9jDgO71nxTd6qhbmXgBIpt6MiVPGITNHy5iqlcJx
md7qsX/ESowI7HcgJsDFUXk9KN7UK0nZLq22f+fZdoC0q7K3l7XeQ82ccGwfaO0ElD+iJc5ponyv
+Z8P/iytCfUsR7j3QStBUoAs2L9U7E6LT/7RxMVXU/BkcWe4awgQC7qhS5Llt/yycrgXQftms/WE
SzylpiqvrEi4w4elXvc4NgeBESSQWkJoGaBlnit7O0LcqxbndWrUFaSWdFzzNHFu6tm1uA187SOJ
ErGTJRUfGLoWnaaJVL8RT3MENOXtsSIJwRJ6OoJYpbMI/NisR5Och89V+5HRuTus85XYIzCpEZvB
mD0fYu9XwKynAbGbUro7v2IeVhVkhfQA6Xg/p4iVrKGf6VXJ0uoe47np0AHUHEEGRUAvOcblzKMp
F+zKNBVbmbxXuql7VXsHSFLtndJRLmyjUu9t6NTCQQzfwIkvnyYJcEOYbhp3H2QQbxg5hM5gM0rx
EtS7f3bMnFBnIn1wqLPlX/TXc3oVmF2VLFdyYrGgRrJYcM+5OByyl9J43B8DYTdt8po7LNBPYom+
wp6NpGxnAlidUCMOHVx1ZfwjLmcLba3y4CYfqlxKT099dOINUUAC8M/WP3yDUtuEQWqU784/lCui
5/t5BaRghwVjPKFYB5aURYNngcqkcUEYyHgBLo+VZb30gF9cTqGJbaq00szOuYWysi6yyxZGXZ+Z
lm/ozRt8oAKrXfSk3ab2D44u/8MOE3IBFdAScig2UBQKDAOWgGLFX+oLRudXMGhpWmySqt9WxGi4
3lYUBEKPM9xlZKDkNhv3HHsjmlXY3gtw7WSgMhmn09paSy69MVvETUAQmaUyIYNEhSbjaJvg1gwv
1VDY/uvWTZXUdoNEhx8gZlY/xUdYn0vnlUw3FsPixqolIdpTjDo+ios8dVJHqz+D+JyDwjixSXhO
SQc8XZHahamZMSfuPIsbPb7yzh6TPQCnF5Q3aruV7eUgQ0UZEdb2NpXe8QQRcX9tROWWUTd5Aika
fxNetRyTFSXdATijrhvMV1vYtKczFMCcHFBqhSWpmXcSUq7T/0y1clqIUiSAaYNCbtnLHg78LqVe
F6dFyVLK1PMmBSywuBKbFSEaC9yuQ6lSx+qaMMqwTuP6saSVUPbmanitJku3GS6KQhVNhM3nIrG1
qER8UtgK/9WzEhw79X4FkAkxnHyhMDZf8gXDNAvmEzVR4UsNnLXXgEaanhSUtA4sYvu04/zk97SG
ZqEdJJbLzS8rF2pZ93edunh43mwyL1T6odnivydKo9rvIQxQL6ypSBqyEKjQ9/+MfPIeFcbEm0aj
3sQNpX+T6sM0t+HH2CbbhH3Y/2PeuJnfu3C9z3ay2V6NoaDgoCFGDa144DjMF/KKqGgjTfHb7sVG
UWkEiWUJVAukAub/53kRptHYuS/0OaCQ3//+nrrkKBBmHeTKHk4fD9GzOu5VL5RpZvyCX0X6U/zu
oCm82EaaTQiJmE64YOe1fB8PzeUn+1AlF12sKsSTWCCFzUz+R7WpkeKvsl7CB0NCg/RzKM0vM0DB
+47PSDULRKSbsxJDKqdJz5H1fduCuNmJPY5MOw7mGgIu1Jm4WCRVt70xira5WGF1JQVUBqSCTwLq
S6oP69x3BvtcvO5ZP8JGEb6aR0+Ug4bmW7rVd3NAOdmzvp5zzYRdhOdy+hygD+GYGmTrzFgsZMmU
wFPnNKYpAfr+ZveCdq3r6lEeMOIafuUQ9nJZoEVjTJoDKk/TaBw/a+nsWH2Qtq1hdUFm7t71xYBB
pdkS0zHlDrENDOrfxf4D3i8G8BFWkyoP1kXLlcPrQu3qLjgLbJzisVXtL68r7WmnLCiVXeqqOvac
SNQDxlo4s866YPZ+XxZWv/Ie5/OEIYmaXioQoLQTs2ZRhRKL7O1PDGtfEGKgeBqGNcwBUCStiwNG
nFREVvr9rQlAjPj7nwLk7V1EMZKki/TqjZFzghqyE8o5t1yuw8JWFuIGum73kKxQMsEayBJDljAd
4vYqyfDblGLNPkdE8w+dLBpv2dLA3WNHUek50/PHF61iz+TVdiDtp9k7mt9WkbcaELwEp4JNOiHl
wugO8algSxgo/xM1/eIYCZbpw8EkqUl6KK1XU5pB9l0YKMkAFdvRpY4c18Rpp52H08H0l8wQ/rP5
ujzfWJkOIDGssXHYCqNjiMKnd6RpcMvbxFIpnC3mQd1VCLSqI27hEK0xq/fdKZTuR7qOWGBvRvqy
2NGGDnsNcSbyIcTmq+SeRoLGcZvD0dwphgIgov5c+/ggJhCoIPUE9YZmDUDc/+1hNqCEdLazwds7
9g7rHDXnFRnFf9f/Sy2W1akMuHsKkpKxwjRauS2K3UzmbtUBNsdEBz88dPIIOT4/kVdKM09I5WH/
UWzOeBOW+mejIHTIAY6OxN3cPkvzKBLxUhC3bbDN/k42n3FFGq7eR3lwtnRXv3Wi9hjIK1ipEFxd
MlJup6P58pcoFGc5m6e7RFDcPI7V+0rnokEZ62VJ48Nejh3kIpD1q5HuyOgyQfdWB3Z7wftOzcgl
0b82WohAvamresxxQdxU5Y6qbstpJAB3K/ByOpnQQEOTJiDWSBH9dqOOTsgwyRqdx35GXaH/fF1K
uDF86kUkBnNKXHkX8Hy0vtCRpxme4XphDkQhB3JZC+Q6WDeYXEgqloyRNSt//ERWEXrEVOa2XRH9
TNmzqsyrb9SesqOaAdLSFlbOHVDo3/8W9lhToMXDFS0W2jFvEVDdnTT6Oc89RJDIOHuOrzsTCaYn
j1dXhbrMeAEv/Sss48wNeXfMXdRrrPRffX2qgKc7Mf1vWVXWLAXslkrBJwDuTQ8mXEURZv7AumIS
IxT614ODag25VLZJPKGFudMm4TKBwsYCsjhuU1K/napfhb46BUrSsmqWynjFxJPZkn++nvUu4W1Z
hgKY8yoTcGom6Q9wjA8olatxmkTSEcqF8n8EC31QHAbQb+vfWqeEhB1v/aM9m1WMKRPnQuspMzWT
ZVKQaEk8qgEq/W0FMBFPz68mpCaVeECMIZHU48qLeXWUM6MPK9hkyHDHK/SEOIgGkKLrbEqBomhy
1oCwtCYWDTVh8WL1ca4YCz/1iqUMcOBEiYD8OijsObgKCV5Z8pV9AfJTxxdBmICVOuiZNSLQl6gv
RZ/rUZm6at66FR390snjn1aOnmkDQIFQZRKTMHG0rdqhXC7UrZUcuYCiwGc2ok8ECGnPDqekDHlH
5WRqvjf0ErG7B04zaBkBzKR623V8fiToe7SJjSDTzSHgCeukhqieI+G2ZDhxBxRUO+gO2mr4o9YB
ERUQrXyf3Q+rfXEgNQFBGRHEkUSNRcnxl4edYpZ7ENWd3y4Oe4w+NSQOzjyLhSj6SuPYPYGNaakZ
Fl1O9kyave9St7TzvWXhkdaWhB7Eip3OZrTMlA8JiQoXsBNzL77oMXM2atYLL1LM1mcnpm6D9U1Y
F4bvnWFAjpKI6mdjp6GjxdEJAk033c8p4qsAAc5DeXR5oBNUpqtOhWR5pHAQjaJl//jA6xnk1B7i
JeWQdarHoVlhAOIoBuWtgOGxFcm5TQZDfUc4PGEe8xE0b4MPw7EK0eVPr9UFr6pkTjiIm04cPHFC
czJWEY0pD6kQ+CIuPxQUeY5ZCKCarAJHiWnop9moudak9WW7i1fAslwA8Z4z/NnEfQADFv7ha0ae
N7NNIePsK4urF+iG6ZFsVyXEiAyJE0Xx81KNyJX+vw1/BXbAdB0aeCx7PMBkJHKIxBNAKG9UBnaU
RbIA10Uvp8DiHKOvtOMPvJLuSa916fmJExwblhRcSdXskqe7MlqrQlBHjAFTIa3o55tXSeaFP/wg
LoSWtSNxeBa+U9ZqeUd7TUGPTNcUKFai+1ZtVS1mSoG1JiBD/0GnV+id95c0FvEdLwyBU7B/u9gi
FhWU41I5coCjw3yaUagBB/q1UuQTK6zXkWOykp3pvrQc88S66f2MF5RXQmiGHWEzX0uwzyImtkTN
7OpIcZCSrGH7ockJeETmqYZz/XOfsvrMEDe0PJc7nWIpd6YqOiWWW03hqoIdKpGBA9KB4JNGxp3D
PHIlEJZDojqhrweu62crGyUVJHO/v6MvA/YlIT3EBMcAwY95fOezqxuXApWT+y77SnbPfE07+hAa
iYW6Mc2lvBF7lXzgszvj/1KbMTKmv627if+COmAtJiIFxB0qMq6AwJItn95VT7I27YkHo6jMLFsU
4h711fBxCNaFgLVd20gpdnygWOFbCEl0ZJyectHIunby72o3tPHIaUAg4GR2UtSN7ZZelJmw5fvG
9jI/haRdyMqS3ro+QtQVh5vYOGIFHZl8qrWVsWRLDINgjLcNXrPkBjetffDU+sbBAtkZqw5Ije4p
yq/oapo15GaE6LyPUbbPZyZitrAoU9GoeyKU0wJ0ROwCef9vn7YXnGPgXbqV36v045EVwWNARzDj
g0iZbsFeYW/aPpCXWe6OlEqmHbDZANTf5C04oV977afWgb/DIXcClgKFgthZ6eN0K7WMXbOA2D03
XDV9suPyy0EjWxJNpOOAkf8qe4FklZa8GGBcyL5HQ8VtxaBTU1EsrXYZQ4a7tjQs5dQYRsA0RAOS
mH1xutPVejypRRR9Z94eXtSv4ZFX71jNfF1hoGnGCF9/7OpINJetRYuT+h76BMk5cWSL/Eh24+NQ
+2uN3c0T+PDcsWc+szE4ooKbMnFbOoasXrKuHl599L/UfxaZSkj+I8ZpJy0e1gixEGBkCg/HRTVg
2YMUD7oESkKNEEAVjvetbh1wGdgPIwgQkTaSqo8LmmP8pi5N+9t/jfy8oaZmv2AzVxSkOUsNqvja
KpIloEQ/rE8HBhKiNpRRpVOyG3Fphla1AMB4Om85XwaD8ZK87WocV0utSw4kOPi8voAGQ+sW7E04
A2OA56FebZ+mLvHdHrOZ831gDq6W+tSHDgUaXz7jdZO8Zp5xlngOcK3S7p2fBcS8WSYw1MTwzbiH
qFvq9A1vARHuES1r/wujLkmps03edQqtViRBF8+ROOObByB/MyxyDJ8HkYSPSGasgRj2+JAogoDa
tzWTxZDIgPqWdx0DLxzo1QMgRLBvxWST27k1vu3Pn1nNNumrEjZquHZIS3OZIrVLxUO7qqwOzAnN
PhubVMHkoa1uxX6wUFnhjc8he2zTw0cQ2ZFfhWH1zCunqTj8Vxb0GjaiJUOa87U8sj02H0BWvadj
nyrQF9MFLCKsvcBje86rf7YG04QnQfnRrtccISSU/mMgsEUdsID+3OKyLvP1T146OcA8TASGL+G5
55XMcYCGZBOU2Kp8BHwPtCxXzjTGpkIulTG8+AD96GS4gLaorzs4WfI8g7Iwf2Yt4Q/FWHy06nHa
XNG6v4JLOLe+gvR9HMXn2FPlHwAQn+dtTaqF1FbaoEh2WhDQBzT2HG7qNPWEAAQbWHvViOMf2qny
disZ0TeTaR3ke/AzzFbScevT22JqEgJF48jLVXaCe+TBxldF2t220vg2GJU8tlmASMRAMnui80le
lrDTknmR/243K1VPaUHB7GMb+ZgP+trSJOHjwqvQsrR/jxI6QhwUfpJxPS/bIaGhh76kYByosYZT
ncls/uPedQJBI8qgtKKRaMN1tlGvRuOZjDoM5/tuutVE9tMJsnqfjb8cC2jsD6WzGvPDmvJZff0J
eQNmaIAIGHGM02p3ItcIdliCmy91EIU9vpLXPyCNN0YgCF717hMSK0YafD3Vfw48ciSgtoj7WQAF
DoG5XHbxHpKU6McsIJZ43qWXlly5V/2d2frf47n8NqgzKcosizQUxEo4VkOr65Ks+HEnzclp0w+Z
3Z/HLjSQHL9mdK0BuRbC6tzFlChOtBeovNd6CZZZOlzMXOMXIOhqZZYfswVxm0MJ4XElnH2FqoIG
9kgbP0Nf6m12wpqUEKCXhhHopykDh5fFk/xZZ0DobvE7ZsFln6QRw1Sidi/n4zLMP7jt3+7qiku8
344kjWm4DOTH6Ga20h3MZoV7JgfdJOe7Yg9TrBHi8CLKTCtdgjIGYdRwWGRPheH+hptp9yL4UMtq
z3u5I3Ml1Czkr3HkBZMzi+GhRz+RhnHMyeKvjCEzSk5qUSW/sqslxjlADAlQjG1IcRk1ozPUXiPl
ZDXFeIKGyeSU2XofKH4V0/kGoBlikNUn6aqY0F9qi++maOxy1qaYi3/El/1yS97wpu/D6IKaVakK
zC70aEIA9Q6SxvNfsmjItJ6p3KOgNv+WwCZR9g+8YhzNaLNH48d0PR0733f5Crj4jsYlH4vdRoqV
3HBFrSzhRuz62Ke2K2pZb2dvCNgZL89T7hd044GET1p2imtT72Kuj3i1VbrkWMZcbXfPSIQhwAZ4
k4xrZjMeFHY45u9KqKCrIVW+WsMpua1Vb7KmlhhGWEt4imqiRa+RhtirBm8BiMppgp27kzUL13b7
dkR7++2/TmZQlxuxBfUArygj55xuW+f7FHEbvjLnNz7N28vk5MFrLhZf0GTJXyn5dDZh0gxyC/QW
VnGJiWApkHzZ0nZ1VJArptUsZjLdu9wA/IRHSLKFR0jLzSXmyi9LcilEr8rMGtyUoF6IdHo+87C8
ngD3oWdcLNXee+bw4N4pSjDRMVL8vUKMn25bqtmIBl7ARJh8q+cbkgt0m73+kq1kyGLyexJ45F2+
rU87IQShj9nf79LmsU8jT/ztU3m+thCs9JcRniJCnje4a36m620X5H3ApfRM2jIoEaepQ4L/Ky2Z
agWR2e6fZWMZS9xDXiqZexC6sr2y2/YX9nhbadh4zKHECKRO7O5inF1zkqrudUjA4AwjGvgE7Iya
m2TPRqTWR5qVmbve2QhhhJ9GPrdRbtwqD/g35eiIf6Tw8QOXrY+f/iaTcMtyAFCAfuspHZwAWBfc
PITtqCBWpkN2TxfbYamFAeaGZRlfN/8pnLFT85Y9rer1cVp+qMdLVGSmoGm/7IPa8JF7pSUUnT7H
oz18SjL266xmzxd8yEVISMd8oNSf1ylPr/C9/qSKg8v9c3UkVjsPGaYUbD1N3uarA8mqLpEYFfoA
BqHGEyy0s7K+0XBVpxad6sD0kcN2DDD8u9R1w6LtSi6P0dlAutAazO6/6A8hu8Ht9ibFJ7agcH0K
6w5WGsSfEwf1e396/HaYqspxvHT8XU3x/Xqc52scQBgFtJ49VyMiYIDExNPHHvOGy7xFH3C7a7+Z
UQmMUd25PzzEGVHu4YatiLEy5gu/vHy9vrvYxXop7kwL8fkRyR3Q4duMH/H0qhnRnvWqssx/0bX1
UbyTRauGYUkMzJ5PGdI11eFqL8iGruxlALKL59pqyODEizf8zYdwbFUfO3njfBYLx4EpKVK+McUM
iuQ5NDJkrYvKzeVn2srNnkbX+e5T79XAasyzon6ypO7BSGjdlivEpxjbfrWjoa2t0vhcQq+kd3TK
COV0eQvFyHMMCxPnZy2EN2B0s+48Ieqs5uSZRaW0VpPfUs9oaa+LXrPdDZC2X75JIpbVX2fPrT3j
AyLed6gop8vhbjx7WhnC16tS037MoassH4nXdrusUVRzd1vMrNV/KQZJBpRmEh3VK4arjVIlUlKG
f/eHhn/Eetulszd8SWdrTPs0D1Pw9BqOpF91GQkkhzvK3sTBY5uFA/QMBoScxRs0Tb5AwLw4HucT
4CuMUCooiSGdesh6OwHoqTHckuDUK5CRVPCFlvmiccFOfQlvNMkkNZN5VmfiFvg6FFedC9Ee0hvq
lJotaUbFguriVQsWNqdEYKqfT82q3C5+Ty1T+4sJJYcgab0gZQ1JQK/91Onm2FyPuLK12hauFiuU
x03tJ4hC7LpEhTS5rde2PZqsJkD5HrDjDDRWYh38dYS66jGBrBoGQxMxgSYgDT2YXBrogvZeioSV
BI7YS6QON4VLVPINQ0SmiX2Ob1m0QaWeV74XBiNQitL/t0yM9xvXVd3qOBAYjTxPsFM6qhi+0FtI
N7zg30gO+tVysuo/G0oSRP9wG3YRvgOyFvq+Q0bNf91vKoNgzCBh9BKULwK+3PBLda3JSNYjPLtp
/YEt3JE1NxCQV747JSyPZPNeTF1FcdSRCut2jEsPm5AtUWSd+qVhvvpup7W/i5fWuA1OmVM51YKT
9qBmER1NXjTns5j6TlSHDxhNLkpOB2jJxEvzu5cWNhUty0nBmV0TcN1Euqmp8fgaAzKwiy4bhN42
6FLakk47zbTEKgrK0J6FMT4Cgh5eNzrZ+BJ+MiM2TxXzRvxl3VQP1BRsqPiW53b4sQ8+G1ZpcVV2
lCut3ANg/W5rtXmuC9b+uEy5Mg3wRAQF9jxl2PC4Ac91WJAqBpInf3y9/me+CH/cJhK4AlU8T8vY
mPISvaw22I8gx0frbkazX7RkXVThh3lUxbjpnm3gsRWqToXpXYIMsQksr7GUrFNIL3sHVHDQrdRA
gp0Wpx9LXoMOnVJUjm7sqCFmakSoLsuGiL45U784/Q3esI4KE/rV7F98HbuL/Rof5pHA1js+831h
vh+VeTLwjvRYvspmEGRhR0v1DEvc/7pRHyb/xMyBV39rY12oxFdBcu1YN8/NbtdqNT+sXg7zQQ0Z
9o/WHem80WPUFPWdu5ykWXMKwyDV3wq1KCL6DLSo3JnhV22L3p56JiaDzXZ23XXGD64lOjCs2ZXT
Fgk5mZjBZGpWctQFict++bw2cJeS0OJEH0Rxrjpf3uIEL/wJKwRbK62rI0CReP2yXgVZkB5eWiLU
+t9HhvW3nYYOT19o1UcioR8zj/8SCuXyQEmCQIUmPAi5q4FtpBF6i7haXLIvboi9IOW73bd3aYJL
GtB+JYDT8IzTP2n+oO/qgegydHYgDNRDjhOiVlcgMDvBxi8gM1aei3EP6O1jFHi8CBl6R2uWEK12
bjPAXqNNySQUz96WmVvwgOhJEib1yjd+xAYcIKYRh+LFU/rIUB/fhTDHuarw0rmJCPOE/NplJwpd
9O0vDiYnQ8DMkAt5Q7obsvUd412U+wO2vdFGgxCDug5a5PVu6bbQWDJeMVnUZcHytOTOCMep27lW
MKCJmmLLeXHGgZ8RdmhLewXiIKhp6veHBFdgwXP/iQeaONNXj7XfvJz2aUMD14cUTG8rFIZo2zHn
arvnnRA/dIb7xiChkjfLblsyYB7onA8yA/HERzGzHRYfRvl5vtPWp1JhNFr/cKFlgjyOSLFnyWEX
uaGIcHOzg69p+24wMlLZIe9hlDq9ntOCnVHXvWEKcYs5HPKEVUGEOgDTOdkvumCfpSGKDMdDV/oP
yMqUUpxeEMZGdSgIByNvnAa3vJCMv3M4gf8G5GMmt7qfxghTVpEpVJ81p+Ztm6XyCK8oUHsgJ9EU
V2GAYgGWUzdA3I8B17PWjryuUk8NG7N8PuD4o56AuZyDA567285IcHB8fLSOTuOwjGvOPY5GlJcb
d1lZ3wJqBogN9dys4L9LP+spGfaLiPMl5R2xdwoxoOGaZSEYouZKB02Im1SysaZ6EKQVzWXZ2jcK
53pMxLvd/HN8phWSKeMLBFFjI/mEpnQzAMMIadr3scH60+Z0GA2nkkhGGO5x0RdRXXN/2svWhXCd
TUv5+sxHc1O61uu96mfaK8oq2aMaFo7Urx5DjxHTdKgo2OwUCawVJ4ASKh8oD9pnpfRz16iX8QZi
HQZfm3lP0cehv0y26Wznwr43iVBfpXRlmuLXMKuJxpAFvTqt8hSq5FZCmyimPtB8o7fn0HUFJui0
P1SBJUqU7g6NsRdEyfl22ZYvflF6pJesOXlyzSA/7TgCARmK/v9wAIh5ZmeBZ72CTni36hDPsNqB
Wg7ShATE/urYdQIBMKcE/iDv6F2zgQ9x/gC5j0uCud8v6wdcZyIM9b2h4+4GxFHgEih1Dw4o5cE2
47cevbGNfHFlKvzixJdj9w9tcS/Nb8qKjaiwYn5BEEO2C6SmVQMp7GklAplURyuq9A21KvqcSDbW
ev3mKtKyrXk4wLnbYJ1OrU6GOI5e+5eBvICW9cFW5D9y+dXclIKQujbSyWehfKmtjlHyPQLbKjbV
G+HylAzJ7fz0tSew8SUd+lmA8p/0s0lCy5RKk5LgY1cjdba16Diovkbu820vwppkE6KQ0qS3LSC+
UPkV9WCIs+SyRM8XJIEGvaRBQaJvvbA/tOLlsMw0o4+7N43LS6uQAGvSIjuiDuj4RO7Yoj2+xMKU
+/rblG/bR2r6J3bHb8WkN2y8jzhP8ka7tLQXNgIweHJzinrdza3ki3p7uurr/WbTj0BDO4y6Kaez
qEbSoKX6WMBcoOR5ZtYWlyjx6M+sq7t2f7+5UVkRPjPUzqQYiwSgpsLMhKZ8sKv0xbL3pHQeLlvy
ne0lIytHo7al/CH7Rclw3fHueX+kGypy+hVayzrlWVUCKZ4bF2NLlpylf5wgAgHVgfC4hFTel4+L
1QpuNa7liheB7L8s4Vho4a7CTQlR3ywjsduqyH9gSPTjFDzEFBkuYIEELuqk6fnV2015yDxT0z2V
bIIG665zqA6999oF4lXcrsKkCthmIjVehIGk8Gf9yhoO4Q/GaMXVaxO9AEctGSqHBS/Te2EmkPGq
I9Dl5sDxi6pJ0qLpgTmLJxKpqYCf++M1T5d77baoqE0BJBwhQhle7daDyvABqjXIQNAyQh7RMrfE
nJkncdjE7stcT033P8/ayJPWSyFTx+VgOyXrkSB+Jg3aMww9HcHa6aORhAe81wgD94T9KEOqXNHR
C082jkWD8s9+wQsHkS6oZaPOGYgSvuYQR+/uWjWMHJLHlTLTYubNr5JQDXH3PcJPZPJXH5ImNHmd
nwEvzfsbOCNFVM1EHbip/TZ0pfRmMOMZBgbXuxD2EDYYM6TPgReIcT2VpSxTkbSaSDHxGKyHiZd9
eLWkF+mP2Jkk2etTv4KK6PqswWdX0vBd7YS00SpfNH1pWkQHT/xuDjIcx2aUsIpS6ezC4fo1j9DG
Px8G639MX9ShvTT14O75N93Qvk0fgWtvHOdN/qRsnc/tFSeDAdf+GI/T4LWdt4UVrwyWnvHqqn/O
EfA/GnngiWNUkbvK1c5Ej6qp/Y5r8LJokKRSCbmKTstm4O5gOud678OTuEUjmdPbUodP5+bUqKKo
TNTUceYJ3iNgYMx54dzj2eiDX6VgyT1rsoAYfHIKin80UFtJyNvwZMbWhTy1MBFjXvm8HCcVTqI+
xLEOyFqKVoSy+UpW2BeJSwvV9ASBB4DnNw+EUq7RFE575U7RMKv8rd8s1LoV0piX2ds6PyY3VQ8S
k3T4VeAmk7lDzVFMDrcj0vv73fvtV3h7r/FA2S5sb+vuPYvaS6g4kpAwVhixaQHtGUhd6A6juQbw
oYv9wten/U3dEBD9wJkErcqJH8WHh5OPLslvxbWwDdvvdmI3sG/5qtgKbjA8nV+BOkwe76W75IeS
7ClirUulYvzvAtRl/RdcbdV963CyGduEVBceGS0BBQe+JL0nafo2q5hRwP/U7mP9O7wS+S7vL6cG
wp2JfEspixXZFZJHsMmnUgMNwA8HPfkh6Q9uEJUbmR1G9YDxJ6LT5HH5G5ENBGNcr6VIl1OFqR9O
BWMyBxoSjWVZpdcUzN9Y8KL6KMo0S6H4T5i8kuUkKW9KFrimroIquRMsyeOBCMMW1g0GOkpt1YfM
VBdIfGaOTuyNSatie81xXIg0ZYivPf0bbHswsGiLpNrO2G6e6PwWXzdUFr9c0O/V4QbxGm1nVbRj
MwYsj5I0CvH9RaLuR2Pb8Ee5MWJYKss2EBr0kyLGQYmBIQKLToUtWRuddGvwDaPtrXkCOsGraJ4a
dtq5Y2mvAyNamG2DLB+8O46s/7ZoTd2VdkaCtUGjcupodSvD4oi2NMnV9KQMIbMjV6ZRS43R1n7o
gS5zGdT5StYD/3s6sYtZa+99/dS/EDymFgOtHnpQk26ovmPxrj4afOsSQBwCu3svoGIUAM/5lVxj
HU2dVc8nQILC7J5PZBAWHkVsaJa55/oMKNEdCT7axiD9a9TSEQpz1TDjgVSLWLF1kBPOygKy54Yi
ytnPxL78J4vhj7F5XcG9gY5VqexEhMkUgnHdgWqV+/CDUwoaPAomZH6HEsScH/Cw0uSzfFDiD0CL
ytlR2Y65o7JKzHB3QkIm1hSHzcOoMXEQsiZrIlmR75/Mu+jaz8uXpzKJSvHF5eJynQCwq8o+9yXy
uqVFJxMsnIxw16ZQheIGPBkB2zQhGFVNaMscyyldNnPC6AFhT2D3KOfFpgGIdYCR9Qha0Wd4r76W
gDGOw2ldgm90LCvj4K+zsKJiP6Gmi1XbqYE35XaokS8m20QqXSoNAmeyKN/H8jfD96EqMfN6M7Ez
0+3Tkgf6g5p8n79PPiWixuzwls0PaxpgG08cKyHHqGeS7LH6rz+eg0zXMDCFU3qE143ww5z/t4qb
1vDi+4pD7p0Jz2UjLzKQK5EWVmnl9fq+ACGhKiM8CrV0tYfCa/53UjDNhYtg4CTby2A9qNunCrJ1
kJbRJwo3UoEJGJRr8kJO3h0NrIG+0qniKQOliOtLb68eBqD3ndg4zNSEpOYm01I1T6rQ+2is0HLL
Cv5BnuNYa+WX3gwUFxEUiV+ace/zhr5+tyrYrzdnsPRCi1lpYYi3dY9CDWyZRqHkTn28/O79NbFw
I0lz1m1pMryz9p8dtQeFTcpraIwRWFUvIa5klM/LRT6YUBQCWBKzpEKJEK39NGiWS5s89l0AlkOp
M3vX73Wl36CVOI3r1ufLNyPUIUC0BLnjaQMXH3TGxztViqU9cmbv8lEcyg8LDxu3xkKuGj9ug5Eo
n41t7BVplNQkLkg6nIFeA7oH1JVDQ5C9LSMMtjch5wH6qxZBOpsjwMx0BQzA5Uu3m4TyNRMape1e
x2ePebWfYK2nrIz8w1klW82jQDOfPDTNv4VxBB+noASpnERmi/XADrQ9uYzn/rseTsVcSW4n4aLc
l1nz6jCJKLbOxSre1oZ1Ke3q3krhSURAaBXShoVk0XMCLi4K6lTn1s4G6o4XjFFC4uQbBv6uzi6P
0LzkoOPgtfQhgq/l0PN6c6KmW9fUPMNaziKfwPJ8npqrrjebJ3tZBJ/6qMZUguGGQXCSnRbBQxEX
A6VpmGvyWLguYcvOQeYPCb/gPOZusXIV4yQ/xdjF2aVET+CbmDJ3CAeN9i/31gGweREJZK+nwaGF
NGESlyWmH+E3FdO8ovXIiQ9yIG71TdfH7lapq5XV42vnQSe+F+RFqTzfyx99JU5Bq+qtXZQ8Njow
l4VzaaZK/JrovvTjif5LiWuod/BlYwSeabZruazUOAefd/XmL4wXY9P1KYyuxuXJI2l+uGasI5xz
wPV8ifKBziZLeIo+YW1YMhApGngOXrsQXqEqeNgKypsflugoJEUlORgZAEzadXWiNbegRRyQylk4
Rycyj8JT2p2O1TYGY952w7klFoGeTcZLB9evzbRJ85zrJKMTsJQEPh/9Y3hCGv5lGGBI8Dh3ZW6c
I5YSt+Vp4/J1LAypx/ASojYM7Bvu2aXH+o+JEbmMZRT7gIFeZ/UgZf6n3erof/jiSrHzIU4Y3Xbr
TRhhvZzCBddB6IfCEQI8wtlxgweF24t+RsSXaXVT9mlm3D1pGQe9wC4/EIlR1HO4UYC0j/csA2Ym
6ik8b2bcmyapTzEPsBPDc37c5K8Vv8jLNSDMpmvJ+Y/16OVX0S6jHP4dHDZyPFfaCEA1D0frbnkt
Af4kmOkDCAdQBQ5maHwKItpVMHAZXs9+ZAZ/j1eBpNPC4tGFj2Tchgtz5JCW3w12DADD1Lr5wm1n
C+nwJGwVu3UbkOmx/zK5dxetyFutKRcdX8rnVS9BIFZsD2YhFZZhSh7PjGvyHVC9yE9Gwp9SEqBO
jLBLZLlGmvZqAa9K7tWVnVN4jyf/6lE3BB2JUgMJyFb2LMSgLi9mK3EfxISjusmMfNDKPSKg0C/E
yl1Hyg8Ugz9zHSOfjUn5tI62f50vmfO0TtdwHUDKyOIpJsyoWWjweDikiEtXARSpjZOF5xJu9Hrb
4g1lbD5D+R7UsN+f8lyOe3oHXgXIdtENNnyUMmhZCfO8Hb+juU9MV2UpDb0Dlcf46C/UCdm2PkG2
Ub6IC1RISaZ8TXRTnAl0JY08vtqaztaYokp4d8BZpdNliT3EoamQ/yUerYILAJLDXDSyxDTZ6u3C
4JXH0acxUL6CmxPFnvgQaDH2RU5BpQ/mOn3Z/gVUdK7GF9eFlIBwJDe6ZgQAp8yJ0j/mOltlZpOH
JmUEcwi/N0wM3bvmYNPdnB04CmhyS3W8nCsEeGzdfLwFfR1dHbWa3ztrGvmX/u/ndOohuFlGBCal
EPC79A6E3aE6zW3I1xa1BGEs70o6vaYySB7+qcaLITnE0CyJpVvF6mgcHDgQWO0TdRuhVd9So1Mj
JcKJwnIQPjFZrBBTq2mPyvYbaTV112NobjbckgLDAU+idXqVQ0Lprd/JsBq33CX6hmubutUnWdEK
I08FBWRIzhKBcKFgPaAayPlEcBjZ2VB6iFMk79dLxBggc95nfDKru+a3JgdCtr3uA0OrNXJWKtQl
ucJOuXBmJE1E9Ft+5kzWipXW2Z6tLA7h4NdljQ5uqp6a3/Oew3/XKqeyXkgRXRcFsl/MaCM4RnYK
y5leFgHT0T+LryyTUzK3BRfmeGWvpMs0r84EGGqqoa96KIuN0LcM4plmVVp2eJo4GULMzl1cn6hz
Q9Vj9NGT88LIWVmARCBoze9y3MW2KqwD1G0ZUizvL7lAlU4EdRmN3YIBXJv5Fh5i1QtZsLljOpFo
hhzaz+p4Prh1jKevh4GRWTCHCWzOwsZT8DKewkWSHijAL2t7rSeV1V76A2VLeOLBlq0P62z4wHix
gV7HLmD3ST1U+6bFK0YlikDe433TI/cf/cA4hoeejQIkHdN7dhagJghhSVQ7GUf3iEZYzxX1cBRW
4rdRWHSKY8L3VdUKtftkNYY7ZCnQ9z5BdnOVx3uZJSoI1tLyKPrzzMiTEDu9s0GvDv/3I385NF5Z
F6+nmThZW0cPx0HukYY+/mo1iRFbYf314S1dJKwbl60oC23qZV9NGMQmDprQRBoBXzuk1aLFEItU
XtTGLeyaHorizBNjcEs1CWQy7CpGSTAOHRP6FkSHa+7uC2d27Yjwba+15SzzATBHtMVBZvQ4+cek
Y/0VBkOkCBqWRyBHJxiJ6rJLwUvOHxUtPWvxKqywM4g1w1U3JOLw7DJhvVnzICSAMU+YjYyietp8
LMtSqambFlBTTVMbaLiGe6dnvtcxmvElsl5vxW7pp7oTwpeHs1vCjS4uWP6XlBKPGCaLKXKNDnNr
e7Ffq6VVCHlT1dc6zsCAmyWqVTkQ7uJ3XO94gZ+cBRazExpqdK+vM7UBK+9/CckseULnnbxw2Qxy
P0y86Mrmq5cYbSVV1vJVTTdNBi0QFXeYJbPyvDKJnhYBvv36k48qsWOP/ttJY+ptnsZRRZ//8AW/
96DBmzTeAwfnZ5Ta0bHAMLDUnxEAE7iHpigonirJGs38OT1zfLFvWOioIneJXAeXv5tmLAKjS2AU
eaba+eyBRLQ4oc4Y6+8CRes0myjWS431MSE14l7oIOc0NLUxCuTw5xBITG6NEVfVCVRIf3ops5Om
is8mm6mUcWnuCedf6JmUEjeH+yDW8hBbXqTUSkIHQypLnnCUACYUsYh63BNJdZv/qBWVXn79ABHB
4RUC6IQGxPXla6a4638PrfsaWWu8cOHpw/l0eZ7qGZSbhFmrg/7MtOKFl6pwy1GqeBomWUc8C86h
rkNBi2qvzztX6pyYgBLxsiA7yW7oHG6x7tbmQgfRYgbP9SQXFdC7bWzU+eO8ydNUD+vze50az2IN
MWamNsQ7WjWNoFuv7IXn/Z54X9ZEVy9PdtTBL1b/28BffVkhV5cT/VPVOP0V0id/iPu/kwwQ/jLY
shYoFrTw1+HUFkbzIOz3g0+IzhD8X5/7XHQsitP531C1HfXLtl/BzC5UReWKNU1hS6sbRGgdZOgx
iLT47wwxCwaJG3/4mXxK3ZpzoS6QrrHnQU/5x88ClSwH2lg1tB/nQYghAA2NN7QFI7itrI3S19Nm
S/ONFSrL7ciYDNYMDGKrcGgQJpZkdct/rxf1DBl6h3aBlnC3AU6wAzWOrZZ46TGqtmBby3LYaeD5
tG+YD+0n+wjJs/dUq3om3JtIuK4/JWAQR7GlYjxUDEzxWb2yLi0mX1P77nIYaDJwYhLJ1yMh9EC5
QjIhVLu/8RBlBaKFt2enEJBW5DfO4L+JEbD1DVxEUDnyk+vZwZP/m6kvZW5pYOlpaCQZXPn3qxzE
nhTgJVoQ1i6btkhBGYhlxIafYOMd2iRSKsm5s+oc4MAjRwViaaizIyezfUTevFMmGnKK2WpP646M
3zoage2M2B7vghXU+x7v6kmuvc9J8dj6RrkWBjrK3KMwpZeSIEr9uze4tnaiuq7y7Klf+bYatpP+
Yalm9gdGQqvXF+p/WSSDwekzLnvvDbg4amSwcE4lshQ3AfmT67pGAkp6dk7vSc3Jc1GRJTdtISjs
Jpu9/wdlICIGItzxXvcm4T3dH2EDOR1UsCyiNMaE7kCw0RgUfDTQpK/i1rqoaz7hQWPpSCP12zqj
a4qAIY/KCh/N9bSaRar6u8aZUAx8lSPdbBz5YXgMwJDrA83CMr5Xf3iGXiekaEodfiD03NhGTD9L
AX33kp4vdK2fGGslkVE1qU+wD7zzkdLlcBLdIc3G9NCRuIei8k4IQgxM0TiXqV+zoFoWFONYhwpr
ZTg5KL/uVLKps1JnNFKhOrF6qaWiqGsr9J962XDTuCVYMNSKaKTvhyaAUS9zXX7DEMb0K8PUZEio
hp05ZH1MgpDkNpPEXSGk4AWYXue6QZQaX7vt0fpCCOV56dDzJeEdUe62sUyoL6QPfbPVFHtzMQv+
EWhU56mib4P+sgSkm9DgQChMKqM131pM/GT22Hu+DFSwjEAxaC9nrrI6+Jomklo+ItI6FpkUsecY
OUEMnci/fk1cD7GssO+pndUKSKtflHc12lLUHdATJ7immME9a4Q6n05K9mxjlMYVWn/LmGvNppZV
agxjigp0s5hagZLL2s/TrWTIugNe5jYUgHF1KWDNhhWP7pNj6Q62pcKAjPV1EqSTlFuVeKy5+5sX
5yt5roDfry+fn7NXzg0LKwnb0VpPjKmA7PQMIOIMQoxNSsSiUiv3Izett7dUsdrBd3B/5WAoGqrc
qOsqyDSzOivu38xyYSxp/ZyvwtSnYKiYtDB6ATHEYxVVxwCLIIu0dn6sLGOk2ZfF3CN7uAT2rev5
+A395LxCVFHw8KzF4jESdD05VpggXz/C8D6ovtj/GZiyrJL+DuHYI0Vs91oGNodcX7e2MPRIoHXH
GJgBZt0quRsQjb5dW0HRUBsuslosq5YDdQjbIEcHj3tFYgXUXliFw+s1vmAOsc/j0bMHBqMR5+XG
MdMJZ2C/Tmci+S8n+f75TcflF1AHqD3c5FNvF+0uQGGI7GG9B4kq//QnmIJc8lPjb2YhsfQ/+PvN
o6+8RExkheTpMPJYnC7GZuXZbU7HWyVM4UqLbSH3mKSVlYPV5yokuUF2ggNH97gXkkWUX4VOsdGz
0UP5oYPKk8xje22ETwuGeoT/Oo5bv4aX81C6z9iKq0FUITKFgr932F/gf9HEWYYOwgCH+051rLGn
gYE7+bOTB7isAidHTEkEjr4rQqSEtPVRco6SmDcrcGPsYIfqyUAFsL8QNNyruiYIy/v0mxOOsEiU
3KBrPPNEyTuwYCaH7ww2En6E2ISsnHpLTgXn528fLlp6pRHRsbcEqha3HRE3hhgx6Gl5/DqlGgHM
/kEesdbJiAO/PsAU7IXuVzd9trbJZj4n1XoW3skexvjv961d4XK7wx6lNddvrFoegAjYzATn7EzF
yL5grLKnusiJyTUnsKuwe2HWvU4v80qr/3yKnSNScYsi0l+U8w5uaDr/WVgdY33Sg477XOsCi1/e
kE3MH8/NRqsFxwNjCFKdEt8Tacf/Zw0w9rNWsnbtYBXtGKX6mADWhmizHWziyC093MJ8Ez1jnOO0
+z3WhYSpUDp8d7/p+X7LpFwrLMNFPZwkiODSZt5yLpL4Y/ZU1f/gDzeWw9FZnJkt8vdPw8Hmgz9D
Y8sMUQ2qtyoOETME03vC3fsQL52Adv3+T0TZqDyz+ZAlfDliybWCHPta873z+NwcYw2UTkAisjAI
t5mOsm/yGxpbWIIuCc9XlQq2xtf2JekfxSdlGnsPVVwZTdhVi4qsuMBh1FyFoe2gZVw4R+Wo9gub
bbtQMpSvKD+7sbdkjr0qB4NZcf5EyngruBodiwY6QkY++P8eVyNyl0NUZti4BlPbys1QeDT4mJE9
c5Jmu7zIvzspGG5ZrzVoH10pFQ8SdDvOSH5B4s1xlwh0gWMLsVeZQN5kfJ48u4sTSdAkBEKRxA9+
ieqk3Xh5AqKapKvG8b560+K5GMbxbhzVigcVd1JX2xZKY9JesevQq7Fx1I9Rv5n/XFw+as7SGeM6
zWp6yXhv7eA23nLLM00ObqOFTS559rMXIAkU9SwFfJtKXKzUJEbsZNuntit1smUWLxGFTuwfgP27
6MontpKGZ6EvISBUzunwnNa54/9j9rW6n+n3qF4q8nqMfv1THdTXR88PvcTc6GDQFe1sd7EMxZhb
cEDhBk6oxY/F4YwvvTU4dIzxEhmLYmQozzKxXBu0HjTIflnpQhzKjQubuzGe7qXkGEiYsmJAuJwe
UBQiJgqRfrQYPuI3R3xJYDwh2Wl3/+qFvZWZAgDmbON43ojdUdmecBqxfpwj9OZyVZKUp5Axdr8/
pymLF/fXjc1/VLKJAVxO6kR4MzFeW2VgafoDLAHUT0GVYJB4NXFmO5Cxp14kPAeJnjTIpIzWl1Ol
ZPHnCi+SIGyDu0mGi0tRjoQ1QgdjT4bjzn4LCQtD1rzOPUgRKnHIOpfaQmRPhOtaW4lvYHQzwI4b
FydnCIU9CWxft17OOhyz4KebY5E0rLapIAYGsQL2FIq9eer5pAEM3p2U5HUhPh9cUH7YaMIfgKhD
2t6sc/s7aBXPlI8xeq/iXGWS6bc/ONa0MDGxhuzavO0PwG6dkiaFsTTUr0bQ+YeXSE8c8qMkjStG
TnM0CgNSdcdzQWAuxHXB0vzAsvXA3IqiYcV9rPOWcmkNVraxl3bP9h+2hOx4rMybKWyrUzDu68fr
DrodST2dRNIyapMkbkzxpJIicuAkHtfyFvh16AG251Z/45nktoWI9uyjmWp+sqkG7bvyrQI9fXLj
Ct9zQcqi4jzYQld8GoQNj9ZbhrKWIaZVICnecLudNs3mzNtKrPiZ+kH9dfYLFE5zQPi17FkDxYNP
qbQuT7NooCFYyyX/M6UckkVUH7+iyHVdJTii4y6QQaiellzgaDfAOQTqoNNYTqJQV5r6/HcieEEf
p0KfhrJgJZUNMM2epDkw1fYAZNond1anzj2SV8j1y9nNgecSk4gDfguuiPIz1K896DMOiySbGEtH
iMy0sbZeBLY/8DtqBE77XXPIjkDSOqAUCJhxOaGReL9bhI6vb+Cnx8IqGpswdtkuwwGGgJGuHMot
cGy7+4mErISY8lYOoy3U/FpwRYNbHvQ4S3ADLSbjUjTViAsGSyyvjewZVkpZlX20y8EtCHWHudJu
AHyTegcVmJv1JYPCKRuMGMAhCvPQ9hvuFWiGNIyedcZ6I3fW+Lc3gqUgXYU0Qf+2FbmCAkFNZucl
VUsvKFqvcZ8Js6GL+ALTR0HtFH18HNwtyj9nr3MVVe9P136ASZm6fjrOgUNXEZGp9v9rC4jJXFZy
JRFaeJeZ/Ynu4+ZW4WmTJrBHXEPKzPARDDd5wpnYJeTpRR8QPtfo2MGa7spTJ7Z68ni4zqM3iXQ1
/SpYLnVxD95eJaICKjgGSF890MLaiIlLrasGNM6iCt05DUZL/83SMJUHsCDI9FxeJauk7o13eUAl
oKBb7xFNSWysuq1FIVqOllHmSnWg6kMaSgAWSMSVXVfBeoCj0nYOCfbc6pj/Ztha9/iQq3Kbz0vj
peJmfZ30CqM5jad88Tc3hgTUpII7HF3mjjy7hRRtxh4c9WxqKxCyunl42T4NLwQaVj/+B6qIYbrS
67ZM54YamTisg+6iuf5l5qZa/ibXVNcbvcPuNt942RFtQcjXphvLCKDhm5SzIaBgs2H5Ho9o+E8j
CX24A0wTMA2lltgxYJvpZmTc6ZM0GEplJXVs95LJ7O1fZ7qo9Z2rtL1T40O3+VeaLcTuse7k0yKD
Azur1acroYCmwMSQykRridVP5U3/M2qcYtxWumut2r3IJ2Ach8guPN32gSv4GXhIW3sDztfqLU7G
Hcxin3OYBJRYAAmvH+n9F7il4/0kcVlGEseYIONYmJQr3Da+Fwx50cfZdYoDUXDkvbdZgSTSnJz1
eJQDG5UiQOLP2ZKeVx6xrObERUcW0THZkq804S9VUjUjns4YckJhCC7+J0qhz/OOc/+bjHiFOUVQ
Dr83md79fcNegoFMLzuchXN+mxxBDaakxcQdECNfCMbSDv/uP8KmDVl7bAqAK2kPpx3qVznbbUk+
iYx79d+J8tGgpKnyaABAZgtG1dAAX1MPV9yp0nN5NHRuNrvRCoztYgAvz+w3wHb+UaVOmQt27uUZ
143nclERr7dyla6vQDI58dXqnavA8gccBzZcu9BlVP43HO+3jT41pVI7gUPuwPutKrd6ZzUrxrSa
gcNzTfispYU+guDuOkBNx7SaqhA0nPCG1ZSUdque/3mBNXAZ9ZIwjyk8SfgFABl0LPcqtOcD3GXR
lL6v7pT4YUHlmHpGh/NAAEGCuBFCPzCvsRltTQHR7MAUYwydaSQV/zSz4X4tXVeyactZBngsovWH
YBDoBs6a1nzWwoEp/m7gwHbHwoMTB0U5Ti8sPN/xfPRmDfq/2P7L5ETY/d5TWbxTpQm+Gk1MxxDB
Svpp6rSbtmAafGk/dF37NwQLyLUfxiSS0J5wm1zIteReD4qGcOAOr85YdjnHlylQX8KuHmKidWVP
0jBKWlKrR47UeRWfvFb6qHk+5ka8KMWMsQO96Eezrdw6prMtcRw4zmFcjsMlN2g7zEsYlusjJJpj
di/xmJMAV7RnJiEgCpICkUTQx9XHdkBFP5C7TBmortNpkVmq3bBzbtTk6OZIR/Q+d/hwkfCGwwK1
Hef+0mwWwB76OTvkOip7kMmA3/o4JMgWaVurATDhxbTQiSe8dD/LYnuEDjTP3rS4/GOFPsN9BkbW
TC3i9GtGXnJrLip45191ySuHj99e84bBLbhG1ICBqwAz4LOoGcBTME9eS+se7FS5DUu4BPN/Npwk
e6sH26D/ahIS4YwSuJ7sko7M5aH2H8EjjAQPAr1UnxbGUtIKse8VSEzR/RouH8A0c+T7S5Z8QvhR
wmzKl/2KNXz8xL48Wf+qSeWb5x9v0G3To9FSQkkZHq3N6aoIO6asSmxhtLAAf7sWBu6w0eQ8LzgZ
pOwIo1lrs3gNENR+YnckjIYf8MQ4Bv3g+Lf3+U3eXbYM1xd16gini5LIz8ZLFMQ34fshQVwKr3q5
W8D6IA4N6NArmtzAuBkaEC8Kr/tdPYOvu7ik95pX39GzbXD5m9tdhCEqj0gqvowspjpIJEvc3mLs
JQxJuvle5e81YMOzFW/GROLfCL9BwHStIH4K95Zo0ZZb0RR94ZDnGOnTW5YgBA56RoYkU60NGe97
BQ4ZTWdFwy2M1mSdEyHdEsQn6HebbAWGYNma/UtwdMpUyPtIB+xsRgSC+vPGKO1gfBV98jnkN1kb
TgvX3/Ed3MvxdcBPGNOLQOc9+BO9tdgV2PzE0pbIukodjNSIEHTJYMzeFNemgzVUfXr2C5AbJzxV
jCg46a+8M2HU5iIeBDutrUcbXj6xQpCKLIAivXWtkmO4qNFmTwIN3yFF0f+OSGY32oCckmDeAfF5
hQp39f7WNKsqu3GB/kPZCH21f16YEzEr3oNotXPyGhjk6BGgkZRO6ggrCdJZ/aBP1KaH16n7kAIQ
q9jvOeH9OPrMh0fBbf/YvW+Url2Y47M4qvDMflmdJo63H8InyfDQbrZsJmia05il1LKsqke2ZfJM
laGRZQKTuyRfWu2iN2lgSNUu0wLm6dhVD7xL5WJY1lbY2AcJHTJsliAG2VKA6/BXZpVTLoQnspmg
8Qt49CQN5L2jzxXv6owRqDB9jxtxwwj5UBj0PTN0zd6KrSJmZmekDx3NV5CKu1Xcg3+rXGkkm87U
TZXT7yFD9GR/UIPtrWSwi9eWs8pnoq9tD3hysOM6EXN+/ls4hkmG4QB5rhf7MHDLQ9UJcmjDi4ga
3klP9ZoynaaDgp0iQiADhPrqXvp9jVZTD8/f3Ikn5Mmzvj5gZOur7t7cXsEWH44kRwL0MKPpJeU5
1lw1jxhve37xSMZnd9s9v6Mfkwjv9skU2wOCfN0LWm6oDborTGxUJRpJ3oQ1OgIR3sU+T5/CZzTe
BWBmn6rN1314e8jAD3UIyCl/kLQLzxs8JKfXl2Gy00h1yRkClhnlm/4Sf0nGaIyEuw4TRTk1VV09
UaeDkKdiC5PKZQu5T7L+mDGiqJ1524AU3n5ibDc/iVkVHdkn5gNe6koxCLeXeiFQmniCrIsSqjtv
V5A6tdFRaxXDVTyl2/iE+OzVk29lej4ITx2CR3AlbGHc+cptW2LgqASIb0BevcgBDct/GZ3pOz0V
idMBQBXp1zEzo6EqUMP7XC66mUXtQpOn7OF/zH10xg3D1j4b1rAbYws3AqcpscpmJaZnnOr7Kn8b
MA/vYP8fddanbUDMSuh0vr6c48Oa/N+Fz8n4QADkSnaAIoweRmhw3/WbiS4nMunmSQqJPK4nBRWj
Bqnb2WWuBtEUrR1RImLwQbjd+eFzi1GpZk0HWrbV6x9bvJGSY/6e5fAC67vWgFrcz4+il8kj+khv
qZQzZXMv7zxzB22WuO4POtd5hU2G/UvXJPLDBnmJOhmDaCc1cC7na3vQEEX+l2+D3u2p2RCZmhYE
3v82/ClT3oV/jUxa5swLgmZLSdjRBkxe9Nq7SNKhvgqUbp8PdssFkR1hkLshyI3ZMlyu1r4kD++4
RjwGzFi5/MGQqitfIrrOMf4gHttPT4VFe8hwvvJAyaPGE29PxyDC4oNtg5KKKUF+5P6XYbQrlKpe
ISZvdL1J+GpJdoqzzkFvpaS25uM96NWtwP+dZMfndhkjYNyb/XJXLhdIcNZU2mm2dzBv6pLL4z1u
P/MDbkauPuM5PZhmmEZxvFH0GLFNyd/ZXv7kojpA2EnYYAEdZLCdI8ZcNzNB66GmFkSxGBpSaVfY
4pCvpJcOio6JfeRybNs1NhTH7ToAPN3fheJubXlekpbjIcHedLKDdxoxcwZ8rb2u7n7qCy9sp/TT
5ps4K57H2c5FMzamVI2tDHueOfO+yP1XW2qJAtBMEFGysickKdyeYtMA8hJxsrMT3nnyFNe9iTkZ
8lEuUqjhyc7VHcrRHWm/2CSHdsoSACStLBCpAJhj7VYLmuBvBHD6D5dlW3qLsMzj5RWfwjhGsEaJ
xyQOMB4ZYETL7UpmO9STEZywFXuT63ufRmD8q7+gOqgAEO7mkXesJ2i/jMhodRG/iCypcLdi/yd4
UwLMOYRWvKIwocXqrAqyl1gFT+uiRU+siapvZI9R0+oecln4EnXQ1fnoiTZXoSs18LHZPjFtGEm9
H8qA0t2yPXbXLnzUC5FmPnpA3JzlLfr8zktyNuI97NYbUyaXBFMHdG9u3Cz5yJ4LxFK90O+L1E1n
fuuXa4Ur6A0aLKTseF7bxnv1f5E9NDHvIchk6XDHMoEfJcDli5wyCu1fB39V57U/+f/GCWoENvQb
O4E/jEYFM+xV399zSz4vXwszlHHDr0jiRHITxFmhljBm1IvnVpod6xPYUcLnBjxT6aO70HEjSWDk
AlPPAmZZet6o0EfC1ZRV3qWQda3jWv/RE63E9WZebi0ielkm03C96W8KB0CpaHd2wxBxgkZ1lRpG
WGy1K6ZxQ5y/f5hJY/jw3t8yuZ4ZeNLMsRleq5pXOguB3wSWACWiSP2XuM14U5+J1XkvQfZZqOCo
d324JZ6UY0Rz4yrpqG2+JXemAS1vh44Okzlkvm6gIIkEWMXa3avS2nxZwLO6kPKuogYLlZBaz6VZ
JWOaueWR7bZDEBcvrEcU6Ci/Uv/mlY8mBDvAnmDNSmuKe50G29gGRbh8RnKR3jGQBfG7V57k0kzR
eEXYrnzyP8mSXzJanuqrlhLiXzi1Msyjtrhqq/NNRRQUHpAYvcIfyGFscHTV/j+58+72IqGvFxAI
DdHLTtqdn57TAh6XkSGfj6xtl0HKa+cQ303c4YsbRIDqlQRUTN8DfuAIEXQ76jGuzOKzHfJCkCGx
XjXU5rzfCqJXfl5akWJdSzSiVMmkD4Dm/aobHgNjqZ85D9EP7tB0IQZEiB0HI0hFXO5z0fJ2uQ8u
KYztEqN/j+zxv8S9YAKOvMvjkQ8XdRDBtdXwt0yyyHerec6yz0drCzSl4m5r/a9csN4VPGrIdBav
7HjEVSKeWEeAHXNK+3daiFp4clh0biAbAVaXDukkUa2Er6Z99JZ97yW2ceZfqX08cQcT88tNntyj
ENOTLeo8ciBFbbsXybTMUIwOY4Uf83vhVEzHGgsXu2GOpKGhCMxcormFQA8xPQ9t9StaI/n2gcRI
7Ft83JU8gNqh4vsXC4dQBlwbisoVxDd48ChRAjS4mm+HbA6YZe3cUBUhp29xEv9GLHUhMxix4qtm
btayvLGhCDaf84/3mfM0nllP4/A61F5IGwkgyLKJm4ZdsliPKTejTAdu7Xr/x4LfjTq19acVOxYo
uKiMXl0Z2rc23Jy+Q/6dUNtpsWxtk8oXXMc0lXRrfeAV/q9iRBjeBlpNdXu5lZtop8MrRtXRx+2O
opKawbLNq3gnmeYF2i+rMhh9WvJOElZmHYTOx0n0dd3fjlIrVDAtoMcIQtVMpXM9sngmtl0KuMeE
GKijy1Xnet0rnbn41etvAr4qpq/xfSCjUPN2v5L2nyrPcYX8OdMzM/9bA5QjnBI+jeQFVq7mzqpz
J8Xb8VXWOSrqEdfogorp8beNxQvwWZWFYiA14t/0swrEaVDSSbnJjkj0KeCla34lH2IdoVvb0SRg
oMlX/jfLwyOKAhvN1+vjD/G5hZ1/8EjnIPl60wPgaQyKiruXP588sMF5mXgneLYynHtzg5E84kqG
gnJ1h/KAEgms7PahXxF356MSqiLSMuZQArIiOCUC2PrEZkWajSYtoHrWi0uBFcT/aNoPCHyvxu3E
gfw9f4ufEUlusID8XhQYf/JCsPQbCmMWySiJkRJkydP1gMflkF8ac9kzdZsuLHL9Z+Tt8Ar/akqI
ZJajsRsRV+f9BwRk1gW+SZqRpgvS35Ak2gy0WTbUzanzvcCSRbTu0pbJhSNXp/8mh9epdTRav1CC
pgqnRMSTDhcHPmXjOxciMY05i5HHwaLOVcUpAf112Wrox5tMa4WLO/4pNGPht58JHvzTGxzx4zvz
mGF0BFV7TMUhNJ7uh9Jrn+0LB+47j/qsKh9/8IAik0oF5hLcurFLKp1jvwrqChzpmqtvuRo9wopG
ExPgQ79nW/zqlfsRdajZ32KsUe3Yjd7HT2sHEvjM3vPNL0CnKoa24p87FXtJ6PhJ0NABcr7He32B
MAbsES0n0wxSUa7/PD/Iul03QEE0+CsyAvDrWZyf4YBUNUrQZltV2gTD2+G1Ahss2D1X3Zk+QhYq
rvOzEOTLpzhWgStgmTsuZvjnKydlbC33qIcqLeAUA5m9ECrGc9SpBqFXDlCj5pzxShw1O7DzVZXu
ea3hNeNzm8aN4uczCQ4ymzW9dckkrxQxwck0gSoQ0z1Zi3h+1W3cwMe5TJXrpYnHHvRC2pCR/Nvp
q24HWtYhLtFTsmCFFJpb2jKeDKhq2N4aB1yzkNLHBbOrUXoqP5CJhmU8OEfSVBeoJ3U5R96ibXAQ
Og7YHocwkpSIoBooQoF7zXy2/BRSjbSoMIkahHErXodglYk6oICPRrmoIBRtcGMZylfWV3ZpcPoW
4y+Y/UJ9UrCwoXt08QySizl5N6wE8V22EVE3UUOq9EqYh7JNyHvcZqFIzRf1l20z5+RXahkmkp0j
t4tZHtLrgZ3R6MgM/5SeVlOo6tyGmDUu4qy7HMpWOH+agZdj2SP4Hq10f8QB/gIhnoMG+NXCWGQI
dqET6Xwahk3DiXj9MmfvB/nY6/UToHZR+6MurkDJitdMg6zh0EQnV28b3Ej9+eHQZn9e6iaoahYC
UuEXav12X0bTO+5uQbxVMkOECAysQvvjp00/AvxEnKHAI1tP3FBioJXzdnKm55nRTpHMVVty46Dg
H6iWnpuXRLt/PAHy9wdozVjP9Bz/Dxkdse1ei1uIb/ZC5XJ9Fj3aTki7m9BAiY3ZQPn5fVoqShbt
o2VKQ+pD7YP+8Yb+dD1GBCKRz1igUDlzVgCroUYqanIJWGI/7QUVl+dME7mTKBBHioz9Q2s55ZNt
rbClodXu2PlEbqI5uP6OIqNgJbKSgPJuDWQJE1UYax6N11x7cXi7Fh65DGSrBfKG+oPYdyV1S+yP
s3fICq0sUk6kPQmWZG9AaoK0uYc/0Zq4CIlvzi/3UqvWReqRHw56GUj0HN7Vz1/D68jI3iAiKccU
LWxFJBbOCm6DzIh5Nzw3a/8rZ195r+C/09cF7ypz7I6Lf8yBYiTXkfY8QfLJKJRstduElZ9Jy4b2
5fhaGGUH3X28VdpmEC/ea8o/9szltGykbOp4pZjPCCQyQ/r7rdC2hOJpSV4GGe/wpTg+0BRtZZ9t
YT2oqEU02fTXyGocPYhn1KxQTl6C3E6pVNzY9BFcdQ5mOnkoVT6lCYw4C/cFVJaajyUm6BXsEfs+
CKC0EWMj4Pd1IKRl47c59UZh4WnIEibmlZNruAF7qzr2GQHQKrhbGPLgRfDImQ+7uE0I5r9qAcKM
ZTjbU2ys3wYzJ1BaS0RFEtz0Vejk4VnI0IMwMnsiF5K9DsBcbDPkyAGtEh/khI8JMgMsjkWxbKT1
DCAhKJe6KtZJ6OuWVUjyfMczFnGFk4/HAUfq/ZP55MfNT/z7UNvueQHLFjn3lvw6y2UhdrzWXnMF
tuC4HrcUCyIRpVc65zkDSXcGTupYYyV8pYa3d9q/AZ63bhPC6M0AEz+py6JDINxaJkZEgD7woj0T
HExW2L/8jEMrKICOngVOM9zb05yW0aRu3cdOoCAenduCoNu8mvVrFJkGoA1YkfR58vs8p+VD7ve+
EpiTEMmCDSnF0EPRYw+pADdbaktlzOn3ZcF+PATh2Ooi+TnmEZyBTTKHfWEdqq0UQKiz3/9tVAtg
M/XR4WD7twBU+2CpyYeOxx1DvpUIiTMQay0GXlcmYGZ440yQXKlZ3nYulUUBYwuektoTXQ6hKZod
XDRmfUGBB42QYoN9cIFLh9rmoluSy2sMiqYAr38A9fvYY4XsCesMMyqTChfNsTlFxbsEuOF2GF02
Xiux61E9Wj5ZFvKBrQRWt4JfxVbEYfVbl1armC/2r0Jg1g9Iqs6t8/EovNdlBckLINKMJ4CqeODh
5+IOSlS5m/XVyKJA/yLG2nzjTvafM1qMbtS6qFdCiTnq/2xGMsl9BgdoJwyJsKpIdO6arJePBfq5
79fMxVxWFlXwu8OzVulDVPcCVt9Rdmpc9J0S9wa0Mp3y5RVds/+/KEX+i38YFDHFugeskUpoHvZz
SKj5to6DEmmZjR1U/G19msm8OwkpuspHEpBlQqpvywjooUKOrmOFHe+4dzCuAfKuTEC9Qzxl8rLm
ND8O1yjJ6v6JD1HNoIwAyjZEr23UWcKHQ4ZLQpDea+rtdqb9UtlvIfCyGQNu8/EbQ3MzggmuDPJy
SaCHVpvbNYOI900mBiDkeEk/J7Z7yAVh+mLpwa8C1ZcjHKtidnH09Qs2bWGewQKLoniEYuaqX5Pf
2Gn/InVVIXhn3sOuAT5hjOkbN3mDV+8+wi1arvQlbrOt2Q3RkTqTawc202BdpKH1CIPwMS8kicpc
0OYCUQt6iD1bg8TYdDo1Gv6YkxwP5y3+DMrzokFRwm3/8vLMF0iWqukUYN4sIYPjnzR3j9SK/W1w
LW/L06DS7EK+DyrDYY8e05VdmrtMYQMxzuuS0tOUuW7XDt4z2wZrSukMv5Wb780dRWXJ2Fq3K5sI
mrmQ6TmQUWUQtDd4N+uxl2j9GQHCkNc+02kZF/9k/6bp5ALwUfNH1dSUipRbEqoZhnjHQUdc7HAk
IY1N6uGN+Yd/KddiLkqsA7XEcUGRGDuGOygvL08ktGf2MPxXmyR+CkAsZP/QqmXIdG5+Vmk3bmHh
XnZikBPyVXugTEBI6l4UJPISafPdpOLzPD6wdKbcNwXvuYZP++QLDMfrXsUFpRoAXsiZo9U/8qLX
X7unnaC76n/DKj11s3+b2xsse2/ifwTDqEjSwzm5gYj4JiIFkfoU3lppQvsv2UxWd7EBC76GsDxY
6rY31qrrHGYHsQa2hV8ed06ts42/dwFjXh1oqPtyg8TLwTzu/Wja+zp1YPO0g4iQjLPJPNNYo4oK
7usUdhqNQYhrMrRPg2FNXuSoeShiG0L3WHFsn96PyWjra5BT07moqOZRA1cK7fGTqxN+DR2rceti
2LkPJ7R5VP/RjKAUzjHjTi9uv+ciH4jWqcGg1jBe8wvdq7O+xC9Ez0Mxbn3goPAwTpoK5pRMkoWt
haAhwdWEOh89IQaUZPiu3WezGyUWGy6+2UtyFV7PvIjfEurhg+sP/LTQXGHoZq6GR7ftI3s/7SYV
xQhwguS+F4wpblnpEzn7pnnF120zLLRwZW/dtCRJg3vPQo55glMEE0yryP6aVyoL+hKEJr7tUN6/
4ag0iUcxCJ/mz6wZf5EcGJmqpizE8Gv/jsMoBQdjZ8aoIZfyXaspH8hZO37sji+ENYcg5vA9Zw6g
6L0rQK7nVNtlkXTgWxek7vGl5WRNFKWXIL1f4kzCo6vyjJmvVFYjuFsQJ0GcRDSd1D/TtHexj67T
i2jrln5ZUrwdCnmwpFLo6yTHSMsbzBhBBCxCCE8RPNDepEFSsyolwpnK1xa3sAvPrPKUAbySXgPd
9P7FHRtRx9xkJ22KPBImnBT03D+7ia4/2QwObkVp2f3xnxGimm2ro3a6DQpVw6/FLgZrsmYB6fQC
eyy9dvr98HRO7QYYOzryTn0hcIJF5bfvz/7dBYneZxHTx/xp3/GDLUy6MUQH1Tv6NR1LNG53gVYf
OiqO28+oTfN2IhaJStlsTPmKRz2gpyaSASJ1ZaCa8z0vtpe9s5W1cuMjbLp5b/JisxAEiaNGzJ/F
47wOzbUp0jFNCXSrB1qG73hTsTDYCkUeAJA5DZiIBwk56vS5AUarx2Bn1faZ7BalkY3rqxznr3/G
jMP/aCjT5Alyv78CubZRNRPQRfo2x4Ebwp5+snXrODPttn04b3YMWdpcE4x2oiysQzr6kbP7gTul
z0dB0sDDosD2W9KC9oN0YVGaUelbgKajZEw0H0afXWB3EziJ1qPptE4Kdl04IJE6oLGKyUkY1PQU
JcNDupK9IiJ/7+0b9lNLCix8xWKm55KDzDZRz2DslOtqElNlLNDeTa9xAulqsrqi0ghv/5ZtB8KZ
Z0NsALJA6Af803Ysvh28AShNo5lFR7jRo+NGrvNimHdinBleE+bCxHYZLlu0FrP6GFOBxzivy86w
n1CELvJI45tbaIQZi5+k1oaXxw5FcZAKLXDPzfwfUSB8BknxoXwKFUl61NhqtWUXxwQf3V4dD45i
DCT5xiahkAMtPhFxHIMSa0vApg6UtjRZ9z7w7URa2oNSQLZyabDt6+5Pn1g+QD2Q20lm27tnWYM8
3fFmojYqsqFtWfyeGtm92hknhIw7Wbwe8KLdFxU/znCj1F6llNRZ4bDxpmoz7BkmxadI1kIHukjl
tVOnGgaU9+f0rmrCtZZT7/Ix3dyIrHIy/3ywUC3txS+V+HJ9dnh6uFnraKe+ZFHjeMptnOPWWqeL
csBxHp5bbafio/1ORpZYDAEhscrLRtnRdUtS0ntIOPsqgWjnylPoEXx//IRQ/W3m99cuorzSxv7G
tEqu5wjaQ+oJCQ8dwl9q42GmHdzEczakWn3HaXVyiIz+ZimDYbQ59GYxWBQFZYVpfl7PIdu9WhYE
rCuLawWKLa+6BgZDTEi2i179j3Zwv2WlHHlr7RPM317fQEJJhS07cgWHfEvDaoU3uoOoyqWlJdal
ospFzR0SJNY4P0gZ5bGYtklcpUeOgQJJGXVEkD+/jokWpUNVVk/fJ6Zf42CQm77asqwftMBc1N9g
5uAyqszuRd6H2YDZNylNORZKSEPF3YXhCN4AM7d3dnSNE96TGlqoqMQwM0jvOCM888uIKHs/U/87
vIJL5aMmzo+ye1lzJwvaGaq4pjglPlP/LRt2qCVynulBCRwsu7tM2RiGXT/Nn0Xj3DHTKVhKz+Bq
yzQ8L+SD2cP2OIESyeYQ/af6+EJSUrhdvL06GdgbfDVh1CeYisDDlMpQnYQW7UeDm7kXD/0Zk1ev
tmar4PlAGVrPLt2cswmM6PCfxCuur/NNW0rgMR7rFJu/s+M24oJPwhth4aN2wBcZQfOVfO/Y9eGo
Ug9AKOln0A5Nm/wbJOzetR/v+oovtQLLH+EhuDNx9HZKP2j/thOfmkTCPANZBWnVf9hdb2smGrcw
EjnIRWW6EI5lSOiJLb+yz2f34BxbJb6QhSIG4VzBTdwYbttyd+AMPNRwTh7zAfs8O7Kc6al3Eff5
Q4DlomdWt/IHIRD2LpxFKpwVnCiuB/wTM7t8g0qgW1WzQtiKf/ONGl34Z043WoQVXL9Pks6JT0ls
zmHO0+9toB7zD+Yt7jALGIdcSjl6jkgw8nSOSg/yyrfMYIHoz9y+4Ars7RuZCVNQ7934ObboTrPC
NDqLWEv1RjjksjH5R9kNre8rXIbWkkvnXlo98f4fNCuljOxVvW2qs24BW9c7zg29tmTf2SZS6wno
HYK7Oy87e0W5LHR3INrzcZrp+czQCRcn8a7ML+784JoUFoSmUPD97302rzbUIWaqUGbjZloHw0BF
NZ6yVGIERRsNp2mOxWT/y7wUNVTaH+LeXv6kxPn616p7uy38O5J6IMgR6IVEw15s+Sj9Yp9vt8cS
vLrruftQyJryro/bTnt6H+hlmSJVd3HlAn+eagHm7aa6+1ue3PZWlXHWzIGVItNTx1U1Xt1RtY+s
PzTPKL5gkYzXmat5XYc3lBdjM9BInaIANAlp2VyaGpf/byo2l/UFHZBul0vVsYJ0i8To26miD7Mo
OuVrXNJDJtyVx88zx7qksejJx2hFBvI1yVY6fU/U+tfkKyCC5ogpG6K6/wiaCXoTQbcxHoN4MEf1
hc4/eA4ai9UV2wIws7jBEtQG7t8VWupfmN4KiMo02YtP5OHxwUdShalGiSf/eZtxGVjwK4k352kS
RREZD8mExHz9f+3KQsPruRLL3Qdbn4+qLYUOgYxvo7e+TSyKeThW1fhdyJSu0mhY+pgcxoU1LhKn
JlyuJ1KmmNYk5VAQrBRnvmH3yB9vKOzMwRhu9PmD5DrzIqORxOLWVh6xfqXSnquCTJswdJsi3QKb
khP2mH1QCEsRwhd8ShTEZhCsZ56BsOgkADh+l98Dk6HzgijhkN2AG/OcubcH4d2hQ6PpedyQswlH
UuGqZfhw3sZlrgfkxBfrA6uVI4mratijTx/uvbjA3QQcCRMwKistMrg9Jt0DdKZjnCWIif/HEgWr
EqaeeJgsmsRUNynHWLTb2f3pAEy5CoYTacT4a3yEagaJW2UX7KRAKZOSjECrnysDXnMtu1NeJ95W
2Z7HmWH4b350SWKRLurJNljlD19l9YimPW/cqQ3Byi8PEUDYZBrdzsVKw4suEy0wCBA/J5TZTstK
41PIz+jNkEH1ymj6wEKVI/lDLtobymF3OQDSAPsL5+pH/PlStEH4hG7HoDXR+dWyqTyIG3AKkpw1
ZYG64m2GltICsor7yjDjSaxahLgxHlkquzh5pm5wUQq0tdQmzqIV63L8NdQDOK8hvFXzjVEuQt6O
wTc2DjcXIZcc03gy9H8pCsbnkxkZDk+9rxbGKvxL6NNdAyoAtEE5RTnIym5vkJycoVohnjkcwMzS
E3xS/+cWfbCDtHs4lPPW5DaAQAc0L9H//qPQTmwxbKCNn8inKsGlyeCBQaplOqrf5aW40L9f4P0r
I4ch4FbY2SMX2AUXrCHnOMjcI5SjxBp+fL+BMfCsPoEuAoQvr8y629RTEQZYvyClVOyndb+VSR0Q
Q9N9+R0q5UT9eLxfFZ/kKzpwy5cVitdw4W8Y0mB7KZQO7a58Ee+NdQXcCqxdmgIFDs9gH53N+8oy
GQPCL297yFoo8sprBSaH18ZAqwaSd0X0sPegK5h/TCsfhKsUh7lXv+IOXKpA2IsXb1YzNPvejB4e
PjrAwEeWWrC4xbMzoNF+8pu5t70BrU/0ro0lQ9MMVwEXfB6NvCZpcTobQAogYqr+ONkhJCgB3uv5
QqXXk8gF8W+B57/fKd+Zd0Fezkq/kbjPKs5VwSL8Dw+a0uTIwfKq0mpL1zpR57+sW9A0yPOiCWRO
auZCEJSk+teu7K7tUiK1ehD9+6/wcP9VKnmmwl1jI5mZSz6oI1TbmZ5W3NvnFjM1OEZJ+GTKwkWq
nSThsghSSZaHe+bijRLbsuJMicpCZz0XzZpaYu1EIE48jQhjXhx1gvNcXnUpOotTCK/d3Af4pvHD
cqvP3J2IlG7rqhHPNZ3Gi2Nif1DC8qY7CFaR+lqAGI1Vva1/G1MMuhxVtiOt1W5yQ+2O1szF3rP8
fGFHdn001B7Di8ag5A0HNL2skrYfCw9HIX+XBxMC2KhQ9OAmB1+zitnYurQm8m7+RtvIhbmzoU/e
snnnQ8CsQol3eyu9+l8yOqibbFMtqvMGfpyyrL+yvoFSH2pJstzXJVyIZ/YoTHd+KtgtZB334TbQ
VlvqHNJCekQC0GEr2yBhWWDaW40vPw8sjzwrt+jBZE7RgK94LLHbTm0sYJUgHNCXSDdYMz8dM6Np
WiehUmtwxsJZWoS8TY6MTgB1tnSdQ0iCZvpRslFOh8WsRUenaiglCCiS0ku0GasXh14e38UxfMmQ
8N2dGKGtcnFSTJrRK1tLTjAsuAx2mmxsNp1YjadTuy1l21TeA1NNjBfXh0iBBH5uf+joUlKYpmVS
uPEQAUhHW+WOVou/yn6aKHhUiwW+l3UHzsTWMlgO0joB/Lk0jTq+7tu+GIk0mHx9jmOog/uks0rQ
lB3jg7tB2ClaDDtkwheE8lSBd/Uirm70xctb+akJAXMez4Pgd+BnX8QzGqYduSkNIuxl9vzxNo04
EJTwKnyBqAXVsupedu2FcDtWGojrI8BY9z9uKaB8qNZ3GFso6GfmmrU1mGydLuWTGT/8yfGHLzLV
j/9l62H26ETEOwa81M0YWctdzQL2ROEbEXKR3YYL2u2TODUsgnJt67xAfifzfa/W1vfmq90pnyCR
zQx374qIcZWcO459xGSv0uwTnea7U4eHvqHt/xNk6lQA5s0f8f06R9PPZNBbrSNkmLbKc57p6/8c
GQRgKtL9G2QElWcGCLDUIf+TQ2vKl4oW8ShPcVeVxfAAjtQGKYRjf2CZMDKkgY5+0huvECAzKX0W
FGzRrKEu1UEt7NO2OmB9oHE9DI94XxXIzzU46HGxJHw0ZtefZB5oT5Gk2cRG1emVZshK0B0mf2Um
jM5fo4ZGQIweutLdU6IfzI9W50aoksyTb18rW9dhkglGpGOnigGAoxqbhArtQ/P5pgJwSeI5Li0i
RGtGyGm53Q2P3WG9ajr4faZPoBRvZuQTF4kgGTmsKRqEFTRH9Hd80m5OvYkPoRETYURJe556amMF
ostrYDDWFxUk6C+M1DBkH2xJuAmnKH2ciXvkUCNfQNqNkTVdKQt/gj9mC/hMlFN5SdJAE3mwBc/g
zt3TbiBKXAbe8fQJONWL22jOv53XTcQOwOG6/5YznejU33z16M7rbpFHap7gUow0mqlaj6TmuDL6
Y1dIdA+3gR3oKij2dVlZXCx0uQxCKstbH/Ozz+k8UDJd+8ieHLc4NfsaJQvIeYABRTCljsiHdrWG
gk257XO36eFuTwQyNPJpl/ONYZzdEd+cv/ITDMjDSQSzkJrJqgaO+Iki8hQ/boJYqyRwOzIQMtoU
y/+zkh4aqwFijuQsjYAISMN2XxuAOzJFIFMz2GB/3RfzLTEUJ7eR8tns98y02cqmnbqKCGIroLR5
g3KaFC7IVCegJpoaC9rUbxNNOWTY15F/m/TRY85AFyCbdgserRl9DIkaBi4L9h59KuaUJM6oGxG/
8i30qm4+YfxKFpTxSUbZPmcHEW57Hgb6rxhv//GFRen3O9NLar8U/OB/Gahg0bMZFQioOFfsbjB6
tzaHd/BiSiCUiZ4/vkg1IHzmFFMdKhZ7dVcEiuar/q45YqfsM932QZWA6ig2VLUJ2FJT8TB6dyyS
8EWmjB2wynNktEWPHfu8CTHffb5I2H12KXLsSTCmuVUAXG5yny3tROXuUtmT7v7AG6BAg4zp2xrD
0Vg3Rh2SVFtLiifZnfguKlIq66HGRHJ8eaERDpDoSo4TklT7TJNBKOzGZ5TdKDWsMVW/akKBGAzk
J5XW6euyuSZVWItx8IedWqfQwz0e1nkCLlRD1D7KFdppE4nz/E5vNGLHjl57C/dh6os6vNw/nuuw
C9B3FWHbKgm8SaBmcuIVaBdUxf6hdtfG94+AQ+VPk9++KjMBmempFeX9ILrdTbaiIxCjYxdEHUO+
YA3lVsVpMKprwbto+tj7+Vs+Xi9IAd2l8OyHfmBek12XaNYscUFTUpx9Ixdjob8WhCRSUpaJi0fG
eXkwyrxZrtNtEWrDPSZgGu4jooqGMq7Vd9mxzAcYqpEP8dtwfzm5b8+dUIfksBQ90zQzCQPCmjDy
124lL/tcc0moU166RdSVzUW/YKWHsnmpHd+iTfRLKBqHPtU7VSbv0EqqdATCzYD2QBmAd5HTIEBr
7J5IDrUCRWZkUpFqixI+6Gq1KsTMFRH7YAnZAJfmJDDT+xHZiRRXKuUjHIKM60ENlzlqO5lbLb31
fkDuGlA1rfHyXB0ypGCw1VZq7DCaWq23V/ipmVVnzuyc+DYbprknLh7x3gi5+YxmX+L1bcJWflQE
e7wI6COm/vY7NTBE+2zqbRuGU/v84uGFK5ltNpGKx6PNbea8oHB5HI+zdyvCpcwRAAEqgUV+0KDS
5TNsLsMnbyqTHno+DkGBKHTYQqNQ4ef8JopleyvdijoQCLrTk2ofJL0Wk/3UzaVY/nYXXHHLgdxB
9iFTlqBy3YS1/Q5Rbdv7JzFfTCJ+BRtxXLwgDMZOhykudBlKVVXGFlzZMxqRuMddGZirk6S8L1jR
Cw7Wo8Peemd8H8mE2TYzar1jVwYIHNvdmSetfysi2hb//YFaBz4zkQsk4dUuRPDhEcDprDE7Xjmc
8SuxqBxsRM56Wt6ua8m1PLj2+adzhluxgW6y1H1TrSWD9nv4M4PsL48uS6QKrvA3dAkD75+bHp6S
t+7bLEIthahsO7H7arY+yoVMamzVNultb5YNjXNMJQKqYu+G+SNJq9hdjCzxYGrc1sacOGuEuPnq
QeZKZ5P4INEopZMbroJsk7OJ26prQ/v7xU5dY4+EtGlA8qoQCWLEV8wSo56/AgxTKaOM3zfiKi+0
aeIWDrzE3C/wr4atGJKibAmiRPlL9Dt2D/8SkvKY5NMNmT7aHkCC2Zy6LdyLC61UW+8dsNJ1xxhp
Chhf6QzA+P2oqKaWP8h28n6vWPfj/ay8jyuhHfI335t7Aoxsnt8OpCgji/FRUEpNvitBjQoRtZk2
cptO/fqEJRhFiwxkGO3LlrZnP/VCdxtihYPbAb0s/oyom3t8x5lnEJPWWoJk3gYb6uBkyrH+GQfb
UfD2T4NZWvigMeZt771xPZSmcjM9uC2mCUNcMfX7d4bBqpQHZBREqiQRuZSGdRZs8BZBv9dhTpLw
cjOt5wg8m3ciQjOr+PWiScAEenJaAAxKcqiDhaPxakbY49uc9aYAON6HFNNiQbXzwv7DmAbUpbBR
2lyPha5frCXYPSQo0D0hZq4Nyz/Q4ytL/C7JeDdGBdmpNu8Vje0FlIQSPf1FLSBusP/yd1SyIp9Y
VlTgWt9jSRvfom9cSo9mTABVG0ve0wbE26CJwU4on25TTREQ8/ahmnMkWDq8/FNmnYoQv1sgQYGM
fjeZQlaLRvdjliFeySHGTIZ3wuONqyheIgy1bg90bR1c/1kUOFPgommq4hx1e7uS7QnsvrH6VGXF
LF0XYNrUcNBtKt4q36vVzMxnW/pOAnMkNu9HHzFes6mG7v2QyB9yQJrOc6XVIFjEoTGvNRQBEdaM
aPcqCyGvtEwPvULXAmRi/D3y/2EpVWPc0cl/dldEulb8xWY9GSGY4fjgEOnu2sxIkvWAs5NUrYTH
fqoxieQ+4P0tRR7pIUZopWsvkMZ6I2C0Vh43MZMVAmFyDxiOy+mduJBxeiR8brJzSF/xEadhLm9E
AjmbcQ1c9WNxF4X0eaQCk94y25+rm+//x0bLa8nXOaUgmIeM+/YA6kPSeheVpkajD+fDUSbnnfMR
J5goC4VVKNc7W+x+TWQ0cNQpMZDdaGhfqzHh1yHnsyXby+PboyD0BhqmuoyTeTGjxL5Q58CJQxW4
2O2ftNXkfoWtXcbdVk7Vddu9SW7j+sB48G3eAe4/jWGFTZbZh00zOELQutxc28jFRwhAil9DuFeI
mcq74F22Lbv54F/JaA4gZ6iwFPqhgtYaTb3NjkpJ1hhWzDQFb+SYvIFOWmd4wUO5EbziJOGVIK0u
7B2JsMZ2Culovfvq9Tf4s9VjkQC1kxfhYqAAy6BZCGZ7MJ5G2ZZbzBEZkFh5BWOeH9uogutwn6SP
M6DUqZuw5eTJigz6jQPQ4jCi9J/Yr344LnXTq8iALBm8+kQIYwt8qojUNWPcl2BQi2iTubFpWB0g
Ifg2mXn2hBCUtEpjoqKDsTISaOWgCJAIXHReDYEdH2LSA7beDCfifNyQVZPvMJIBfS3X+XRK1ZRl
8dWqCVf8P5LOFTgQdSUulMpFYPYJhVccAKklkrD1wOcc+CQwMleazKY3N6WLvzeJBaKbEs38rjE1
57MreJm3Gitj3Sw61Ckxg3s5qY/GL3xeBbCyNkDE0PGv9dR6GVh1E2tGKGSIMoZGQEW3fdsQA0Ju
GLo6CBuZDfeMJojJ3n4JeKtRyFeqZpFCJV/V3Cnuh7GsHbiutcYLvzqrwF1e4sDQOzWwer6c4XCo
Mmp3bpl8wgZm8NT5mxIbFcpzYd0LVy22k5VAwZMjhWN/d7itzduL0iM79Pq568Ga5/1Vq/JTcIaI
yh/5AbkCrqyVcH7iWFAj4NjiwU9VqddsQjng3TDHCokqtKw0lUZ4VS1erKQxEFcweUBzgRiyqLb+
LVH4kGFvxzgU+GEDYusjzxtFeByqB671ix14uCfxlWVf+eY6yjRRm7FYVY+B/2zl8AVN6an1tf7T
3hgZ3oN9rNUxngTNCObyWuhp45FmdQC08zX8nJZ76RsO/+Rjvvkm/upLnWy9AUiaiUe0Rd4Hw7kU
wRq5LZpdRpQq/zBdXI/uVgaan1AmrrS4lTTl/0iw8G0snUbDVPI9XqcimXZZlgI5LtvSG0NAZ1J/
uvW62OXBuQRHbEDNN7EIOxHVpfgCReggSj8a+H605BhxgO+DfNyZFqB0gDNdgQJ9RSGBMXyYcy1+
TqxHnwSl+9s2une5Oc+rS7odNRum0LAjtfsiUWM9MadKNlEr72CaqWcqCHJfr9GeWTi03SbaYFEX
cDtN5g9Pu0bdHM01r8BAHoF5JtjBtGfjCZ7Yvsq0gn7ArJ5Z8dMbZGIsj7/6dd+nbdKMSl0tHACM
L2PA37jmpJjDKWpT/Oz6Y2spiHrI6KkCgOI9/rr9tgD/5vASdSLpOL4VJMClzz1x9aTpN699XllJ
WCdrpUi3sGvG3NC/rfkijAFsRFei+FWeNOlUVs1Vc9gQLpVJpfIbC3nLie3S3lBeuYP2DTDA/WjG
tQB8i+DGYjUMWpcqOlEYgn+XcJ+6E4cGyDFN8Di+zRxR4rUs9NPZw8cqkPeut9WhB9U3KDQJOKJU
LghWqPquFaPQGc51ll/sUBc5/1XtIph7nuWSwJ8Ot+/LKyly/wrc+ciFaee80E4JVZXj+sdu1M8R
KG+eHuo7lVYYM0tjmJKOwgxYeDjz8n77qx4HZSz0wbh5jyhAJsIv/hgwYizBN02ea3Z3AUkaukLh
AXp6TuKsZMaI18tgtoyFZomGarrznGUE2gUvE3zxW4s0lIPbMTm/VCD+cIMgu47IwT4g9Se9i1Lj
n2twTX47d9XwD7ZuaKbl6muUZAt8ywRhP2p1jADAWH+JOp71yMTcpfVbwtSVjjAMosqYxARhbGAg
zDW4PCrsycn0ysWU0Yg4iLAHa1WUufvNbMsRBXczJG5pOmwRRNBUDcjPZliQDIhyAmUqCwd+vUDv
Bv2cz8GaYJWVxpyxzPj0InDkdMDP7AmeD63pYKgwfPz1w7qtqtl2CUv6JF/Y+TWqtrt9vQcbL0wc
kin+nzHtTv0Pt61RJQ6aNNmNlEUTkxoEH90TniiotnQqDRKXJF222SYBv98oB584+jk7MrRstyzJ
rNtnY0ux/+Juup/2hVvEn8EE0vmNsJYbE14qAK3VeAcFtp4153oWwQAVlptc7NL/umuoDbaRqAb+
G7gdvPpdIKkAfPewR+oXO724a9ACjXbSn9kwYq8SNyf/j3mlbS9unUYTY5uOI1nc/WUPgqu4O8i8
XYcj2oE1QN2LsIqgsuSZvWQlc4rxSTfB9EhuqDA7C5ekrD78OEj4XW0cnuj8/DJIRGJx54x2FvtR
Fk+3RE8A0xDtP5sz1Qml62Me+35iDuaiIq/EtIuJ2BGGu8dlvNSncWQ1O3uhMbSKGEKRE2vNJJ6h
NMCRz0FcT5IFxoVebcuEIpZBsFRomKC9oFrCZIbkLWOSZuqgkt4xcrp8ldkUYbePJIh6wpF7yRLw
67pt8LIq4Y4RqSbeEm0dCrW3ATlwp5yVNDADx4yZvlgD9xmWB5omQYQnoUMCdhBs/VmV4gTkJsoq
a3yTKKJqhedvxe3vlN+XW2c0UuE0UYkPOrUk7UjTxX0afCSfm0K3Tk9dLT/1NW8m/rzSKhZSv6qH
qtw6MHrvgF0cMDAa1gJVUS+XoMSU0CoFI3aDz9Fd9YEGuq2l8PdsvUC3bA+B791W14y104Vo6fz8
xJTlY87JPiASB4yu/CGB2hOgE2g7w6zq4Zz0jr5YxOa9Ff5CGgR41r/Rmb1bAKnpHeJjDrzz+sEB
JPs2+VG5BInS/zvYPK9aKrm9FeqkslPjW4lh+WrVM5Gy90XSuvD9JvBqjvrC8eEx8e8dLpEynOz1
xhVBzScTalNwRGQdRj2/kHa0va7SAQNZ8Mfu9rvr4ALAlfab5ombHtMLUYOI5bK5g9bjo9fOqcSB
Dfu8HE8QOTIbFYwgZd6C6zTvxAWb5fHqRq8+cuiu257n9r30LgWWjT0HL/p3YoA/7+RYMiref+j1
ooKpdsIIYKOy5g9uygUGaOhwjFW0qVboBbRM2uzEBdA3Vm2L4/Y15KbD65k2ZRzFVzEKNxwyow8v
yz++XI92GyMOo/UsOWBDlLyGc0kZg+BaLo6wMOEc6naAo6ztqcwt/Fobsd9z4VK1w7OvXmUOd7jG
Fs26AtBp9ZzprwJkIGgKZELqvhves0rpj/xl5PL0YfnJDtRJfEerT2COcGFjMx8hEb8JyyTdi+yQ
Eg3T2fhsq5Fgss+9brkeBDbbdluPmRT39hl1mW9NV9wOHi82uC5A5/QOvfuhsbPZLodg0gvdxVlE
iLXQiRnpuM6Brd6HuWhEIGxOd6ggKaGtcoKRmQyaFhFpApROm/NeN+KlYhuyBdg8Ppm9y951TiEc
8LOssSVI9OocmuxoDp9wvPMAxFdViCupDCdcyq54vuulw0eqjbtcqPCdaWP17wYK8zXp3ZtDDyuP
YVdeoRUX3E57AG5q7mA5RyIpkr7EkViwcRSg0gTjV3k3Nc7sgYjDqlWzdyaVz1FEckPELi7LiXgf
8Hy3wecWDhx7YHbCEgOFBU3ZAOr3AVJeNDpUUrmKQknh6o9DpEv6cJWKaFFSgy0HmAoxXtxy+2/J
D2dxIEeulSw4mFUMuRT0xKysopr2bucCZAArhG6lX2oDBuMBvvR8OBd/53qECeIEVh2hvMCdhXFN
+3plgJyb7d0GMoyibW/F0EAafOv1dirSRi6+lti1cZy75MbtfwzyVOfMjSmOk3RHmM09jZvh/CeC
ARM7ZFydsxeb0X0eAKYkdBXHqNwqjP0nUsH2cDKShgsTWG7nnmzB+nSUIweErSVoBw+Rfp7KvR13
Oy86xT+AsQKOxlKR+X5gtJgYSVMy5TK9Zc8NgDE4dzC+acb9qX94tcXyzBmQLyBbPKtmx2/vurWr
0Xt7LIBbDj9K2b5p3C89vsP81pkH6yMcaHHgdKzwu6Ybym1p18wG0xpY+Iin8SWXJTqdJfWF0ist
c174uY0JC2nQN/i2snC2dOxUHJDvPrzehFIYmdi8giom8k5v7ot/oqXZ+7QyEN4aYGks4jz/sLdT
x7RxVFe7DZfwdeD3+rxLOQRn0ufM9qoZAKepl+smwBvKVe+zukSlvsb7o13x3zXDP9nroaqL/V7Z
7Il2KIE/YBK/bMfbkobZAOllywLHnYp9enunGiD+0SuutWp2yeo1ShL/btwBFa+W5MMZ1k+ZEYxa
eyrdiBqEZ4Eizfm/yKjNT8wX38Q4k4rkih0bnxbzm3mCl45y8wvE9iOjCcyzOmJ4hZPW4pZ7vH67
V59wXNOCM6H9FZepK/Eod7YJ5ptHoybn5oD+eWPQibeHuNj3rTtU0Ei63Iy9yI/oxcKC+4VFx7CI
Lqx0sS/7qsxdAb6GvxJdKgR/c7eZg5Xc9n/soeDDZjlxlkls6mM2hhbVEHmVs4qhX9HqObWaa5b+
IPQnMt0+0w5VAMgt/xLlARorzDAXiThpnnYMozdSLrhTeBdyo4b9cDV430JxWn9meNf9HpM2nVlq
nRrhqSAnVrnqHQdtZ0qHkJMj+NmY0F7/zIS/gQ0Gx4Hb1+dMquUUHAhlBAx03IcLvFLp9jTmhTSZ
IX2lcVL4Mlj55ePRHT8YnLWUH8Ft7u7uTSNmPN8D4c+3aafnLjjLG/uv4u9JSaug1dy25N0KdZYy
HvTvKlie0ZCN0IF8VgdSyPTkfjRWHQrRcTlreqlQqSDjtadzT18youCr0fovBJ8IAZLrJVRU6pNL
NRiv4N6UfJBU1oOKMhMzj7+e2/ael7KmAxJ+4yd+Vik6Fy1H/4YXkfCYGGo+zkqE72LgsQsiM+Uw
ZX2+Hi3pcZmZLpkLGZviywj1dZpGAIvq7mXg8bi+A7gyEnMR2KEZzT5siUH5HFS67JfOu08boEQ+
SZdWkQBrfir5CWJNlAg+dAjzsDYUq5jkGAizpzoFx44EnWe2deiKagB32BzxPJNWlWmaKJAAFGez
EHsVvVsJZzdk+RBwBzrpe0YgQuQ0SZxpXbhk9Kp3mSHx0zqvbs3kqusuYbN9nUwRFhDVrtPUxRnD
DBIVHzF64iCfxgpGPvklVaDr4MUwQb62w4ThzWEGJzKwOAAjjagUugSdJOhHcsB88sUg7tp5rn4U
Yt2E488CVKgukVd+Bl2r+IDxYFSrAA/j/7pqlMiTDJmlNNh/Xa7qZd7qx3pVuyiwjy6rw8Ll/VBz
j/FMRxaY1xMHhtlAQ/JhI2jT8gKVeZIYLEq0biGcHQNEY5Ud4nxaq3L0kJ97xY1iwGIUl8XG367s
CK/EAhKjo+lrroFVkelicECjRVM5FFVvH7iZE/sk7XEcFSNk8ltrxvS4pFmjHw47V4BZY/iloETi
8HeFAdwvalBV/J4vzcRUm6+Yl+7FOe/S8dPS22UPIgpCu6QRoKT9XDgRdJTHUpD/iD2VfmfHU0+N
TzuhId3FbprnOSXymLPF9xiYvC7xDD6Mr5/BUYIHnZOJblGx/w+ovh7PGb8fJyrqT3DiWhW8ZxX0
+87L3sMT0WL5KlpTcpJOjnJQJlcTcu80Kx4InKdIgs4LNFli0TCzkX1OtyXGif9CONO4jkVEDG6u
hqXqdU4F+Tog7fupfxXw8qHtcny0eEUa9RkWU5tm/1ZEHTK2UFVIkv3PP94y4kRqoJUCDVscG4b4
3l5dxEZ6FX5/i+L7+8uBXpLippb8PvYz95uZo/2W5PESO+0jrb4CsIMQJRVozpCfbWOeYuGIOEN+
F/mN2A1isWHCdTt3dC5LuI1QzqRKLnS1JWY6Mg6AhBGkouwbRzO76KWuBl4PGJRiP01WIzFK4duv
n0fLqYDfiWb7Om62cODXWsZNhnj8OTB51NM3FkRiTgkKb3WkJXjjRWvwxF87/ohiDWY9mHzH5dlo
LwLXXIOBs7Z7KnR94ikiPuw4omepxayBHJFikpCS2/UnVjP2wVXg0HDj5g7mH+XC5ziJ/nHwxMKy
IP/eQ5jTGzJqIo9TfLvQItO20JHLx8eXM7Tro3mOLR4NpeEELhLirxPhTfRHWMUkqOriTZoxfQZC
+KLr8EGGRQcQb42SZOEgg8qy8nbsEwv9N+N7IyDTzRi85pw53HJJnLm5rJdNw4FvIJmCgB5EFYdJ
dlWBXCdR2ylWs9CgajSQ8Kq6CXuXNTQi6pWCrXQV9xtaxQmy9Jjf+uAhoX9pdrQGmU8OORjE5GYR
rxKOrvOdEqHrEPjBl/zU5WbF26loQnxPKQ5WB22ooAvTuWAG6Vwiec/7WhhccTR5BklJGD64dSXA
Iu2Cn9+j7LEy6/Iu7DRpHP2os8CGl/neTpjplpvHK7vV3Sr/SAwnfrYxIaLZTI5d7FyjGE2YTCIR
cn/2PNqN8NlPCtNyi492cVxwROD+2FZb2lQt2TdaVn2ZTgqFPCzeP61mVdcZbH0R8cY/mV+5JS/t
ATLmUYO+Rd8I8Sp5TwS/xyyXOguSJniU3zbA12skHCMlDFh0JSf/Zr9hyGUleMlD3LiRpuJPwWzX
yG0BbtglX+AbOSF2PCFYfEBD0mLjDVReFJ8YRU65ualolh8gE5EBxX+FYw99c09i8ECgA6VKnbCh
sN+P4ZOqXbjGi617R9Mzq9z1JzWONHhqkfloJxCb5SqgDQkc4zL3Lc9gMM4TrDOmO/3nBsqPl4Wf
t3jGWXIAVqTHZIwkQDBWYR9iTt84WwOapAk83MzeyjclWhAnbW0XOGNyfqyjwGM1B7Pyp2S9fNJk
adWOkUzJhezp3GW9s36OhyJ6jq5DPnPpTh/46lMvIiMsob34P1Iocrx87ExWmYeaOgJNAQkLlw5E
Nm4g3k0CAUxKlnTpqgQi9M3xuIqPc0yc6RYcG0e0VYptPruCH7W2KAZMgpbxV0InMTj5fXAkbNm5
/U3sywcL4ezOmi7H5FENDTGRe7/xredbLcb8iEBe5Ohu3Pr6i+icnq9YOluDd8qjJDHaBHBoNt/6
zBA9AlM2aJaMnbgCo2WDBL7NYV4BpBxtodMo0Byd4GmD7eE/DtfGGj7sZmYaxoAb2/Ar1EnmiL7h
6lwOXmhM1amLI6lvpuyZZ5iVNvg027sXV7u6gL1OYqsFbRCVzhf6p29SVHXrZ3oVABMNbHUPNNe0
Gpasc812j7ux1v0W2DAxS3E17NFHv0REKXTZEZB8d4M/dp2nckheSw0o8PB+zbQnUPOg+vhQfA6E
6RqBSmpMWLgJ41vki31pyeREyZvhyn6BLUelZ3dBzABXCIHOWwxUiBjcSOALKg4KPLAlKb6b8JdY
3wg4r2UZDFjfffJeFC619k9d0X9win4D+uLGB1Nic1Wl05s2AyLRfyPRYO3vZTPwlmPf5rNlBzny
83HL3JTPn46kqB92OcveteBEDgANU3fGr4TGDDVabYWSTJKry3++UDiieTE7a54M528W9B1TYPKw
rL3FQea3iG71nqZdk3YSCU+0WruwNul86TnJ2U+jthA4TVKhtIGKNSGs2Cio1iKSw/UymKzpRCqC
KfJlwrBGGau9NlVpCt3I1AewOUhp3zT+La3fxRXImiiuSzLY6UPXHssP2Rb0ucOVSPAWe00RpngG
3yiG328uwH7XZGF2fv17GVEEwk9bQ1XkuVyLdLA9v/rtyKnyAgS6xJR1Bu6vPT0UqrtYlPDlYYVb
Oo6jr8wzBZJ+/tYANDNaPJfloNlSLhpxU2r4tc82+c3qMYIFUHeIfvEFDZbNK9091h+uLbbtesF/
4+31Sey73E16Y2V94IJp7AoBgJvY0X5Ea2dXmbxwdqzXcLM7pI2prnEKlDgmZH9bu/IjWbsxkf8p
7LgK33H1tUti0gHUJrFzMRL+Wq29nrH7c7JX+7MTtcquovUFWsQvaHZmGgQYmL2Voi91wQ0twLpu
7qAXQTxIQBiPTI7V9xJKj+Esxnzox5sqhIlwhAnG2jcWe5oOAsao9kz8ox0Hpo7UDanFvKue0UzJ
p2HS9niW2yPI/TLh+aguKI+VBgWlI0c2JraUFZ/ANqpkkEyQ74CF80WeEfKdCu4R1SqVTY4E7OZ7
mgcoksnmfdZiiuNg0EGjxrN7bCVaWSUtSzY8RoOiv/c1afb1I/em6zErCbqvEoCyFxmzBsWSg01b
8MfZnh8OtweUyZgnJEogzyGBy1xpuNcDTcJknwJnaTUzJWFu22rr9vIGcm1DufdJlLpbv/YjCdAU
4qGxD3ol1kCcA0prlPcB0dzGv/nPvkwtySyIdymQRZY0R/wY0rKHvQ0L6Y5cWcrLqulw2rQVLcrB
YEWl1BawgPSNORJWEQ7sWLFMElRnYSM49qT0SCzRXWzb43rwn2Sooic8ANNp47o8eKTSKANufsIO
Y1nxwwwqGR0XK664Vot2D/F3PcMp/Dq23py969bqg9hOOrmudmJde3+QwHQF4Nr4b+p8RnG+VlmF
QTjx8JTN/j+lIDNomcz0tQYQLnBRVSO7F4Fdft7aUpyLX5Pj5DC0YKluymGW+xpqCfGp7LW9sc2d
iplRufEpya9A5Jylr/H8uYkmfcp56wGrm/rf716CZMdcnZOmbeEHGkcl3rWE2KYJVsQKsFV06yUE
4SGLit6Qb1e34y6ar5eHhy7j0HpiaD84X9ehGUpoRghGaqpeib94d/1NphqmSFvRU3wfBtVSxZ/e
ERV9RCpuYMlBKBMqQi5vGbed9Eso6hcxwXckCVpQ3f7p6uNZ1rAg9nyXG+1lgt5peHjM/JNcNN2C
YAMM6CQJWIq1WkHxsEK652f4bWgKqqKRS3V7Io/gt0gb9pIHnDfs++zYTVjnKYimZoSTwyrhoh66
NqwQ7UKALSqK0YYp93ieZ2ClMO54VbSFXOYcSArBklKUE9y5uw7polkupi+oRnXewNJ3mIf+7AlI
0jO/q0ic1lvhHKj8tRVSsDlwBXtAXAbToY1TtaqHLcK8MLvJ+S9lQgibzy0Apw6iqmgjB2GatjzP
uvj/RSZ+JZriHXBFeA3vOzDY69h1YGwNK1PZRCjDtIzff8sDiynX0EIyNRh8oBiCObsPxJK49f8d
jJ1tpU2teu9s58FmK0wsajNhtLdJpcTcCKJzOUcFxONNPU34nydl9kEW7UsCcwo0V2pU/9PMka6+
IXc3KtWPAVMqwovu+cVEs3NqZ62f2zTDU+pOrhSbUnwhmF+6ghgrsavc1bylY6sb67W3eg0YHhHt
rqU7A9LTnonbSozj35zUYZtM5aPbfJfqoKcqCSCGcKCngvalJ+rGqLU/4fNWy8i8ID9mJK7giQgx
OzrCbUQ93ofnVOLrEZS57/6avnze0j6e40c8QF98p+XNbf1Xvn4ls836mn+/m4fWsgPtXbHyHI2N
whahESVggYTtSXvkgF8FysVmvQUM0/hcVyGoLRKiIurk+bKlzEr9yZLbbCYq7gneP0XwHjpZL2gg
q85xcyzoBlpsl+eidKq7BxxvOLvu31TVaohHzWYzIvifqhTmqCI2L8IPK3yf5gWFCYI9UPJwViED
upPGnzD13cofl7uG8t6oMXhisdMID5whczKyW3MtkOnm9AVEn5C9c9Qlw/iMYz2hLQ4Qn2KIR2dq
M+UHvT/jSZZZo7fzhWHf2kNAnakxcM4Qhvy76SzjWOnhP3GiuZj2r9l978zV75xITXi5OP4OPZbD
hwEjjNYGUmo7BEtKzDuBH60Z9cY4t7/76uexX+Ra+hSdD5+FjaulG1tnbuwKJW/TKBFUJULFaNjN
oCM4GuxwqSidpEWsDTPqT/POTaJXCcFRDFr/ts4EI/Huj/FEPAcHrqtPyyxMk4u4g+Ohd92Onnul
1Ql2efkvT2FT4pcwqshBAaf5DSEXxLBgElFsXxWcZDgUfIri6tAP3X/hUvcgchTBDeE0s7uVsNm/
FgPTCi51BAPYSyfqzRz3RSYybQ20jdRcIlQZ4F6Or3Uv45JHsC4HeT7Mn1TC0jhQz4JjQcYMIZxH
6/X9kMYsFq/4GRbpRFNca3outBBhMSiUzQrifC2hnbpHpLzlo04nzluywGd+qK1c4Bila5R4fJnI
YC/mxTwVJZGf2fgxg2qbA9vd80OnrUz10u4pPfDDzWOIWeMtdzTm3OcwIMC2+phhX6QMke2llEwk
Ihzy+4v8YENHEAzM4Pj0XPt6XGL3GqpQwc8rTKk2O3Z6CMOI/soLwlHaEtwyzwKPmtUza0xkYE4G
wmytHTB/OvYzDKHfIxqf89ntecpuDCDxOnawrMK/2YT0KSQTaVdBsCBzgkbSYimOX6xjmNIp69Jn
YqOEy/qKBDx9FIxyonmVhdT+eTYABNvIDI6W5Saw/HgFi/KDbxGihiijrsKZ49uedsV07b+BD5/H
D30KtsQR3twh8YcVBX2fTlNGiXFLLRcZk9W483NJD9DB+0OPMlQXnuoL4PC/eYyeDaQ6YShZC73E
f3JZD3podmV1VWs3uKrCGp5K98Id7n3M+RrkiLsOHyTf53Hfrc1xpKs2+bwIZD69tL1zgiombxTo
RtkYo9gYZPuQ78ih8JWdtq8ZJlXeIosYDrs9d+uLPubKv4F9Stjr+js/E80zNtFUCI2JdBSuYF33
G/17dza8a0IH2S6wL37woY6yVjI8L3zCiaTP1UAHX5IKrlcWalcoMJlZhRzpQsT66qYdcjW+cMnD
RCq3H8P2dV16zwOClGUdM81iBGWDu8ctfSa/gh8gqFV+qZBzHWU4kDsDULaeZucasx1sst7kbGDs
VIdn5JbYOLXbO7/xwH/+bvev356YJ+inM5RffNjyc1SXaWUhiB68Gx4caceKfft6AaVPq0UE0nBg
z4mPUPn+UUTvUfC5+9nmoqI43kNRPVXnL2fWOA1BjbrS8VDzqXg2Ysp93cm6ZzBq0aOcu4udGEuV
vw5FQ6aWMfTBfqY8p0qWQGDRg3Vm2GQ72ma7/Ji4epwj7wl/HPS+NhyHW7ndekbkdQA2Mp9GDbO4
eAbAEPnmkIT58Qk56ft/fHdJtBOWDs+8FgOwZnivHZIfYJ39pm+B+H7+9HiZXz9+IB3H6S2KmJOn
J7AVHESSPg/Un+2k3pIARspzz+zFNb1Knl8VB0Uv5YAJxdasWNcrb63t1DzM+DCq5mWDuLGR+vyu
8Sndi2lNM1ldUWcR0A7TyIn6AKnXgRgGEoredXDqeNbhQ7FCS+pSwwzhUfsHDxxOgABC6bWhu8l6
EWSWBy2hUUOCubZWV1G0nSkWP9ghbmZGgWHZIxYwBDCNUMSPrJL45R6p3bWoXzMqE4EBTwsrqzqK
6bmO9napADGK2wGoG6ZUZL12QmP0pM7E0BkRm+EjGFcOnT3AbhOzScOdW+w9DxzUOHC5gdqqFbZ8
LdqMGn30d43NY0QetrtOhBB+e282G0R/WAlndSwAyqdoWal2ladQANf++ZBqCGBVGKtK65D809Uj
aH2qs1TKSGJV1MMt0KBxwBgD1mRh/kHHmTuFWMigyqN9kb+HyundBqMiV4BSPl/BomMcisrnWhSe
cS4OI9sXP02K00Hzv/NVEVF13x5fO+2s1Bnvq6fn/PfCcGRVY63bORUJF2jpQPynesIcs4vY/cpn
p10iiB+N2kgKdLuFnalf33ZOHr8Od83iDnMoefNA/dp41szjvEBgM0M/jjeb9Brh0irnKiR799um
xMqemmFg8LJzvayyLVha+WjfFdSFo+NvRDaU0zl3/b+Gf0nMGR+Cz7GcMpEZyREojfrKyBrc6iS5
/5cmdckWCYOxiB0OItUl2LyMCBAwm4djm4USxkp2Vr6oI7z5ZQB3W0oPumVRzx0w325pI0MjV0k5
Sp9OSethBS9dEMGD6V1d4SePRGcLvqnJ500xgKeHfuSXkLmNAutY3T2Pn8+XSqxJU5uIG5RXCbWR
V96MygOaPblQGkKdOyQpctnphkLOoCAjbGaTkHk3VS7dnGERzYBHGKsW/+j+sDPZpijYLHrA1Dtv
lXZjjgOVB/XEsMFwvXD6xbPFZ4aSIIYZkO+nWVRHCFZL2v1sfpyMCln4aIQMyKJ1AfxdOaQlleWp
GLFars+gYfyzzIQp+L0ZhQQ04oNO29kMv4txJPeiHiU/cHV+i2fQe2YJkeQM7znHDi4UeJZh5BE9
U/sATpc+CL/xeUG0mpg+V9aGX5mr2dblsesvG+GXEx3m1NWFRUzfs0WsPfLGBPQd9BQ/1cfvYqZu
gyP3JLvz9HemdrYx8Ovo4m+f4jqJAYWAkVv7YGw7v2APhZ1laEY3Rjos23HNdoLhtrqaum8GIx2k
5IPwSbFUn/eBjLnv3G6tUxntuhr4Gq3xah+LRlj6d1UJ/K2tyRDd5HtU883hwicLlC9Vd/UFC9Bx
h6ifP9BksKT+vXGjcdhR6cXet/xcAXVgHbSL09PnoumIgxLEXtamrCQ+4nTIZ4n1IZGzv4RaLR6G
6sVbEWJ0+iK7i9ra6ncuE/IAliqPZjcDXOXRv4ZeNLuomWMI7p0gXrCDaf0tmYVetWSlP+Oi9Wh4
vU8cX6/SWfcTGKsOwkNWhg4XvT+VL0q7rpZuSR4j8ks+XQrxIlE16KlyKaemAOG5EVMCF+7HRcff
Rtgo/35XQuF31cD8StlDQSSihUifS4pRneHd9WWcZf96VIdceIH10T3K6GOck50LYCd5iBSqGQWw
s30AJxtN1ixbI5zcTEZb8mvB7h2KLgX1juiQ/P0l2yQBubWRPqrHqKlKS61rkKHgK+7CEyeNo6PF
+xfiLns0qza87ZANfWomz2cKXupwW45r+hO7/T67BI2D9tWTJ+SNIfw9dzC6vizUi3nscWrCNkpr
ViSgfSqxVNJqQjta8m73CT1BHybM8xxv3FayUn8GGdYqatDICchxNzKnFqiPiYz1YxQNRf15taE3
VVVRyOmsSV3C5YsdSWivausLKW7elTaw81+74ezw8nJqHYAdD0VRFmRubFJOKiwS4eRKlLINdTrC
+LenPINYgq7HM+/PqiLjjs5PVTv1mozWQe+p43RRuEROBBBsrZZSHMkWxOPRa3LR6txLcltunxYI
BfLwdzMUJyc+vxZP74ejQAiSOWsG7RgJio5yoZ3xDEfRvDKq0bqNR/Gw4VtfFfYfq4+rqybdb1Hf
rAMUrwaPCZzwSnrL00yepyZVVkizJppsshYWkgVmDOOru14M1rzgHvLvjLve+ibkZPb42BCFnZnT
foDyYoWXhXi5atX12nB3jgOrdMhzUPJH73XP4izHJI2T7XNhZl0H9G+GM+DSu1C6wodxVfeLgYzp
/9vRlfkyLZRFVDFEog+26AiqJnG67/y57BNHN0l8qRyFqSPQLPInZ9GACOdZjgymaoxzTdbfgT9J
NO/+d8nC6nG7vkKgj3gqqvpnn6kyWJovy8oqLpWnsbOyEzzI4OVYlzF/VdJXe7g0Ca1ULXeQw4OW
mQRLQhO2IOA4Iek4Cd7an/RZgwkOXVVQuB+Z575Nt8k7atul8YdBjxv7YyPNsQ4LGigL6tgMa9X6
ALhSpFmKNyrWqGUHzH5GVgfbTnb5AAkE23zv0UubsmLTAMVFZQ/ESjy/95NcrJ6QzUb1XGLs3ubI
vmZLSMBrmxBrlhqly1V9XF+tn8ykot5AaL8LwRB4ZpNib3wTAZ45ggYayh6Dd42GY8Gy1vmvnysv
au7+iJxo/1c2Z1Hl1Qpa/SUwfn5a8LF41pR8IyabYbT1CK8taXNQ5suKXJo0BvTs5WYlNPHcd/g0
sVsOd7O+QGuDxKx8gzB10DZ6E/cd2B9G2zw3Az19hvmJyRXbrUMMSlW0SXGEPIEXec/Bsz0R7IMh
UnhkFqQbk8t+I3xJoKvABvct9wX2EuAk4XLkDWRE6A3RPRgCMcRlgi402phTv+RV84PDASLYpuDx
cTZVT59wIiF/N7Xdl44N1HvWAxb071bvPZiKTfQOZUuVZbdqT4NApwQX00h7ph8xESxLYEvL3juk
6hxu39wTU0UCHCIGWQSGgzaA10jCr9r/CNK/oBVNnL1XUsG6tH69Iagv2Ur8WdtcOtt8HDMbS5ro
TlwKEIHJKbSNuYpxdn0bo1efhlevLIFHckVeuJofZKI+kf6ZAnUSvkwtdGtmD6rb09Y5kafyPjJE
TfZXTUm/tkYG0Mlj1E6zwt/FBSzaglEEqkn/kpNUboqgSG0LJLQ8NM9y18UEMjYsK46QcRUo0gKH
JSWch8q6tmnyb4DGOZzN3yx8uBa3rSLMVaWJRu1mdGabTa9LT7MwQKrjCflKXexChcQvnLGz7Ns/
keNkZ9vCcJA1gl9ANhvV9PGqd5dOTrGtjQ07D6EoWRO81IAktaoyHG434I2HJEAXuSS9AtFIDVUc
TEh5Zk/mqSxqEQEAMnVIIGLhyTQmblJpQo++uUxbofjKIzMfLk/QZ7ie/CLLAB08N6tPlEAqMkKd
L9bLLLzF758v+EbTzkfDmNnPlb6QS7ciSFAi4vAoo7BucJh9rHqZLS9xccSDR/lY9cOIyWusOuBb
acE6Fc2yQgGGHykDMrToWCctv166SRDBrJ4oDLfEI/RF2/deAD9xyLLtfwInyagOOyebWFtkI5w3
0ZRyenhy2rHIL8pooYgffNnW4NdZ+FHLWjzBqagyJQAQtox5gdmUUgBkhRfDxKxTMe+zEIyCXrt1
N5bQyWKS5q0fpGAmsf3GvNTcXApYJJ/8Iz4iNkxqIyMBV1ScNrRoXlenJyZJXICe2W+h5yrhhEyC
Dr7d0ZNyyRKi07ICiVBgJxK3f2Q4vYHti4dYCEw2M4uF7e4G7yFsrzN7JqY3d+iyks2igePYlZn2
JP9DLfQtis6Ow8TeEz9zSi3RHWG9PhBBKNtos4SsV35jaEJpYECAGqTBNfUsjTmC8Ir3nJ2IrQBM
9AI5xvXTXQMo8DSk73a37jdz4ywY+aBMd9j/zrNsIr0HzmWCORFX2jSBmM7+D4TxHDc9xqITf6ug
LZD8hoRsFVo9mi1VBTREW/wTU9zd0ft4hrWDuM3R66MOY7jOYNPE/dqbq41OjV3Rd8Yfm4VVu2uE
JRo1IdCN6uoWFuGBCMYQb4K6ZuQmrBQ1qJM3VH/3QghBj16foa46JmpDaAC2OGAjLtKtL9zpipOl
O2IbuzQOKtIEYTI5i/rMHTf9GV0CKMxheLUPVANy+5v7455ffT3NgYyGscDaKD8AWX7PHAhcqYtX
zaBLUOEn3sZR9pAAx0yckwEEGVctlfTHu7HbUrRSUdmua/6BwS0qwTS6ZKqpQ1H/vsCfbL+MiRdw
+r/QLXR0s60Pj2aXCkDsptIbBVcEo4MPFKCvjy7HelRffY7iZV5+pe4dUDr/L3Wh7tUYqoM5IbnJ
rMWte6+BoSmKTthCmvF9OtM8vg710sYLQpV/sSBp6yjrkztZoMhUmnaZnItYoJmzVyEVt45W7LGq
KXWtm4RaOmO+ESx+k8UngP7edFKch2IYeNeWhO3dW3UKO6mP9QjBys57jzand3ATeAeqWngxxHBe
3MIwn5xloYoXFjq2qG7LSHBp37C8YM/wG4E8ADEgsS1it2mR5e94sMIp+RTCbY5mEsb+4+1A+O7G
WWVXouz1Gj0FJgzKmsKBEZuDSI5s5iFIjI0WziaflX11jW9ZPD4nEixWIG+UQZ9bCF6E1H07gpyy
8quEcmtpFh2/agNT4BJSzKR8VVCx7O83sXCi+JO3mPBByTKWZ1SAMOyrR6Pzwk3iI+VwC+iFcA0t
93jHDKPgtMCVAnQ22neVaiplBNUXDZZMolXzOxCy7oskYD7X2r61x+VC0zG8QLgl8ON1k4eW3B0r
rvxmCJJ4p4+UKeQhvcq+o5kvzR9tAif4rc0H8U8RTO6uTmur5asF7oFIcdL+W6VyH3acujHZv3o/
0BFnU4E9YWdwnRmE5lhf7XI2XSuqMEkDWrShl4QDZGmjT+yVqDMLg9Jp5pm5KjsOLSbc4yWMBNIQ
1+j2TxeeyORrq6zX7EVbfitODoThNHJeyH9LdMNBGqM0eEafm56M08A2S5KUORauP8x2l90tGup8
Fs5lBcuu5gIb2NRdL0CckkjqLaZjrVEhdis5TIqKgIV6uqYtD/a6yue69Bc8CubkB+xn5WdNfdtx
l++dDqyxkywlymUu0vYuOfhLlkpC8syekS6pBdme3Wi83oPSejI0HetUFS/qKCb46KDd2d6s394X
p1ZTQt3ls2cBVE8qbKDQwfWdWp8cfoLBkCC0o07uL7Ci/0OyOv2OgDNVSoIwYJ6K4rN28Niwl8BL
mcnh0ceI93nwZ5Qtlx5FJjf9wyvYk8QOr89qGEK29dXw9cxTbWlD20e/zzhobNGpBd2/79MbHLzw
AVvrUsEPiuSqdhORydJlkEbPBL0boEig2dN6mtSyhCKrPt947P4CyFzmrwOlabz9OYPTLFO1ggpR
mqOaTmt81/IraKTmLiT//nVbm6Ck1L/p9sz8JqmTn80oMOV38UqdMX1j0cGisGNpzK9LhcJ8EaQr
UmgZ20j3XNXBkVukomKEs+q2L815fw9XLsQOrBcDWpgl2lkBo5EJYc1X4W98Jta8rRWMJVLSmdQW
W8nJ72fnoLS1NPhL6GvISvoTFi5UBZUZd4vl+4gJ7qWOfH7IAGUV15+UFUkdkrWm0oO5yycgqjbO
vPKrK14yPzjB9STwHW7W5HCxvHqIs/BMYYcNg+bX8V/iSyffqEFI1jPI9wLVTdjD/RIK0XRvYBRl
0U8lUjNtOW6v0XykQ+rOYwtzl6gEYToP9xvFQ86YUR1yAlPh8EMwR6GXXG8g8kxFqzCyZp44pze/
4pnfmnBxi603S0i2IZ2hsTAcTFoVjYq2kMo+5VA+P76Sa+Rnh7Tz2MVX7nk8J5hr6lmxkBS1P9AE
twO5OkNzJNWtXl10FlszpNrRhsW8IOOsRHmYMGKRicF0G3nzI/Ih3IkstfrK8G0bJus2WKAe+NR4
5bh3aKbMGCHQnoLiTvhLyrt0vxTySVWujvneSaPIeLRmlPW8mEUT/Mv2dTeyr2UABaRTUhr/YrqQ
yjK6v5wtXYaN68On462iZU+Y7E7nnpmrRRLP72yCWChOGV4T0mcMrsmBxdHu75fb9v8FoPH9qTCZ
DH5sJz1SriwDBrOpO6lnMZWHiGAmweGN2Hqa064Hi/H+QG7iZHhWTd1tX4DcG+In14nME45fl+TE
AL0vhmxiZPHRTSlbQkPJ/uSEyWMEslBvg0Rr42M85cL0JAVv3ggvEupngSmcY9jU8mLteUhRTH/l
y81mLQmUAemCrNlkOIf3bYlWPo8TPzp/bsDlAsVps7WhHWhvfFZUq0PUrgv0dw054OsMGgVYmF04
dMPLTyQYoQbtNeWPcJ5SN/TlhUKpIAg8w+Bw8/WKXECndTiOoZmEg29+ZjFrZJJKyYD1HOJSVNsX
HjOPFlViXMT6DFzl+CcJ/e3XPiLK7RMAKifzTnBw1ZC5vtx6L+e2KNZV6eAKYki4S1V9xGgD5szg
4NGGpHei2gzajKPFzkrR0KYjhCA4nrsfiiyhsPP9JqucjqHSHRDKo91DvMRGN+6icKZXb3pwQM/l
lfOsO/XLHXlnwnYwwb55Uyf5obnh0lQ7AycxXc0He36Q5ZzcRpQTQHp6Dtvn9l2cXocm0coa0/O9
pFqTt7OidEb8dXTk5xUCyyRdcE6IRTq44439v0wCjg+mpjgbyC6UaM2ip5zhnyMgEjeDxVkDQx39
K1CdPqLmc/IzqS+Y9hC3qVGduGw2DZxLJLt9LWVu8/UR9Oe/NKzoN+PlcMTgITSwapRdWO3cAfJp
FIsk34IGyJlg6Y2YDxWIr/42zT8dVjCbVuFXNRzTlkqlZRkwCK/xf+QboDW1DN9rcJwcaPD5kCCn
zGEQpCEJIo4lsaIoNAezyHJ6ItlXnOONxDT0sJGpgLL+BulsCI+aPH+UdyosqH7xjqGuWPene/p0
OWjm/GVELtm1MdkYE3HogXmvF/uGNFlRWIu8CCJO3jKwlM/EpwuDGoY1d1hJvMMICkdzkJK/8/lk
BoWhPfEKv3X75VZmaa6LfFzQXpWWKboEUCuNNsqKpN1lWww30CCqYpJS5SlJIUkZcyR1aasL1AVr
MVrvmQtOadb36l84TFooBLmsT5nCAyVH74AVGmwXnmA10BSellCyGYb/+p7kV2PvSbb+EnH4hXqG
w+NDFeOmUb1BCnKhyL3EQzIFnVwGKvOj9lwiDlKQciV+xzdXC0gUDaQasP/H5W0vxDeeA/ahac2+
o5qlX5X2kVCc9pIEdzKs73FzGYkc6u8yF98TCIDKXGb0YRtoo2eDb/rhhtkbWwtsan+n2/n/cG4Z
CSrRaQJ8X8wxJfRB9jfnpvvZI4vPGR+tWWRsTpBEQHKZpOlLKVjRpv7fhwSEydlx4Pf26lby/8Xx
+AyYXHkaano+bHc5AURV86pG2r3GWooEejfrMwcuUyHIPwy//se26u0AvVq0VzGnfQ5WKQipbpmk
WtlL9b8+QtKWAsMmKuefCkXdf8i80CUaThlJtCLM9eY+KSVZGawaRhLhXbR+gAtS1O2SOBnWhD4s
AvvNy/hMRxuDCYk85etJforUOlkTlftQBwx9QNimAuERxlXTHkL8d6zR4Ps2xTAKyC20HIm+4vJM
bpfqYxfNwKvisRxxZTxcBn9fJF9U8r/a80dfhXixCVmj4iHpu4P+acfA4vN5bGu35aZtciU0rHnN
3WgsdQPS6VxqoV6VucQWM/VKOq6iZCAqoNue4snIWp39B7yafmRIgN4Zr/EH91L4y1R6nx+BBkj8
iBhdc/2AOiXWxb9pnn00nWDmyjxBs0PFN4Ls7UEsLc7MnXsgW2R2Zm+2RDgjLVlEY5YLykMAr7JO
tDTx2c8XvtiCuRxyHKAxrhaJ0g0rK7NTyXUet6Fl8cZJVn6N3TU2STAdwHiNKynxr6fF1/JCybgp
UtzILSGnw2gJB/YuMP7maq/Oq0pvyQKTKv+q3g9X3wYAgplR/bXkS5VsN2vfAiEAT+lACXX1/9A3
I30ONeQLrTjEAm+GN0pX9YTuajBA1OR0EhEgT/Sd3TPyGNnmLTwaIDHbtYBxDPalkNxBvKlfp3Nz
ST8BhnpOc1APypbuV6oHeLqF89tbv+jjtDMBDyAY0BcUEdomTMsDBcnJmpo6L5z9qOVCSIiEZ5bo
loohCT2Q4p7ecopShxImDDV51T6WUuWhK/o5IThB7nsM6DpXa7irv9TkefmMCFz7w0M5W392XpNz
99TqMdg7G9YRzegS4B2c22OXXOvA9c6Rmjt0Oa9Z+yS6hCUNM6espkP/0FCvqCaDLXwVmf9z/nZo
Rl/ieCjLKLRV5F0grKJgLxboieSsfz0JVVCC5N4d3pkfgTZAh2g4XWmueSWAY+isoB9mxfQqoNoz
YEuAnL2/OLPfGeLxmAWyxO3yN/Ou/Bwngltyh2HVFyElYt/RFrXX6ndChErNvHIP6TwsU4fo+X9a
0Dp3NLRAMsNRGkKXFj4gykdU/CW8XIvbtnX9M4MLTkvVRRrkBR5dAibsHSqZ3F9geLG7w0Ae+ePo
zTgH5aIqMrjaREEThLkqFcwxueVRHxgU7LupAOjsVlAt/YtAioO/1UsmaSeP/GY1hiiD+/rOx8i9
1JEz7nKd/xOv2Vc9XjKidIzZA7KolKAygZsOT2J5ciFbeXCFukLycDUr6aVMSz/Mr0WFgitN8Rjr
6h3w3syeYhtnG7WzL/URMoVdlatbqL7st10L3jVSe81gOnMmdUieBPkdUbS3/qxyGDjf9HJGnl2C
8JxW39hQC42Wxg+cH0FDqXZ/8K1BblQDWej99Wj5GAzFEKqEbGz79umfiGjQQik7XnRS+mSgCcNW
6JIDMIcbvVup+2lycTGBM3CTazmFhur6pSn6sTalO49bhD+zx+nC2N934qVTdoZb27TVDhzroW0Y
ag9XKOGyr7eKuK3NoJDVVL7zaaBGCQJwrLdnwtataPNvCI1fhr3XoP95Tf0Ufqg+8NsS9lBO9RSv
s271L0uaLqZi+e2e21D+yYtFP1UqkcPNjTEiDoxJw2dLDP8DrBjSgHeQ+H510rD/nnbyXgDDOeMW
UwCzXkYIu6OeR42TwB/Vs7UcfiCqsyZUkdgKDj8JTNM7WkpGOoNNFvtrDaoXVvF6RyHUHo92mGHp
w+yRJ5q6axMLgM+5BugfNI5IDqeJU4Z4fSoDPg86pEdDUN55vG9FEvdNy/E10mYu3UhPD08VvDYw
t+xaILBqsT2l8by28PR6RA1V+k69fO0u/GuouBOvQHZ6nvNnMwFSbc1ChHPAOfxWciLq0iA4/x5T
HEV6ve02CHTjUvcMGX2Jz1E4WiW+ntc0h2XOOEgkilpoU8UpDtS6sY3uUUjLj9hTpCPxDPCdOMAB
YoHjQK+HwR2rdiUncGUtxIGgiatCyncv5CEoaxN/+/zeIkxdhdVHzkP2TXrhWg2VlJIxB8ZeIRLr
KHZM6lh3mN41FmRivUMxYoULUSyPrF2DFp3/Yy86ZuB2yNnB8xbaEnp+4PuLcl4b66zFlb+GM/tI
NfxT6pVsa6LUvd52urjnaEcFI9Rh/rCaInlkj712SIKV7JsEIxDr3f5NwSlmEKqSlKd3Nz2LtKgR
oouWn11tw76XFGhlnWg+9kA9IAidVdHwoTGO8TV/+9eTDlqHJt50zndG11eIBgcHylW84Wi4PYYL
q+qMaAuCODpBdj/ycMWDqduAw0qy2W5L9VOfeVNdwsg9+d37YGLm0wdjPVAPPJhcBcYzZqdQ0ZlK
EQkgvq2ohVRJpCQQi5tNgmvu6yvOZZ4P6pe4fzhXlo1O0GrC9PWuOVkILMsEpkiOPlX7qIr8nWhq
zxbNaDN4pZ7Xrwy+EXAQVfniPOGyNWUQEZUWLqsC0HS1jq0jAzxdcWAWZV7ptO20Bga0rpMF71RH
ZJ0NrSBsmxezbkyUSXWSUsHdwwEpW2wqeoNbF3cF3K5DQFuK1U2j7sID8iDRoAiiesfvEOyUXZOn
Btc4hy6/KQowFBscryNO61AFsJXV+bXx8qG55Y4C/JnI/7np1Tf5VqkUWL/KATXwOka9pHt2gjC+
zulOAx6iw8R8BqkzZ3VMfDQ3fJT58w/mB5WJ5rSiq3jtubt0eMnEIdmaVUhOuWkNBZBcKLHg0gj6
/21A0MZFQfM7qZlvmXIMsnDaDbC69L4fiZ7xOvp/NjY5owTMyn/5QfPdTXcgRKi58quEurPfPVoR
G9hSzUgttPCopAgyyN5nuGgivR/aKPXTnCl8VMsbK59WwVYCDfsLqJhonlOePydAYHsVoHW9X414
uX8D7tBjYp6tkehsPt4EstoWCHJSUMLMnIcJCC5/dQQIe857/rQTFaiykbpdfh53BkRWvQNjliQa
6PDC91KJOQRMThCeGAtFc1hG9SalEHFF+jf7TWC5lYEXqcOfHLTd7UDLOQLGQ8KbKSNy0CNiQ4Sn
yrHMZYxgyuhQQFLBKnDqoTyV/WMR2BYjB8P18AtMRtuTYdtsyR2DPdgl1umx6S1ZVMFhkBlTva7B
85g5yKGBOaVDG5nAxuTAOpB+Vg3uFgLeEszAvBa+vgefGM/zLOwmbg8Y2+zh9BRdhKlBLklCoXy/
70LLnlua3IXE+2dKsKNZbVxYFnmbhP7qwcGrxTv4O/SsUWaL6RX7GKg4CScgdtgrz6hz6KdXIKEq
DReRr0X/u1AyB68k8n1k7pHEYVE5e6JBNP7LFVpET77QNZp04oTogN2OpCG3uYOMF6IszbNqFUwV
TVOIQsAyL8l966rZCp1i7V/S6cJyucOFc8G9z/YpMs31CqeDces6g9OSJZXGYE5vkVcgB3CMKmIb
M2m3xncuAlRo23zVdG5hXCaWideiRqvepb52R85SVeB3P7uxbvk3ReJtXLaqah8Dl50mz0R2F3sM
XF2E990+sD46THxkv8M6UwJ4LcBPk/TUMZVUcjTs9kUc6GYF2HuaxuFHQTt1hJ2rKz0HKRlKrCg4
ljHyHew+JVr4Uviby+1yvwwXIStP39Q+bFjbfiVa4Qr1SG173C84WOl126JfgwYxh/vviT968/aq
yV0z6kf5abzt6bZo+Y8JTCVWbuL5WbLHPpc+5EouUTH3emDvhbwhNE9zCscZndSG7X/xcUbJYbmQ
e+lVxf7MDRT2Sdhdb2CQ3nfQmKg7Xz/g2KntmmZ/dwVUi7nnQcwnvrOoKZViYmRtUdhXKw1mPAYn
q2giw+rLSyTMhVSOkBxIGEfjibxMODjT5haMtGM9qTz/8DVI+pNweyJpr61FjdQdl4psT7JSRHE8
8JWZa+ULcR/N8yHxdHmOxqSPiL48QOS/+0XXf/ibAuymd7t1mWHvtuz9u3VrwT622RFtgfj7z5PN
4zZF4tkwDjbboo5PjXZJ38KW5+GoB5Cvos1T3EQQr0VAftb3+wN5JS8/6iCEwmeIJcE04d1KD0KN
0/kvH/VRHPYZ9zpTc5rmQtcgSqwZ3+BY3pj4lm8BaZfMPbmHVX+r72RKjqAd1V8KX6E5bU+dCnN8
z1CV6csGVCFTYbIwaBZHK6yrkijeBXkJvJtJdPw6v9XFffQZ1KZoinCRdP8uKWMzs0zYe3pRsfQJ
y6Lb5VCk56zZuHEluKmsWE52cG7wc1x7oMy0UcAph50Ejt4JpM2FeN6MM21eNtiAc6etBNAhdSC0
maKuGYUIyJ42dhtqPKRuOe8oeaxLV5V8DjcVdarCrarSAB7VhJkugWf9ZsL/EO4RMBxYk0WnMEfI
BcW+/tsMEfsGFWotefpcV+HV7hNxxB3u6DknFDNMbk9v3yY9qsq0GJHuipDV+k/4hBnwGIaF+VAi
709NffqndTEsJerDVA87a2Ad4b7zziYpCBi3UxgHc2YUsx+PL06097EweU5lnG/c+SCOCOx7trLf
vl5vH443eEHJbgncgBII1dK+6W6XLwYQ/tQCYYuRdf5sQnIWCt69yT7jg5vxFRcRP5vLw/r+Lis7
UPN6QOhZVChkPQdJjr4AQ6OhYiVd0z+RRwRI0YEniQ5gU66fb1nBL0vEBvZC+t7zlphiY5qn1aOx
VjZ/iNz8zq8GoFzXg99DDCasD+5AAlK90EFV3E6xqbhGek/ArlmU24fNr+3d6BCfs5QplsJPR2m8
h2zQCkvpJzUzIEoU7Mktt0YSobXoRrZQRYmGaD4kgiomfVRLaVHFd+3bcp2E+a1236xWIeegMXfA
pCuC2Nvgi3ZYPig+ak0jBG9VBCFjfwJeYXl1rQCM0SuI6QwdrHrwJWBfTeBwufaHuBy36uTDXddS
OfvmoGTc5I/BPh1h9fXPAvX+NQKV/xaoK5CfY9Lw/1LZ4P9aQtDkfp1r7tlEIEcYVfDLWzgy0/0A
okqyJxZ8Pd8Wv7OgoPZkLOgKrYFZpJlnjRHd+TUOEjFL/cqj06eFnJJ3bXC1KqGAUfNI1J63VVV4
qD9JL6o/bnrXJV71cfAuMEkfL5g/VZoufpP23dpj1hMO2ctmHcW9boOCKehBSQMMl40MQM8W5DQU
+9Z66PRz76xqYMGBvX72cMPDYobXWyuJz/uT3epL5tadVf/TcpnUucYrnmbe8k3B9ZIOPz8rWuvU
K9k9VHr1kJ9n8VAcufcQvdvhEAgXlHAbbL+ZgPwtkHB7nTsxPc7PmqLeYX6Z1+AcctgOL4MPMWz9
S9rR6sWqkCQdh0NQbyDnMSyyqygbYSeJjgK5fO/HKK7RUGiZ806MaUgd79Yo8DkONdtii+mZEg3+
X56QZOCUTofwL07h+vj1HvVNayCaGLTJV0N7l+rQUMLFUXA8odKxgdyowajSHujcp4wahzXkBVMR
nlmzXtjXizLwBg2D80fRuLvqGE8XaqCCXd9TxFKKDh4ObLEYWG1mwGjLZc+PcrAKeJxSZGtQ10Hi
FoAZHN7ZgecrR2Nw120nk33CDfsrVU5iHKeusm6KBxt09lYgwOLSTboKs3KJDLoluy2FPX2xJxUc
dPO1qqta/JF7yCCXsnEVbniIZ2AcODaZoqsZuRPZxiKYvgmqlo0c9wZAdl2Q8WzlnHVbpItu9+Ui
i1Rxgx70QfTGGYPo3VBfBVw19Wiy2FlY7cQaFX487RMGULvE1Rb+yInLKWuY3cAoL2r6lG6PCYVG
WPnb1QirufV/f2a9lFQUICGP3+3ZvC4GGvJrwqdXt4AMXMXWScEByagKGUF4dFQSMU+mKtKgaZZW
r47JGbG97v96NHs/I7LNM51rZG9F5093Kz9OEa75b7jRbPTBFHm3PRJXYOwlbNW3ihzQ/HmeuXS3
59nZJL4y0PDK8nrAL9j6Yey89bmI6bxUvCG4XpI0ZAO/qVGFJCSLr2hKtV5exbq79T5x1l6OD5oR
acGVS3b5U11PfPrxYyszqvKJVwgSdufmAULDKe8wGiqOE3c24IRQipQ6wWQVJWIIWFDb2v9RRnTV
8O32EkrL+VEcBM6gMJyPPBEizTUJhpFnXWb3aySuOgSRnIQGA6uB6x6D3DpHkdzCYx/x1xgxjOg+
uaq4EN7d/zXGiBowK1Tqv+XpO/9ychZF1lUdPYl1A9DS/WJnwNV0dGY57l6ulItJ1F5kRn2/7J5z
80Wh0aCX0GjdnK8QXJoWHTMvBaAnwkvlDuHdmLzE5lTiRY+YyGdomm4JgwpHn8jtv8AbuBBYLpzm
DDbFnVWjNkudWBIrSTl2U8W7rSNvazOO1+abOcBBltSNc6OI+uNwOxfwH/a9UMJNK0nm3+FAs6uD
pix51WmGa2NirUkYKfaS6ZC7tUK6LiNaN+zyUUdwLq/p1TaOMBGRHXldgyWT1kba9//K8LjC5BZW
8I37sdhTvRKQDUb1l3+NiBlJgFPBxiEfHgWni7aVewGOSb7nby2/6KeppTGExavJDBUdUGMqb5Em
m7xJbf6DE7hatt1j+/wHiRNn1LSuTHxGFavpWX9mb+GnB7kxY6I+35k9WNn65Ut5Q7727RfWeMOg
7+oiMaS3QCeM9aSchlPDKyZuNCCCd8ExilwuT5k2UYNUepsE3UqSANUwiDdci3/M8ilwkmY6NhS4
KX+mJkQr5WoXbS1/FhZrqenjlV56fYZQ7jqpEQCquiSO1rx8+Bacfcu+Vom4hqIYE4N6gwwB1tAa
lQhfaCa3iQsBLGn45rgSDCfa3kPGnEYD5PrLCAjuDE4jFJZbrbvAxH5XKM17grKjwcAMYGfCyhIU
L+CZI15ey3gp8VA4e8T6seMoALMvKqD+XNcaz5+iftpCmN3bd4Uu3TDrrxI6dblRhDDKWXG8OMgP
4Rw37ycTFFJyuw3pnYmefj4e+TYMHiTimAwVAh99ibLU/xQxmnGseZUTeVWV6KDGuRrVkJpmYD+m
jGlCsm1tzvX9GPyah5QT4GoB1r6XJbUdYtBVHuuYV0g27P4ETxhhAfjK7apQo9EiovuQLov/JHWL
8t7VwiMMU/eMbH1FigQHrkTPdjzXrdjh3jShoOPmC9nmFnAeB+BGfU35juXooh45fD0z8Ac9wiFB
qJIkpk+XXwqDQ7ABykjM8A3YYL1uVuUXn/VBRE04fW4dCYsvlFWK7Ayjpxf/XwKKE5KUHA9vudDH
XvCnpx0csmd+7wbfhG/HblOg5KBfN0APDMAsJJ+kAZ3qpeQqLBs5d16LJPXhly1d8Bp5K5GJgBiv
An1F3WjkoVlokN5NmZ8TiSB/3DJJO3zyuHl2Ax1aQfiXeMS9qswYwbzubKh1uNPjAR/+o/NHHxyP
C9Q5j+qmk+Mou/rDabOY5kqzLRgcO4Z+W15URSiCA266UX0OR8QoafDBNu1PzQhH14pk+7P2kRmb
TWxHdqnrhXY6XnkmGZjiRp4dJqymSig09flqVqmBnDdw+aiVYr+tD+txjEP1VF8AdVaKB+l1Urkb
hzKuAzNy4a7HKda2v8vUXn3/Bo8ofgXwJZxpSNuf83junWDR9OL+7+hcmMLZKO9ZlKTh5i7DfVSN
EAXdCGq4UMxxOQVkmkMJ3CktFRNRhsLa0rU54Hv3Ev5bqloMMh7lPWc1zCSJXlO1lTTzGE1bwD6I
AFwJW6SnOiVBaidFCJxKkm5K5ChFmTWl2+KqvePxTWZ8JYjAlHLO5ucLHiyfmpL9wcxqRFoWuq+2
U1NjEaiSje2dqE6Y2HgN/QVM3VXTDhh3p8qMreSTXWO3/g4b6LszPBDKlnThzsQz8/pEtElwGrPB
3yK7wCVow05fWmvl8iQzT54JHTltjqJ8fpiXEpVtpzN7sE7GRmGAYOFaXDVX+yxnB+Q1fKDnZrqU
3okpy8GypXjfu48YwO664lGALQrW2QmDV5x7y//hW2FWx4+nTxeVkraY3+RpIkzpYBuCZnQjZnrC
knQSdR4O2tDe9ta1keyOwpB2lE6JN9LWh2NoPlsTt5uPan1LUC0EkYZW/qw/5vCMFIThxkXixgs+
WFSLbAbucAi+KWk5RWv3cUpQeKpRZoR4qn3zmEndJKv4dQet/ssQfGfOn4zlKpk2Oo5xh/OSFIY2
1kR5Oc/66/paQXPsfZnbmN5nM2BSHqUFJgQBW+m7KNQtcacummJShLm6K3fPZ66uDnXNyQZa4EEU
4ZfwU7ECTM7eNOgDVZyLTupy5uZGcvLg/SQHEpi2XZcAy64Vh5TT5njloleoiWsYT+3bVxiQ66Sn
hHKzMtUcU/fqXKS6nEdaS0gOgSnFdPydl0qeZjOVU9YGoy7mra3AiEvQVnp7qul8p2mJvMK6/C8u
9y65mOXbu6qZ7Jkalxsp40lqeAchEzIq2rH9+guwAUO7+dhbMYmTQfLidPWrX77GIaHjy7gmJIms
ZG23/d6/z8eDWOho+Nyn1ZsRa4OfkGDUKtG/qJ5Q6curb5xPJQyoxFzwep0upjZkwv/gwV+nhnej
guhBpv3o3oLYBmQxeVAjy/wPxlttNw81McX03vfIP2zdkMVLyhkOVAH7R552S+suIcbPC38Udsxb
0lhXReHjXzTw05SKIOViaWGEbIBaRWgaxMX8Q8o8TK9wvicgqwtm/a+b7lPU1g6ZWvkZlGZQzs+B
kHs4ULXcjdZNbwXYAwqsvPhC6OBTmCr8cfRVWID1k/u6nxDSuk4vXmwXdvr6CgIyP0znuEw9VgSc
cOYxp0kRPeg7m77J+FJ2O3t6doK+tklbUDypUiFu5ocZwSyHeveW0BvSeQrnIfpDq0kN3nLtlAUc
eHe3hUQWL0EJD7tiCeqbvEvlTPTWJ7VG8iVimMT+k/vOgUkm9RwYyCKR23V3hZn/+uCW/1ExSh6H
+brDmAqBFsEt/H8HmP+0UUS2gBLpE7RD596vLAvnh2RpgRH/p/7NCceMhDcYY4F4K7VWlyNOFYvG
3Li2/5ZlEtQmFdSh6ztYCHCaxZzcR++8P47DYOlb2uhEUkDdqQbwNC5o1ci7kTZLGZ99qTW6l0Y4
E2UjdeRbpJvXu8FcfhW1BJ5gtglGaNj+rHgj9s/gUz1/rdaR+MkezPuNWTQta8SiCYlA2JXStutt
zijXWppRMdnrAkjAE4aSbci3fIcVnIbapy/U7OOLH0dDo05Hu5Iz2X3hvKXCDMFzFgZ4oZXCVhkB
DxvBn4XRrilX2M/AbJnhkFhEUitm5S8FtP/0E/+yAXPljB10CaXRQRphrEoRAjWowMsqV6bLJr/D
pxnmyX5yyOvnNgJk4HpqiYdF25Vq2Yox9Ib4rbtAtKVk7z2yQRg2IiQfJJTX8Gf8h7whYAGwhRnf
rTEPpMCu6EsazH8w7TC8yI4QkWf8Hx9EOl4jkQ62quudSK7H4dB6NvJeCA98xvJjfAIUiGekNkG+
BcHjDCLhvAlcyflE98rDudCHXvplGVd2eQTYt+q2oKRr1h5JDVMm7OILMrEhb7oj9Ol9owLu0nOK
aH3e4QSyQr/ihGF3eeyLp7BqDC/RKkvP5TWkQg+9Ib1kQ/yNq5GtE5Jga0zrHAKmVNhgnEseWJDv
criAtuIlrJxS57qq464j4AlY3ZfklANnX/YZ4tuWZFpQ4UV194CiJg48Pg+Ls5iptPQ/HzLKDj5+
jGba32AccjyKJzMINU3lPqKrO6HTt4RB5f3+HgO7iTbKgDdlvbdSwqdtKmeXjexp90bI2mOJdU6E
T4+4Nd7k+a1tQZYs9XrftkueprON5qqMYZo/EFIepDVzRW8pf39N6VDJxwsj8g5roydjmuoLbKL1
qxitNwpL7BUQd2q7Xkq+eRBfSo23phWetbenXrFcy1rkIciKYsDF5bEov92QT9SytTfH9UT4ZqDo
7hYZ7ji3CBKsQhBxLxQvILfHh+ZL1mWWtO08bDeeyJ3PY9f2z7Cs0eu5K9wbVBMiKxDxMgUA5ZUq
p1DnF2zOsFDWZ/9AcRptJC1zwNpinS4lG6LcVhR3oHJ3lKGLmpyeOM/IUfGqRw4KCgbR3oGd3Itd
zrQdFbTg1yt3UZmprYGhB2OVqM+EnkE08dKdkUSnEm5fblxZJtuVawHsi1HDzJommWDcFYMxtgc0
urteuAqjARJWgL25hq8yO7tXyoAjidDcgfbT5qfM0f4hT10Ra5OFQpDD0V/9Mt9M/qR7egy26jLt
9VhUHhz84dUd9Y74eLeGsPc/egBV6deIujWZdA4jVtjgEPOSHSbWh6Gui3xC1BR3VhiajBpRu1I6
Aion+3ITE3ubm3T2oIpKGbFAe6W6gQ0QHepQBvqm4hP4qN7pHzlEKEbOdNxgwblWJtr3RGwBr0rX
PoWYKaHJz4H0b9Owzy8lbXRXxYgys65syYYsm25bBN7OMq8oGZL/OSCbWjp8IcMfXC/fY4+kI2Qq
M4rngqfhvX1DsBmu7CYduuGVlhOwg3cFVGSU9r4sEgW4AgfEAh80gDCxgk6e5tNGJgwqmdC0qvQn
02YDpZU6Bw1zSYmkJyX8l1oNZoj5Abaeng/zb3fx55Ae9WEJ/z2uDQElAPEYazu2TyG0BY0rkgam
zt0pq13jlq6fYpi1xWbwuySy0P9Wrszu2slFF5mmVHw8NLguwOfWplCw4/wpErMmMEgmWGPTqeWU
xYWUu4awgQQIyC1yVmjK59cR5qif5D6KYJqLtXI/jUbgP5+xZGqsgILD31oF7vtRDJ4lSJNFbzZZ
qt3288kuRHm2NyaVvhPu6iMlKRLpekIWajh8FJYdLrrCHSxTgigTijggqEzwzL8+fTBEk34yTiL+
lV8vmsnRG4mraacSHG9UcgI9mvgTTXAy11khGZVIUTPhj2MKJ8RzWS0+6MzP0sg5MjBB6/debpcQ
98E5ZUurU1Rh4TIz5nWvLYtB0nQ5a7oTCGyGfBc02FUr+zY1KOuaEEPYZSY3D0QVtbEm45MrgJ4f
+yeWC3IHSz5QVrUTXPB3TBRRx7TouEuAncONxHjp5JWnsngIR4OcGXlnXukPe8kEjQDVcgwo+6oz
V1tG/t8SV2Q2CKUziPvK/D5nt9olJWWPyOTjucoGs/wDQAAC5YGerqIn49+hSaz81hhyOtLq213V
IEa/xFptz12z8mJGweRA0aJgDPGIHyovGcea7XBAa8Ou4X4FcmlCnmPoDuNQ+vTOxK8mtumNvGSi
j46k2hodJQU3IoJ9n+bvZnGun0FGM8K23VczA9E+mpa3DpikwNwoJgXmHCzt7WTFw2NWCkiekgAy
JMZTp0OBBAUNlAtbsblDM/CV3tGFwxJhS+sdBLs0lMj47zGVOodS/PmB0qNRY/Q+uf4ZagFdZaQ9
zv+qwP7tx2rfA9T2ZM87iUpclMFqJ3z6QpXa2mrexfiLTZJdYiyLjfBl4bUH5RqAX447cwywZ+wd
FtreX86keuRt2hfIzhW5Dvmw6iMni7CRj4PuDqaoBiIOCteu4fhKyDWMsjM6wLaobe2/cpKEqmMP
JglGrbP321AezYC9JVtBAwi/ErAPp0ixl3Tz4JTHoqMu0IMkS3wMPX6PzVjOwytJDcaTneRPAOVQ
nohTizUyN4r3lLo1OpNjuGE8kw7pH1JBOwVW+u+ovYUaBmIC5E/bljNNG0Kyqxvniz4eyohoh4+f
P+sLTjY68waaBv6Jsm9vJIxH+TWWN6v0yKIFPKm7ReVjpl1NsI8fLo6R1GD6popv2aG+SWqicDBM
lngH1Hpuqkfe+5Unp8tE1Xl2ya0jjSGLQhs56aCDuGEWRz5ie6qqE4s7/e7cC4NQb8bikgdB8E0C
4l99BmBvb7M2P7ylOVUkYEzqulc0/XujbQH6pehGQroljRm1975JAoO98EPrMlk8hoSwAo7fyWK6
KT+Ie/SlPcR4PiduK9cacOAp1LdOCnjzz3BgtNFAl/HmouBaQFINQxOQK1IFkB7jC3NAFtvCL2IU
69fBAx5TXbL4Pu1tgsvTWr0IVEjkRHhO5yxgfOjm516nCfkZKw+mkjCqFJp6189SmzxRw2RcAErB
Fb0TmWcK8lYVmk/NBJMBgJxdqtfjetlYUmKkbdxmCzydc4IqK5XHKJcC4u5wBd+DPgixKsRLOrgY
37U8UMXZmK1wq1IjMD6LbRUxIPrhPQdIzVHljJEUpkW/Ey8INZbk5otI0iW2Ln0vSBffEHJdz/iC
MKTzfsGzQW3bBgF08juq6FkCaHjZJ0ysjB5N/C0QbdMAZUXIU4CgruJdolscTXBT//uD/hjWDGor
Fv8DMByl3yuJxbm59Jlnj+VFvE9OSbQGi8jgCJII2Ox0SDxdnuu6HHo2WEJL5qUWYZ5ApVWSp1sR
+lMqzQgigcQGQTrEg7ptPWp6qti6RYmT7RB00qg83pRFU24pdww5fUJeH4pNl2lw+OPNVr2Zgm5N
zsBXIAhCrISmT7LZXt0nLFUJ5dhUDxLuV7KkAs2Zn4ILALJFpXXtEnhWX+uZJ7Mc5qN4nNWkZSG+
KPcuvJOsiESOL/YplndV/BTMKZrQv869VwxwvY6BuAkrEzXy6gf/uAF/M3JcIl+10RhYXXDnG0aL
0KM3+YVLUviqkZjLMVvOpn6f8cGLrqTfukfxVmIy6g9j+MopIQQToyuqSGsw037yRk9vdXcR01B8
v/tTcTqcijNupwASYRPo0+B0sUNsaFAp04ewnYcLz98FutG5tCxNCbeeT+AKy0wOwLb+S/hUPpWF
VvpvDRDipUXipN9zDcTB2BbFZl7BivC0o5AZnr0vrs0TMBrFXskQgLLl3OxIGf2LVX6AIKLRLPeF
7B6bR7jywupnMgmAOgsM9iBhSQlVKWpW0FKl7wzdpPO45nwTTYZQodoCvKLuQDBr7fz9exeBzXgb
Ka1iOr+u067WW+fLOdhmOQY4s8mjM6nbb+SJ8c/SXkQsSvDvImfXQd+PsnDrVNvCvy9GKdggUhCf
vlh3zrdqHmiS/Gp2tR8buZa0bCSTeS98QMbB+v+ZcyeGue1VF1lwLVAqZtkUAYhkB0uD5jDQmw6+
YHz7PclSD+KVoEoSW8P9xeAsy0HPM0PtDj62bDY/dtvm8AEO9l2MeUGgpcIgjK4Q7YTgS5gciOwH
DjiG8FsD3YigbQfQxNfyJZ0EUTdLokmaGzhtQaWRkI8Y0b0VYgWJ4h6LeVVTG3YNO3RaMeOf4gfW
pfCLz4zxOoAmrpx5lBnApbs9EP2QCp4TBlLrf8IORsMfbiQyZmHzyJttYpTIketzCNsCvaR3SfBx
XP72M4S+tj9LhMnyt5Bmngt8uQE7vYGzYKOxc6gqr4HvGMG5dpDepe7DRL/wqcdOvdxsKG8pFSAA
esLf20cEy6bif1MxyT6sKBxz5Mgf9G60ZrXcCr3tRbFHWivMq64rGnlWYk1fYxmhMCQdm65YuV8s
5Bu5bcF75fLqjrjdjk7AojPajVYOIzZw3C+ye/cssvFurzzIJcJ6RmpBPgHr8meC01b1NtTcYmNw
kJ2HHKStyqPwSDtLCF5YOKjZngohMpiS1gAR+hoW2ozgqbMWoAmXkXAAVQY8cZkKQD0mSbJhlrWc
KQbcOemHqXwSaepTZhU0YarKODhK7h4BDu0831NZLG6cuUnhPr9pVgH2eHSLQqfav4V72WCjGEEu
4BmLzjdsynd1QZl2+MGQQ+5J/PdDy9lEEZoP7UC6zi6meZ0utGss9Q55DY0AfcZgao+d4hm2M93i
t9nAfBo7Hs+V4Fe8Xgw+FWovE7eeTY4Y/ZksIKPwEmPxJNsYVCFBAX5EYCWq2OF1gUoPicuthgq8
ggM1KwXHTZOxifJFD0VxLuf5S5PG+ATYJJ38XmparfVO0azA5qRndJ2PjBnjCZ5HOODDw/QidZxb
iDhb+2epmhFD7OX5Ja0s+whJ0d6Mp9h3wUxAsWaxck7NKUEPYswwGv4l+VXkPTVpUl7Jg3mcUtnZ
2GCjP/LJMyLefVPFhuC8RnXYBpiPncJEqrL8KTep4q8z6dvF3HtlhgmcestnQNM42dtnStTXoOdE
+9euFXd6T43XrilYIto5x2P2F1FCR7HEf3b9Qf1dVjzTW2lcboeGv7QO4lGTv48I6Ju1yoWQm5Nd
k3Ha67wOwdBW034ez44/5tV7me48li7vOFvSHXl/NfAxsly677+azFssCvZ3CiRlz4vKYQK5MAmf
t0aeYfW/r9GHK0NRupWgVjyWTd3H70tquXmTj8yRTBR8t3JcwXDhsNlohfaA2dG/dKU+nsUQZkGF
vu+F/1gtC+LoGpMghF72F/urSDdx5y7O9Pifx2wvJrAvkzZ52ihKTl5bNXq+rcgs+cxtxLKDPJ7i
kLWIAp/DfSUwq3+CWOn45WA36Gfhtvee4PFUr+6Cj1gjQ7kCwPHDsv7DnTO3QMPqlUldtzFORkjj
HZCCSpf2Sk5YUdUHeDo7Di6wft2ppZsoYPkQv79AifXhFmbjl1VGvZTqXpTBaT+sf+lN5nL4s1tz
kFtsXjDFPgCdJue5kRWPOu3LpZT38iAMUxnwEm5ZifuYJdSpBLCAaIplp02Dg7TkD69UhkIflWJC
xz6kfNRl4a5GtvttZgZNv6LOwuSzq62qPPZglVvu5iVu9LcTkkPmJoEk1hkiGC3h85RfzgH1aTGY
0/vtkVaFP2ac9oDYSnq9qPKilMykKkd4pkZbvX4qazVX4v48Vdy5kDPNIcmsByPEfE4dnwEn8gcY
jyiPM4ZCLs5pHy7BJqk4CwlAiLUk1aAzPacQ6EWsSSyABPyio7cqTZp0JG2MF3hmaKHPbF8WpMEd
D815MdiH6HjfDR+MWlkBU+JwgG2OIpyUpRn2CWUKUnWEINslZDJWg8h9qs2fQa+W7JwyzRuDTDOZ
gKu56qJG0dvHvK9Hi8AV47QoTb5y7g0RpAcpMA5LLf41MBZoVQOAG7zFEaSqfTb2ee2zfVMXHkRb
VqJad3PFtke2e1V8UcLJSPhkFiGNyI6ZFi4Mu2eZgJ3/3Jy1sZhk5FKKlMLSlqcZCZy/xfEWWlV3
VDnBzoxC4xbK8E9VYVjzo2qjhg18uaR1ZYYgDMK9MfdZ2lbN88Fn+MiLfWUyaDo+z5sHiPyI+YkP
cWIINWmjcMwtC1DatoyA6mtF7eqIqSBXd4UieHxbuVXP0U9331nPVyucGpYKZNbvDaTeyLWCD8aM
f7FXLBHPAmW+OS24MY7/OCCn5xwbzyHVHaez5m1Uyho8pDqfuGBY5YMCTUkxFRg/aAGxxgzdj3fv
bPD0mFvACHdwo6GXHwXmCRgBMeIJWxfl2k/Kh2q+VS1KflRRx3pF7zVxIyMn5wH8LowfA8oT+G0c
DyHde9s1yUTk5Rup1RCVMP6TdirZaZI8ZUPKgpKi0Czb8UPODLjPTk9vB/OHrYFDBXcXeWmrl+gX
mS9SmomO116Cnk6fG4eKTFMf9jzkRSabopzm6v7WY2M5y1cdl6k20DhnomDBGXU/JoalEM/sHtL0
nnENB5PJ8Rzx4zCiUSQER2x8tBeCRxDwgFlPq9jz4BGJ9pvHIIz4Yy0qStMGlBGYQ/EzHvlB8j+o
yw92NKCUONZiwDvtrFVJAvXCKj5goY5ungzJiEHT4ANCD/P8mBpdJLfXwpCxxMVBPXSaRHWOTrnW
pM/9FTVt78C57oR7SiEvufGI9WmwUnZpBxps6R+KCtp8VYmi2qvX1swfXpBpfU5nQBGVOhBq6p7z
h5zkHPEtubwDs3QOLs5l/pv8i/FlRwZ/E77yubUnFzLb3I0mtC5zTLNOT7F42wlPBf9Y3ZOkc+Uz
oqttFWZvVMnaS9MuJ5C99j9q9hDFOTgylZQvkPV96+n67G4aqSYMUaMgZZwxnuZleGGe79f6NjNI
8EALFL4KVkrsHwKGy4TdxKx7pRUQqMpKO2ym7PRk5aXt3i+Jt9ea4HK7WeJHYK7akzJoritwOWTj
htiHmSQaxg6Oq3o6XCu2L2zslxxcy5TViUJPG6haQKGl8X8Mo7nS5XSuWYQ7nThNl799olKVJL9W
v+omSTxcw4c+MGkb/fEyrNK18s4SvPNvHzY2XcHmcp6N6Dn5v/g8gxStUnrWNOgdz7nHUZw2eoJr
ZiO3LiSs2NY5PbT3omvqy7IvV0DIw4wjiAC+R1Er1LjGg6okP2KvHY1OkdfukM13iKcnog2kaYrt
e4A7R0zpRWwdZp2DQyMC4Z1XaUBVIvtnvlrr7TKeRnmt/rOx8Vf52wtsD/02vW0+8ps937HSO6go
5Y3B492h6V1Gikj5Ab0hCHVy7V/A4dh790kXF0g0rk59PyuvmQIPmG9T1VC+5MaZljXUYMh2hltz
UnonSah/daMkgAE7FLg95UEM6SJk1YtyoITQBDLg7rwLonrHtCQ5jSWzvVkS+h0hvkW3GRcKHM1i
mKcByjc3g2zJruXBO0Cr6JD2+rxuy+Ta0bJDmR5RA6L8Mt6gm7UEvpGBRDZQyUrseZl3EuyxA/+l
fq8kCfc1xSLnco0DwUwC5vDLnZ3d4D77MM0RytnpkqfTxQqwS8NwnvChPi5t5tG76gHh44WA6Xa+
nqThPy5Z3TMhdgOPcCg1n5/m09qUgsYPs5oWtkmJdSHHFUeyFa1QsDDobP7oR2Yx7qZF4uVZsF+K
Bj+jSt9o8BBO2nMgPtp/4JQvzkUbxmAf+/sXR2tmnrbwyxtBVLTH9b0Yiusw3hUcLYW38AihejxC
hPJiY+RYBQmWgTWOJ9ALYhHOHEP2xGiA2wr9dIwx6RhswPnbxy1Sbk+1maM7bBjomquECt53MBlD
zapYIs2lJMa7snuA+SEIlp2UwoAHbntXueL4ALWvOqWKtD5Bd0lMBOB/tu4aulmk0e9zc6xG1I+i
buPybydN0IedXlDmVGLd2VCR366Fhh7g4tvadFJ0vRFhwSYPsau10iudx7I76gXthzwnPtY872Ln
eJrAS3L/NwjXFD6Y1RGVYX0KCluNagax462EzDdm1n/RmcOJ/8GXXiNvzppCczBYm0CMV/9RArVw
npOHkKk7nXX6k3W0Myj4zBRFVsZFsEAcZXlcmsDtz/3HWpYEEmCiJjvo7tN7vtidgzF92fyvMQnY
aiYOXj8ZpiUFIFXFw6RciVdAqOr6La+2Inb33K23imlxHmG8tif3M2OSa3hh4L5p14h5LIlLde+z
XP/scoaegAgsjS342x/kUi0MMXq/GoUtc3JmmPicbMUUUvqmI+KPSEgCNYhpPGVTPVY1X03dXBtR
gAGHuENsi34YL40fHze+kN4gkgH6ZAJQ3qLqoB4+G0u/54XJS9bY8zMC2kQmoaE0Mi/KSxXGi4e5
UqaV2f4mBjX5DG7SaHY5PyQCLmnj2X/adhFEzDJOzuzWJHNxwS0OtvTsftH/GvGAbJcWVtK53g6Q
6FdNGb8HZPHLTDmA7bhzWxuKo7ccPtoJdUDAg70sLeUGPMBRS98nx84HWiBljwBUNyBbve2PqGae
mmauCmSuE0BAcc56rDcA/BDl/7XYg5V9ZDXwWheWHKt/mrkru6reZJ3QkyJWnfJCntZaXLKmrqiP
ptUixZrJ/NLb3aRim56C5wkN9QmRruGffefWj9y7IhNK9TUCnaKtGyGJFjjlkXszcLhVsXCpNtrE
krJnrR72j8nudpoTbuUU3WxKpUD4FdwNa7fKIgW4h6a5ws+d0z5QYHPOgTOYXr+lGWIm97QHDTMn
9bQ30UU4lVx8aHIxaORaJmu8VjP5zPwl+L8ZBFcziBEv2U57p4/MxkgWqSgxF/h+YMl/MvDq73u6
LEteMiuV3CJeZxEp/dSBaNAaxeSLetLij9Vg9SVQZMepqrUg5ajoXze3yzQsLtUyQGIVY4ESdqqi
Jtu5PGsD+YBPiVA6sTqVXO0ifDe4WYDqRmp9oiHBD56FkNBk+kxVFKqR2h8PBN4AY7dQC7oNACZD
8qlj1U2D7Gc5BfquWPbylAhbh+nBSfXyHV8ldwk1SmzUa/CtGtWQpU+D4PqKMvnbBNKWvwAjh58b
vsXrhfIwlRUxkAwsxnhbhgfi15xCzgg7Rohqc9vTAAkh9je0yfVcdVF2XL2ORTW4+BET5JCcsBBJ
O31x1zKZQw89iO9tYRX0m0qcM9mfFqKQcCMHsVfJjTW478xiVK6l8+S93FS/vT3U7QLmZkBDaJvy
lCHW4j6Nmh2SrK0QtMAwvOuZlCZfsj0VG+xK24zQsvqnoBbG7B7B3HM00YlpDiPMSHFHucarFyfo
NXTXSZMak1d4sFseFGHB1ZJKavc4YBvW3Hok0xdVM6Ot2piqYLazhSmRvEUyKSeHdgH54Cj8h3sT
ImcxYB18r1Q3zbrxZj+i/RbtQPV0tzH1n/mTGYqft1xPhANZvxvdxacSpfdAMsclKOpIimeRN80d
zVaB9EAbOYKg4yi9K/J/peLsWWP7R0WbPs8FkCx2HhYEBXykwtdOwvd9nPlpEhUaa4oSeO3oHLf0
LQNs5Ss8ZxtxmX966efwmntWZJ986SxX3PFrEmoybeqIZdDig07+CsWKhvbTAJdFwBZ+zqHU0jFM
gXWANgaJJmfJd5VjLjwgwu1cWCWsfjfTu5sAQRGVsiiwsBmu5gSd1r2Cad8xD77bqPvZv0tyMW3Q
F0dvB0hbC54EEvDLZmG+3t0ePsqCWk9yTNCK7OXEh6QKs8y5qkzG7qGtb3a9L2P23+6eZoofISmK
j4P+hN/YST+GOqVYz8M6pnHtyhSjjK1IUGAVr3xPwfCb9yloicGgxb6c3qWHslNU9j6p1J2Hvs3Q
ppY5KFzZ0M+5admE/zK4MIU6X9C08DTadTns74L6XMRzY9ICPZayRKuRmgVLNHaBdEz1MtYG4CW/
5zM2HFp7Ob+ldKmTQIF5NnWdFryW717vueRq6tVaTEtUVrAa80Y7nly2niaxjImZgA7l1alOXo+D
PaPdLcvS5KKUiaCcLaX2ChWJoqkLQnJNB8BbI8W8yb/J2govYCMUDdzLLUNcjIaejz7J4yFq6d2O
noyiCe0lk4dw9CYitKFSlEUNMx09B7yNlqOXvnxKKDgZ2ErvfCMMuV0rvy8lybBvS5+PiBby4wEx
td3HY4cVi7OVQXi8ig3j9+n9aO8uuG7jG5G6mC6NAZQNsb9VZ+tjjuhJyJ/8gNFzf4mhe3dIsIev
HYA1L+FstqvzMvebQPxGRA3ccZq91d4qmIRAAe3eLg3t7//nUsXPnrYIrrHc2PrnNYRqHbM0l44A
zJRUClDiy/8eO6+er2CnDfG+uKe5V3r1YoPnMsRRuR0Rzd0j7bAzZtKutEETXwBItEOG0sN93fxU
AiFKp+e8LUsi43oMHlHRFc37V2OakrdJSjH7GlxKZfokdfZtFI+jWPsHAqbTMoT9KOzaCQ9gVlxs
Rpe64GzluBwRhlosvQ2CzetnucPYh0VTNe+E4X9/UfuB1n5oEhMkz3euFMUv0rmoG7Sf3NHmoc4J
VjEaCbEhe+Oa9+OLjulhEBkVLegLdGB+VbZxd6OC+0nk+rlUO7BZ0PPB6foioOm9LY/q/6Y6NBCI
Jmzzmz5Ot9ZjmEfUCR8KdcyMfZU0TGZogKs3CUTLX6IVMgWDPY+amg2qNwoTAEdDPyduFF/7YZhV
LbeA5rfVNgiFTLPAonKrgt23EFijmU8xRgVia88utVVlP75WruZmv1cu5F+H/VEcZrtxr3xoe9gW
lX/X8oZApKuzGGNVxiw0ZV7Fu+45Szxplx8u2G2TlEnkS4vJExs1NMwKdEEz3sq6o27jvAiXHBkv
pR4hFiAWzwCs9nmedbv6CQZxZgVZyUrI1xoYjYGjo+lyqzDYr3m1cKSTHEnIRfMVHc/CGopZ5Ewy
LjcOTi1lyYMrguj4iJc9bV40OZR9m+kRoRBqCPouaZc3GBj9zKaIyVate20sNF0DGQHwrUiq09MC
mQeyGzjVaETxDZ+HppnjjzeLTI00qBEUYIcIw/RJO7GfsTv3x35atTpFbDxY0QTKWmDhJswsVoO0
Krwl1N8AobbZxdAc1tF3qUmI/SLFt1pYjiVbuAee33mmHgCATgXPjxUV21rCffSY5nvMibT7I6IW
KnkVd5NutSRCMZNLaVIRKRrs6THNO3BSzlHe9SBdz3MzMMPzG+Q1syQ2cKWfeoudHO4o/WU2bfLL
46fj517sm9AqOTPSbCdb2RxAIu6kjoq6ockIjXpMlt1/ZRXj0qHLzs+1LaGK/w/t0t6J/RrqYG0x
euWNLYLun86BDQoD3/FghKDsuGPd5h0oNy1dhpjW0K8xUv3ZcSpHeKzm65CMhECt4ymPqJHwWQtJ
1Urr/DRuvt6ppjJFRr+PFPcAvZUWKifjlLrha0bSOcswxy8zKRwA4Vun5vcZZ3HBaQBUn9hQyCYl
EmPnYoD5RfzPtMJmZlDCewHwQrzkmmrhdtHHfg2QDft4PDxef21+Z9e4DnMMZkxVoByQOgms2g12
BzLpJ0wbSjEHlmY0UWjJMqzMqp93EpuxECsgibPGMbglFsfqP94lg9HSW1M+iaLNt4TGtLW8yo89
IBwDxxwMnWm3yJGTydzKjlZFvmfEh2mEy/Y44X7kubpkdTaFzyKrI908zi1o5FlfVyICmxSWLFac
RAL3ksWFUOGcUkl8ji92n1GVL8rRT0iVRQu7LV+eksoeqaVYtHhAAQK1b+Xc+NHWb6d+CABG+1Ip
lt4dyuOyYK6lHD/BnElLig2EJ9w+Cs9qOSSMDVmprHFKfaL/aisETph0w35m5O2mV6Knk/KlZ9eL
48VEtiHe5RA24vMIy0tK25ylgPOTsb6FuctYbBKKrnnDUOiiHfvuPqSv3eyEKa9/WvCcIQKVi1XG
6T7FwLaflKMkZ2JRj54LMUkzdDfZ4MZgoDgu1fjZduWnwIGcowXWX6zzr1AsemVxjXRWRbJFuuPe
WLRrdhjnVjgIgQpbhFHTo0mBYnbGJg2mx3oka+8hdtyxzmA8SHY6/ROFS+46phVxGBUG6oxZMzqm
x5nNtca5LsmpQL+kfG6pHKVGRp+YRpYb+XyU2XRTrzqWElleUkcwYSFiHy47B4S3BuzGP/V5MEdf
3cFFJOldwVXwj5va6DxCpc+5/o/iSL4a1cMHT2w0pgX11/J0MUwkocPIM9gwKP1i6CtsSj+tCZEP
Kd7lByGGvmq28W4MduNs/TqOBSX6tpudOhmPBEVffa/jBj0GZI63hNhbt+tTzhHQ3ZBj6jgVy20/
z4c9ceoOgeq1gZdKRc7c59A7VrU9wCJHJTQFCVBpJ8KO7C0pO7gmSy5r/Mu0RCN2Ng5dNs3aBRXA
O2LRffpnipnIelWlcX05jMFOIVYIWPgZ6lMufunZG/LSsnCZUOqUbiCM0y5szH9St5Tf138y81Fr
YdFU24jBLWv9+BaLmx+USrsoNrG19onCzPIN7upVrGskHwOOXqpws+0mbcZxRmTL8W5fRn80JFlB
AVsJUauWI+rV9Nk/kTVpuXjACaGZaD+ionCIEWXkh1AHfUCH6zv7iCUQUKncHP5UAQWy5IZ0bMNP
At7f/C2cX7HRBLmFGgSLrqkxPXcpQiJIaKowPMyDpkfI+2WG6vTMm6SaItzBP4Qs4AzV4C/rOcGx
oUFITj+KYxE8IpY3pXezhZQLpJvnTr4aOZtYsB4VHIY9CiAXUSq/Oe8vVWKtuJzRH294+mH/fGav
x83MPNOQHCpRjx9A+EI5iLnsb6vs5RBzK4W6HPEEKA6G65K8Am99e291XIkiQzLnvfTDlJl/zE6C
W4wK/p4E8DlaNfbQ53sxGKgj1H+RIVQJmhMscS+nZm52yDcDvFTVYTf5bi9ifzUeOoN5+weUgh/J
opJqL3MbHk9t+nlsHYc42OC/MTCpUjDPQ3brGk74u1slzcScrpJPDc5zMD/dVGZk+8p/pXMBEh1z
p2OATYSbtpMlcUXDuKA5fHYBXne864JWM5SIbp7E+rrxZ9ZECVrgV2mfWfzy9nkJqcJlyTDduIaw
FZ4OqcOZOtWkQRM3ObcRDCf0O2DN+onPCcEjURkxs+c0edui6Ggf/Cs0z8Z0gqPjpGTUbTLDFOYY
7TL7UhrGFt3UNU4H3nzT9TqEBp/8MiVrnp52w1OIMsqgcDNHBBiiITCx2IeQLmbDXWKqlWIe9OVm
6z1KDdst5YuhWd3yfF9uSv7T3DUMLzpCjRYuYFWo6+8BqGUmLR8eLSWFvCQCFpLd7czaZE5phAGk
EmXw+Td9J6UseVvVx7cPWt6UHtiZ6akQR6mDwMKbbWXE/ja3VEGJW35WFzunr2c12a0mtM0sD9zV
KjqX3ELXXLp2205DW3GoC0VtZ6pE+3flhDCiyIEfTwyHajXJISC1Is10bNj9UVabKr+Iup3bYB2X
7NOaRjmctO1DuMhXXsRLK4CvfCGKg+APJBK3VAY/N7/QXSrxRzTrPnR5qPrhHM56o7moBXGE4BxC
E+ye6gvzyIV+bhcmW9rh+Xw80Kv6o5wkmLqYp+hwZHuHxUY99ZNYNjuPg2Qrbv0CNoYRX08EhSfo
MJeovoTkZ38Qpd6A+dQB86qVnEYRXgNwm+mNDSYAdkOTSULjcT7HLZ2m3hadYMSeIIP5TA+lAzXw
h8eoGk3aFSV9B0ESODLnoyeS44QreJF2fYO4UbxCxb8HfncwI99ARgy69sEQRaPTJMhqQft0H8ae
64c29OZRvufBpacO6jPJnRKilr+i3RAcUM6your7a/LbMX0IRp95CbcHwXvRkCM9zEYhbNZIl+aB
Pmq7/Ci66k6r/uOjRu1zqXjoH2c7DS1CXuvgnmTgYOLWJjrfg9HWzNkZ0RIyiMK6L4g4GZ/66fRw
K8DkBzbLSaV15j5vsGT4xSE5HOUjUwPDanoXyZeHKvdWEnMR7yoZvIbPdKBE1AS10LBy55dHNG/y
9ZcYie6fbfh3vYAU+u5i68AWlncYjOXHHm4xite+juyTy3xZvOyqcKx/OnRJAtZe0mVhrsqPwFVE
gYm8YyEJwHbUEGezA0RPQPKEGC3a2Zzt0VTBp2S1SUinlzqAoXVrFtWjlhBYgxxW5E6BwkvhxXUb
RMka9eeklHjNXuYYPA9tZUQBZ0PlqwvBAuBPHKb7d1169eRDkiH2W18n5ii84Kv4iqntmSlDxMYE
9qNgq0NA5uVPg7XBRAQI9KfIdZB7wHMKRug+y5qdUnToqginZ3QS4PCJ/cqp9CFzc7Vlv+tg5iGp
jT0htnuEP7lp5/pGZJPe25241iSE67aGvZZUJbDExluY5A+4Qcp3Dk/VYthiL8/yaVzoQJqb+ITN
s6ZV1dEFkayaarXYEdW123ouOOLn7JyOsqdwnLH0SCP5xvus0n5DWWzqZ0LMG/kyWygU1GP7PQov
gnVLw82p7FsPYc0x4m2JoTV2qUtV70573n/m/oyDGcYibIQ/O4hA6OzErOzLlukcPlPnoVbFMbnM
W44dmVuNMV53BlFHMv+awDukrbzANYD196p6aMu6N9/tdMPJ2TEuyJDlvrra48oK4pX34lH456YN
h/Gsmc4bXfzgX76e5FdC/8e5saX8yiy9ErdZSm6VNooEgowTEt4xNs+9yFEwMnUrTJgnbbmXhxZl
q7CiXn114wR2TK9EFbGjtmvULo32F2ckXqmijSea39DeaEtkyFIWM5axmrJlC2URrn7F/rv87VkQ
E1ungnRTIP8EeUwq26Msh7r7LxRz9HCPU+ki4Zk3FAHr4knTYcofJji/BOdgFtWLKjiQ9iOIKiaC
+fQa9UQLk4JldAUgJCsbLs2XdR7r4J8c1qhUvcSMXRRihBxyw68msxWnoo1+LfWWmIejatkcShso
tDIMdgsTZse3UfN1sdpn2KgnGoXXz/3m7nc6h0xKq2Ozonr/A0wFKogER+0FRpH6zo9IX5Q8qDeu
yiIvUe+syL1QLh1H9mkvWSVIdKSg5SlYVOsYy/eOic/ZN8tYpRyBdSHBlGYmaEzrq5ypf8U1uMAH
z9d/VGQlDdUQLhhfZQ1oq45Y28fyyDTP8vibLoZSY1gql8weK+OUHfxRum6zniTdWkyTXM8k9pY8
cnRMDFUAnN/oFJEt/oaG5AxjZSD3soHF3CgcmRMn7lJeCzfCeJE+IT26b4aU3u9SyBzt2JiMsl2t
XjBbmCutrFld+c/1PCp611d3WyAlCfcScCEynTdWEyjS9ppzB/r+YNq+0OgDCHVPO9qq7KcgGMtf
k40hc1rUCuyVelhwX7fVdMjQ1VwB+GFDOY/V1MoJB9qOZ1fHN75Z/BZEo7DgcTFogHbsfkn92WZ3
9OfHKDoEqripcwO6LsR8ubRZ6RoPCNMR0lulbt/GK0KVwIl5+v2YZYX04Av1P6FZB6sOa6xqlUkc
Ag+NN2uVmfLnaMsX7WPl8k18Zo0UgmwHHlw1dMwgS7MsLkCEB9tzMXbOE8AP1BjXWUj2OyN/E/ub
UHvyMidAm3fWdY+dds6nKmKE+Mvwt5kyiq/ePaI5V1p+jO3dCA6bCp5yL8DlwMxfV38frazyEXIX
I4F5Ve1D51ggvRI4a8DBPsYf0s/lFm6EM8r4lxhsAVXuxg0LEAhbOvJbKzYMGWXFyQSGITFhNaqs
oiJyptdAcWtmd0ZZ53PR2pbD1i764OiJU3nPwkdfZPvWB2J0V39RQxFxCVJRRpQjHQuxcLi3/BI/
hFoj8pIWbTJ+5zxgKU0e17fguR0l7sSYAPRT3eNaceHehRaBy802Kr50P+730WfDQwl0Z2P0HFsj
o7UOLfpHLuWqDZlYpGRxlWPpzro5nA/WMvtXEkNk4ntGIoOO+UK2N/YrXhgYb2e4Uy0NrhFPOW/M
+QVd4ESuqmvHI0IW7uPOgr18XD6EmueFBMU+71ZKN7gor1kN2jCqrM8Q//3AGZcD7ICxFSz0LY1n
0NQHkZw3F/xBCXirarlN5G7o0tOq2metD7kGYuz7y66VWr0I8q4lnZBgwZEDV9O027H7umA0wsJg
TuD6jiSdmIrBv/SrZXqYGXrDkNkby8kUwnwrrqRmYFDz7UzRwcquUVjptccSFTp33/XMKhAxqjcT
E1Koog7hTH1Egrg+1RRrlKclGRPIewRLdqeEu8kGt66IJjtSF0eRDI6DemoV8gAbXroJ9P1E5Y6e
+dLdz5FmzI1CWyPz+l94cdLRrKIttCTZFCse6p4HbT4TP0htm5Wq38hatReO8Yl+jOXEhJbJc+Qs
0DYy9QKQ3En/1cQlKcPKQMdNWs+t7AXsJiXyQOoh7E+ktdejnQHe8lS1XcH/IlJtx/opShGjm1NF
92yufm3kLFf+vs7g3F9LFK7CPrUeQes3WGK2Srky/Mhbf8WgdZB5BmLEyu6rs+5zW4/seEyzGdMu
2B3uCjhu0dBzDETodOLv4W/bgsWyUpTj+DsXme5XNn41rufXPJxHo+QUp1d/DVdVeJEJhRCpljB1
a49Obo1nH2OBAkY3SsW18d9UwypR5RWTuApWy6X2vEcdNb6AF3/XWmMFTvj595HpytWSq4K2b6CE
bdP6od09BZ5uxPjDeIGsxg8qNw3MgdJtWoDQ/YezG4Y9xNG+eK4vj9hbX2lzVtCkQ94Kt+9d5YAR
BnMXmqr4tyMFyY4pBUhZwqmetLvswUaeVbCAqpiuMVakwJ6AxE8HKIFZg0X85b8mhLXi4k7bZNdY
C2CdQDsxtwTBtPYegjZsrTT33Hd/EnjeNMP/JDa5UOWYhrwXTgq7OXBFz9+lGDSVvnqLspinLjK4
8U+MCiGhbaAkkWrRvMChPjTWujNmW/pFQv5YPuf4a1RbPOWCMKeS0Bxlnznm2gpyjpOk8pjsYkCS
c9+liMHSR+mBieBwfLkvflObhmck/aPvQdtKcekKSnWUdOOJWNEL7+jF5zsFRS/dx1wWW5v+slTP
8rnK7hg4H/N10dE56qif9v4ixMyE9zETSHOR0MEVADdKMLKO0Ne1rDq5Q5aFGUh7wlRdTmcDoASY
EcRYkWy2cZ/KF23KTeytlsKFLxoJyIT2YTvXdqg2YIhzpB162HPrGpVpsy7DWM+gGfESbC8CHmMs
JRjBXoB/o8IC85fbBbLA8R35YMH2BV6LERira80atqkckWyrcU9wJ9ABL7zLnzlBimhyPZrxqNJQ
ntLp8hhxciKDjpLWbck6C4fqwe7/sxrU+TSAs4Ub0YoYWUk0YlFlj+kWhVeExubGeeC2+azZw5+Z
TeIBXRCeK0XnvPDIxHu+wJ81ucYQ7ej5x0bMouZuMXlFUMfccb5geSYerswxfgHnKbTYLNc3jPuq
NQQJl5uvAoWnD4Qy4IIqhbnwxNjp0gxylvSLB79RbP4/kv+XBk8z7UaT7t+XjQDUSlpSMF5ewTsS
WWTY/7GwWdU1XcWLUBvJFNL2/aXP2dEymPd36rm2r9KTOS0pSEf8mdc8Gq8Ka7LJ31YRWhU+eXlc
eKhKF2RNc/wkgsRhoYWb54Jmh+OjC8YLqf3W+obU2wNGL84uWzUlNiEVTG8Pr+bqzwm6alhr0fCe
0cdKeLFTnYh+f00Dw95BBvYAS6jTDKhUPIsdDTwBWRHMNUqg05PUiNJBamS1r+y6Cxn8HAGGPPvv
Vpgkp7A/aawmY5v+qieHD4xocNtFHTjh6xAEQQ/SYVa2nvvJ/hdjzAE4/6a3kmxhe6JLVeAGV1h7
qJQUonS2lDPksLAQL8kbBBLDTPrtzHRQDQNvIMGqJk+LRqyCP0AmTF0dSeCPHVct8gq3mIxZlU+T
GhV4TF7hd6VgNf1z6pPEMSs9BvVMayYzPW1lYxBk+/ukWg3tUpSqX5jZQRT/AFUniSIQl6M7DE9Q
d/1pCosti09VbaTyzQ9dTRiTRRJFyTPhOoXTXLjn/j0ckFf/TodrRZXW2vFiq1CWafv7zHUs1PMA
YWZbZ4qRykbG7jMHiq5RiLBebZaqWAlZLYh557iCaRgpETAQp47Ed/f9xA3H6eWOLjqRVRvfP6PA
A/Mb75swM25uXMl1XaHup1Jc5ji4zGlKx1D6cUC8HqlVMZ9lH1tXABWpg0MFvFRqOAljIf2fQ83p
OCOn9BSPfdq5p11a66D/tnFIqS0jQWnlBgtGIWLKRL95DE0+NiwcI/sqxN/lZUGMbGRVghGq+VCM
nqpU4q//a7q2Ufr5eWSp9kcDTXzRuq2R86W3Mna45iQpZNUf2nx/YXOKBFMEDh6md97wzGXU68Zw
NFMOGFcE6xJHpBjdt33HOd41cxVRW1uuk01w0uHPewyaSsjNDeqQMXx9PohPRGRulE/xVA13jaUN
kKkE7igSy54QvON/O+Znpo08DyyYH3Hm18waitp1coD6BfSLEcuEXIMnAtDHovzHYJ7UkfLGHNOF
zjOJSILVZ+t2zv6jH2Vl7SjF2u85HXVyiDe2a9bpkb1Vttv3hrZto+yXArajASsfchf6+5hwlF/n
3+USHbqmJ2eLjxw5HHvR3CDcXq0moxSl1IdUe3BuTvABFgCBph0y8x4z/36VBreDdZBlMH+hvH1Y
ii2Y4E/85/3dSFuhW1gBEnxFV+5v1hohrkeLzL+KqMEpg13AJJh4YCwibcVOM8APISPrppBzBJQd
mYu7najySyzlGjeHAS1qdyV1Pg/a0lSUng1gJckDNfCKmdBDRsTEP7ioHYbfIxAtgwfRpjQa07df
vhEHwHutd0QbGNJP1l5UBQg3wjukmXEoLIDky+2PDbC3s8eCznvngvXqSQe9010X7SCI5Sbk/EvU
S14s5s6k6GbfegzqXqYRpxYHm2GGAomS8ZaCR6wPC49Hu/LjhVTAT3ND4neNcDutuPN0I15iCkTW
qbDeh3gHPWmy8R3kMqHT8Zly/zNGUrMxORh+Xg0CXMH+MFpCBzhATItA6wCjXzjiCIAhvc1TspCJ
Rca7uJ92W9fHnr9CK8AZFub3EajGhNEGxnF6riYUc5lY71PUkzw/BQKeK0lgeTr/ShVMGAOm2p6i
j2pvMldgnhYSKZTum+kaanNWyUJkjL5kbmCcIZ/vNH4G0YNKikcIKUh/ldwyLB9GsyjvEpX19vTh
qJEb1wHBYR7QlC2Pte87dfjvV2grlVsq7eVpRGYgs9oRc6EG9BtKvwl/PVAOLqf/3yeHo+2uBJ1l
e3vgNblEwdwpey6nVwgaZo048oDH9/sBTZRLxTq+SLUUz4QZca8ShjQ5fB3RcExsYNuUS2X9GfYU
EVtfrh+AqbaR8PU0psFEJZDTv7VnC5cFAWec6sNOfk/cg70OwhDzpeRShzI1RW6h4C+QbyKqyO4+
A+8lRE+Qr5hGr9lkMFAxQ/fmUNEno5u+fHl9EfVhT/zHl3jMH8eh51YVcGcDOnQRsar6LplqEvo1
BvFW6zTqUUvyhJRNYnPXpZEQ0xFPVUYdSySKd7gMlgAA11Z5de7o8HTbAf14R6I7BhDmGaAeY7ue
IDPxIEZgfk0uuJj7hj6FNsV7k5S7fNWFXe3kV80TCQx7HetHRdzOe4yRAp9x6aLo7R34dDn83vt4
dFDNingPSaOP9U+nargN+44/LMsO9lim4HHpSawHadR6xAx4k1X8GM5LCyI38UTidztP15MG3hEg
CM9Duj29AV87COcvUJmGRxU/gdWWPaaz9yN7PrKX5PKVe1EiMvIPCm9E5tJU0mcRet/utnxP8kIZ
PgYy6QdjDU1eh8/EyVh0oBI9jyrqLUxcXpO5VYBtOGTNSzfWg+ufb0MKP24tfhnz0rAZp56WVDCN
mdh4vdtyXhDI8MjQ9kKO7w4CvJItyXtaPM+GEIRLopsZAIgduRZGYpSXjgIPCd/mCFfncbwL3IcJ
tdcViQGER/325vTr1U+cYbkK8SDqg591Qh11fJM0N2OEcdXaNP2yCZZyn0tkQWAlScflVvvgv2N8
0RdJVWScSM3/5yVmnCK7507pB42tImGb2erqLRBCcbl+lNxCd9EzNZZiLQUsvswn8yPgcQeOZi2P
xq+3XdZm669E6xkk9o7GywefDWUZNn2mIEc28LcgAP5SyLhoc7duWpnyiCwhQnDVlxqzS06oUCpX
glrSHuwwHd3PS9NidPKhd2/tiE/mhck17xfs6ttHN0NHev6P5JB/2VroCCOoJYnK4aOdsNv24ox7
TkvbuSGN22hgng3/RnfnAu8vHE3kF3hKRWNxDS19P3db/dPj0mpjHYPEJ4BnmkHrCdQpc0X55Jlv
EB/IzVKetPceMVBEPnMqP30R3Nb/PYJmN9h0f1kMRjpDMQFGHp6lwBE7yPSzxq3rLfmlyqGFhEA6
9s6M0Ti78QwErQGVxkH6XizOEu+cQvHTMUgsmqmgcvyg3rA9Frm/28L53WZI6rrVgT2vorLAUbXa
5vjfdgRYCE4rBgTVe6BP3AsEjn1ZsI+Iw1pTbP//jUHKsFUCXkIjtsmfRGw+ffwN2N8G/tMbvyw2
z5jRRlctmdGKZyd5RcGtelHhQjMb+GKWtDarrJiA2r/cmHIRq/MEe1RLvRUyY9XfsOrowUJt+UtS
LDHxuL1wUjKUuYaE++RG+c0G9NY1rNjt0h6fE4sXUZaxxgrOF79EQFNKQHiw1RBIwW7BJmchBxBj
/3K3LqcFnkmv4B+xatHJdR910hJ0z07shXobvshdV+afcuNmk2Jxw4gC5gBAs5rvfsNh9ReKu6AM
mZTqgv+IJoUdUFypu5sHh6xU2hgJni/Nuhhll0rsPbb5B9SXQ8stSh2DLlblUWgv4UtU/OBbvZ56
vNvgSW5s7hb4wyhY6DUTDG6+v6CYTMHVWhR85+wqzFmQh5khpPDgs8OTJXlAGp29WSutJucwrmfW
e5drCQk2jM3m/aQDmapUZr134zInLC5kTH4hrCE5+xsinlqYMECPiMQax7quRF7JXKyHxRTvZDPd
DkiN1dbztNqslpD5BTx9Dqd1dPNOM/d34HvLXFvwHONJN9z/NiSxu+ZIHK+qs8qNGSUPBrw7kiQj
fZnKSsVSTliG3FPVwgOsAtaV2O7WOFLvuc9slyx9P7J1fcvEUzYCHS05NXYHUzBws8g7RNT8iafJ
8JqnSr7J+VYzYZbDWDDgmH4ppGLHuSwJnA+i4phWf1Tw4hLbik7Z8HkbeYmYcLjGx/VTWIOhifgV
rQG5SbpcNGeTg+csgar5qBFNVvkEgMizdZLigAp+1Jp5CRKCnxKX1VwlQN/prwN+n7XoXvsO5Wz1
nEVQko6DniLix5P8vfwnd1eG6Ulr6qX8BevDgYaNkmNwQ996eIVMUxgJsi/RjbGXOTZa0Fobupsm
AHk+QjZf7MosgFp/WjHv3ilPSbVsrN20CIzaTwOTlk5Oy329JwUyNPiP1Szpj3pVT/4stZJogXhG
UBSuJu4eYZ+PWm5Lx9rscBRQYjRYWlnCXzxBAsO29sHD70u4+EijMDN0w4nS3FbhHhD+87ESda4t
kIVOfaQ1bovFJWBN3raLwUEkO2L+ZkA/RKzCgHY3xRYxA+IouNCwTKU8RvGtegr+unHyIJWXwkVp
nfIV/trV5e6KZrdOB9r/1TZtMVgoSH+q6X27uLJsRau/JS0/VrlZ5dKaqUFeOHFvyX2qWU02rSUF
88FLorIf8GXQRYDKFUKShZBAFqu2A8MVwFr5Y4wJ67gqSLwxW3je6hyvrdP2r9+Mc06JGmHfIURo
h/5bV5pQw/ZNHbXjm7fb9ZohZKGBnWFSw35vgxYTEkJUj6ZZAr9WsNaW1K5tj4d/0Fvq0OKcoXyv
MXyPd9vHeNFSM9V/+PXnVH9fWbjsDl67ymIvNMx4RG7ZcFJkWD8SAGsFnOyy/Vjk1LFd6GgtTY0I
zjLVu37XpNC/KePt3UMeGduCwpQwHmXUmL44FcpVmZeZK1R70XCctKCg57NKZOSvADkE+vScp5Jt
uGZ4oXs02fe0OnVKdV3RBYLwEwE4+2FGHFbfyDjLTtQ+rbkNKnEnTPi+G7U6ACoOYmiAPNbWAL2U
oy2zeYqPHdo6zgRfBO67ssuFhwgUaKF/Cy/hhlderCgLI0MX9+Qoww/ELESzzzIUDoy8N1EmPlVD
SCCUaJ37SZvjCduO4k7EwZEnUsGqklqXTVcHysWqn1NomFARP13HXhMvhhDeRMFwc5yC7/If7ZaY
GCXNHpel4wJHvI4SqYvuql0yp/ZtOJq7uLFx8v+6mz2xrk/LnB/AeRz9VjfVYOCBjV/PhKiwxSNM
i16j4jBQ7EUQg2OaU7Co2LLxkK1VLln/qb90u8TbSg76HtOz63QyNInRrGoEq9lpaGJ4fuFE2Be9
7PNx8ci0WXX8FJYuhqdYqS33gV9zvFM1G30tJRpQ5PsLrNX5SEpGIe2trIGYMx2EnNQgL3L2YIa4
69vVHItLHe65Jmykni3BIVIsMvUPm6i51C+mXhBd4FTxoRF8tHFECSVFEZQoVjiqANnCYX41Rh6t
yWsXXSqHqrve88uF37CVUT7qhqW/6PLNBXQcNn8kryX+YhqzYu81FWpGaEpbQwq3r48jVg2eCJfN
41rDKPsU4osvyNTMhswk2w02BSdQ0sGJdPwUOWL6NU0DMhxVITFKjj80cejeW4Loel1fUiXKNYtA
cTm5Yl+Zgjq2HNxdJoBh7Ovjp+WBZPog7cAPfZ5dnzAX/HpRM0yCNRiRLeOf+CaF3HNLHDjO3Y45
yJe4uSRWCmdMFWa+BaheQcJ/UiHEgTPhbVhoczd5nzQYy29sCxN856xZEUl5q8bVRkITLUgS0oo7
DM7ij1kXI43AsX4Nm+E7IW6uKzUs63wilpoCMg7deTG14hMJEeEzRE1AoTh9SpHvdAfD5RPZ8zfw
GkQMcunqhIGe3DmmeF9VAlbKOe39wo/kLnmvpCzC0RmB9bqlIFedOrxcIM8LZ5rYztl/rYxdSCZb
CjLSdnCHmU0h+9d4wOu9p7WQV8UwBabhhIDCPZVpHSv32YLUfvWGo0MFGXd5Puzq61W31lGONdCP
GkXUWEQDxxFyTZtM0v17Wzs9zRnkb9NCgSDj0omHtzy7uD3uUWaLZ07x7ui2SNrSLtE0QbAOZv1n
ZieIdv2jmCOuimpuYa6GZctjTA7xNen4YU9M7zwfOxTXLxUGUF5MRVtOU90sR8A4d9U+x9TGkRY7
TKbVp9Sx5sE53hjKWBccltzcBSNAv5mQuFDQFV+3DhKJ3Mp4nIXMjazZ+9E2IkGXOIsL862sXUG2
2DxTLpK1N8vVGfV3djSC+U+65tjiYfDMG8bmyZcmVGNVCTvvvVU29IRFgydj6h22pmBhY5yH0VZR
7O3tKPEm2QkqNZt55uNHjZIw1z7Q4218kIF57m+n7p3ve4UcWQ7eVuPFnA2usBk4ZOUT3JItR1Ul
Xfb1DJnv6MZb71ABvFWw4OzMn/kqgIzq6u0WQrUvI/IVC5TzgWx6ohgsvBsj5AIFQlWcLnfDE0Gc
9hIdSw/zSnWVlOAxBC1NFnMwW+Dn/rmmTfFc8dn9M1BJaP88eb07o2ykjWpk3gt0Z6jF8fRS3xDH
nX11wPVPM+7yvrpgqAmvhkJnO5vn4mqj009b0xvYq5VqU9DqS4qcDAubNige+yDjup5PnpMvEQ63
+sPbot3WXtqo+QJYjuSMoxkngcDYQwU8TfZQ/odPGCXdfKo//eGuxKR/MqRSE548Sh2UVFDRZdYz
sYTqdzA+Zi0RuVLr/c4RX56gHYcBvMhTcQX+xMz5s+bOqYyh5C3pQM+Q7JjDcDVK35TwXQ/4Bots
Xlusmp9HuvIj6A2UeUraOs3terOEDeqg46wm1KB1xNliR7pz2vf0zPkCi6FKHJHAxKWYnEEIaDA3
W7YWAO2EiHlVxsyzmWniwRKuZ5pFcE0l2c5yxKEEHqB/HJNtpaNWQtw9WyqW+IHaZVNqc7Pm6U/H
udIyMZgVOZ2zL1Q7JrSQ0atZtFs672KjJcX3itarbGBR/52HvEFyVRWQYL6x7TeIR9Jk0MH5r5Xw
KJZ4Y3xvp+oLjkJeFNzP0L6bB2V1yctm+U8iV7Jql/zeCcUlwZ1p8anBVuA+T/gfvKj5eNUlXjDq
WVIOwIBwt4RgrG1cT972hOECcx+n+FrXc7x7FwUfvI+xCmioo5HtpcqHmss5bMj9xZbnej4wjkEf
0WpZNfc9FQ97Pe9qlv759y/JO8v4UQn/JwquM6/cnZkJeJWPenhLujh+fKV5zrkMOlvzfcf2cbM4
Fc6WOwA0R2idmEkR5Tlpo4Xz84grkzdGvIm5k3A+mto/dLC3mPorUsH1EW0Gydc0CVG9FFFQV5bg
nCGbfNfpMEVvrXiFdZf6LK+zcM8Egiawzn99nWyR8lKNCnZjadC3m8NpjMu2vcen+FJeQBJzVNAo
hao+46kjZb0zNokuRNG8psRlagSdC+DwXp7mUhCn2yF0UMdc/WpsjOOk0W6y7qY9s28l2GRcm4AX
p0CCcIBec4+t29dnqt95gk2LiCi+8gO/sFH2Tdes7JhA1BJd43gxhI/Eu/WDGKtg4vRGy6YiZy+t
x5s6LbjGW6Uz9tWYLxlG0c47Tx1lfH6KwV/YZZNGJUMLAYswdh+Yd2FIfRlr6pHgvj6aHrO/NP79
wYKa+XgPXL5OpG9gl7gaU3T0pM1ql2uW+vANGbyQgUnKZCE0IL4RuBWlg8Tma1uSFmB6gBM0py0b
ewDKN98k23mOe+ddzQ9eWCinJQQMhyeUoTy2T9eGM4MeT3RK761AZxEXtdkUjg1AFdYd39Fr56jQ
0deBMjIs0qhCvJbWuQgi9qEA6DN6B2Ht71riXF3SbhMtMxE0CdoiH5h5iauJYqJGahZUVSNTtwnW
q6LNRSFOpXVnOqpz1pGd075Rzpc7VK5oPAWRQ4yQbdL3KMRq5xF5xltDq7wjRobyo594Bd0D13Fn
Ber+6g/euYu+Cxu7TTPIIaDVMZH+5VyT5+9Aj2lDPxc2kHkov8D0jjCYhifFF5TJWJfwCYDpI4Ad
aU1WxxLxEykS2o0tdSwbRLFXkWrxkcIwwaFv8am+u11H/z+cyPawF7TKiFQ8YAy9iqQo8rF0/DJU
b3ZAPSUH8P4Koot94BmquPc6mYTXIm3W/K9U+/Kncz3pFCw1LE8Z5Ue5h0ubsZBuJ4yRXv2bp8AM
b1ZEJO/9dejqsGBHcpVDyst2CovR1YUUPy1yZLqknPDf7OtHCU4GmHZyGarA8UJaNTGTjX3Ls4sW
0AuMaSkEDsb9Ev2paIDzEj9+wzuvawQP9TmhBABCg0HcLgFTxbUujQS+SekJ++5uBPWT4nnD1wv+
5C4lsXLb4V699nBTlOm2xYIJtN7LKcFRE28u9/hCLKdcGS8bo+jMT+0onmDOg9grAS81GgZFqsTi
zhjBLYF/+QRbWgB3gyF0YJerECfGrigmX5PFT8TYnU/95f9ZIp+z3o4LgVDoi3ARv+/a3lAOWamd
jr6OpAqRpmbhpO1H/WOi7wawEwWRFUY2S0mZMEfRKNH1EAwRLF9eydr4O0XEDxQA3tA4Htbp0X62
eBZLXUCY4yZBPL+7X4PixKkPHnyVhcJKogcvfEtmGtpjFHLw3z345DHkCCmZcYJLBkDm0ghOfSp0
15cGLCUy8lt5m2SlwZQfgs/H+WnmqvwkQd5bhpm1AFUznlNohKAOgFkaXxjkRYCraMZtlY3KMx8o
jSmpEv+qSM7K3Xvo9qENFwDV1lg8sT0C11r3UexEg+7ndtYMnjkrqoJqV+l35ALCvB1xOxktA1Ma
D7iRpI55tys0Lqr69JNx+/i4Vpu0QTPja9yNTGN3zDtzM4tTO6rY6GNW5M5IClSYv/wXlIhxbgMn
p32acWnNiTaYXgZp7AVHwkZgKrCrmRkzYuvBQ4zqV6wgc8q4y575GtJizq86lxfFHhg4cZcy8qdg
7XteQmscTDY9jO9DJmCrr8r5MsYu2kktjQDYjBxNQ01zL6xb8ACa1RPaQ4bIql56kaZlFzXKkO7o
1leXQvji3UR9YRi01LptqNSjabZnhW4mSa0viywhbcTFliq5EF2md+hlQBJXYYVbsFQe73bk02OH
s9MwpaoTF1+A1r7qaA6bjcUA3+s5HzG2X2vgBitgfrX3im4j9rR9YbgjpF9j8fqeES207qJjLpWz
+evOH1A68MdaPYxkgsU2787DLdl6R87o5FE81S3SaaMMzLH4x4UAk8k9PfAkfil1KAyum2C5CAGO
FJ+4ViiKHjvpq8d90fnTV56PHuC/oA8MjihWXBmjImyPxDLX45pfFfz8lA/EALD5ifGVXg85EPye
JuDQJs8YNmmBmz+PFA151ugSUJVOocTNusb5omhaUb2gFUSTvbW9IiuhddUbPdade4usoKFPpohN
sXJW2Q0+3Crt3+QZck+KSrwzCsRZDfJe3f9s5S7egIDMtD82LHf3gQYYLzBzmnjuirag/OLZ9DnC
bQ4T3G9JLSRtjosqG/mLkaK4iUEQv7UMQnTOxMhe+qp+bl0L4XjtxxF1/aLpExzfpLuGJh/5UyDw
BSbq2SIMn86Rgf7sxXZm4pW50d3whkS9Pa+WaUL+hqlDOhqA9axhhmxdfzdsWxij9T6JEw36j5jh
UlGprvJEgOzSQyrKnv1MrNuQX7neo/YApHOvxIPglfz01xK7ZlkhH2yjkkoomU217jXP4zKrsnLN
ofwksCLmBfYdjq7+RMapYLq01WYMiXYpk5SbT+qT+1k/tXg9cO05lU7T7EQBtZLY+i13VWgJ0xAk
jbEu7hj1hNeikEuU0JaB1ckZiA4MpuwlxwjeVkQKMp3ip4VaZSji8krGfTRGJyl9lSFs31Yifa+7
lxSe1EbKb9JqT1+MnHHRAr0bK84dzR6CfeIPER4Yp4BHVNIYJjKYitXiq0Ci6E5O+txgSTnRSTJT
+d96s5yYZU7XF0arfjsKbnVYdUtJSR13hUi1vVGmV9vOfKhS4cFKeltIiDzqJE5SO9YAkEr+UYxD
rkSV/tLvdVf99tWy2pY6PD3Y1zRPJopO2yZJG6S4xla7Kza2C8Zukfb13oIBHQDzz1A5sg4PRC+k
pIXtXg/3nbhKFqa9MR2M9qlY50julR+Fh0CRh4YecGXmqkqFJrhTgUwTnfspu6VQoZEOpcHxnHUR
Lvijo/E3pRQsSjDYdcWar9clROr63nm6pAtvlIuZRUJCnuqmRjrAOslCFZ8+BqsE5p99LdPtMKSy
vcWVHEx4XlVHia4kOpOT2RBfyg+BzwV5LwY4k7tvkFpxfaVSXhhs+9BpTbiABn9btlfnKWyLwsWx
aN0lW3JlXkXIzZT3EEXciAGCzwqWT3O1iNE0DQe4LVjS669idM4IK2BdoXe85Ot41l4k2Qx0wAL9
EM8StozB3r3C6LTKkDh6sCh8NiIvlWvZk2F0GVxEPesEyWnhf2Gwtvo7QivviyllSbhGx3Qs9IWQ
Bz83uTVOTf2YuxYJCsVcwUz7FgwQz3mirBxj0BqHHRuXy7gaDRqRdTxjPRcsgD27dD9TpWyY/A0A
yvJm/gWFO4QK2SRDvrPjn5KfuJFJR98XxWkGeVUhOzU3L4AInd64T/U81MWvCO5PIIa/3NFy0zEf
Hvpc+mAz2fOpdkGCGCd35NdbFU2dZeLxpSLJarXJQOSCHemdsGVIl2zqw3bFS3SV7ZL6IRKssBpW
dx5TWTDXA8/ZW7yrCW9FHbCOhoaB4ZyaLX5BXGEVsVA1iGPA2yWKpTpJ7gtqFzlmu/mt04fe5hTI
jg+5KggJ7/JnrSOFHVc8UdCeGKNX1reVLZ1m4F3DQnFFqT9HTKZDGeA9N0xVhPhxo0LcCWjDOtRf
s8CfkdyNpFnOizoEuq88go3N8G1SCzfor9NEMKgedqRCc/RzOKP8Q/nufgPfSrrDZ1CCXKATjyVA
ZsM+lwXtaMIeUeYVAULLL82gQD+mSRVKOzPdRUFlioPE56WfebtwKeb0UjnW5MRrDKcM5JANIF/i
IR6PVelWhBYSS9snNTtUdlc4/gE+qfSMLkLQP3hXnVxRiUzPpytDuXKXH/HXfvDxyLr7jpy0E5yV
Gn34PU2o5vZ3FY7QA80Y8fjGxTKGHrKOzyoz2f0PIf6HP6Xxkva0+TXsO2vAwsas0UaQzUIUC0cB
g4KrCUVnA5WAqW347nsYfMI90KK1Bmnnf9dobjOFWi+w+rxxqa3Gnv4KX2mZehPBh7TgHeoEOq3V
hiN3T0hoVamMq+DFt6ROEU8HeWZDEd31dn0CHgrUYPT1XRTxcB17YyI9sNuoRmn05CxmZtaTQvnM
XXnlkw3TQilc/30Awsn7ryYUVCvV768ep2c4wybXCWx5t/bwVmYZ71j6I/lZo5wYIDTDaSmXq7G3
tl6GYNH5pg7sXX0/b4joyWhv7w5qWMvKMUAJIUS0I0JjwKBTEmHfFLnz8F2sneh/kLVCun2MxWzP
No41+Bfk6Wj5uq/Ik9bCWFuHcLMTy2wMreY/FP1pUGLsuAcYDaVU/fKiToVrBQqIHg6XxngL7YTQ
OuPMkh2Vh1LHnAYut8m5m2HXfiPq6m7Mc/uQELQ/v1QAYLZsmfDHfBNXu+p8bGOAOUsCHjhms87d
2zT8rRZCQQiVIPpiHgpXzJpoA0XOWPZuG0B2UEaSf71JsLGoHzu3+nLCRGMVotPUCJ66try8iafL
0sG7INe45j8XpEGZgeH7tyB2nW79UC+Tgo6sDozEgjFtW5Pb2sbnei9xlbBN/ZYsHG2jkuj5eU+4
kMVlI7XDQlIXCAqqJ+DRW9JJEMMLLZH1CbyWAyafVGLLvk+5WeoCEHGzOWD1Q01dNmK2YFMsVlbT
xXzeTDOqC6FLnkwL0BwN1VkB79a8+lCJV+tiHwi0xc0vcjnay4JWCaRNvhHHoWPJzsrHknJOs0XM
+PCRTA+E74VT00n9rQQ7pMgDQLSO3siAVoUhqIYrctNqBKYSZqwjZtil9661aB3FR3YAJWlFGotg
k+Rut88pd84+oNKdSC9e0CCEKRtnXmgPwHMcxVYpECiaXElsrXmx2IAmtDmv04PqZJyyEABM7+3K
gdkGP5Z+nZPU/eds66Vu4sOGYrgYJ1jh0UnYpYZ8/Dw8/5vXC8z9RBYQsafC1XnAcjO4aMoZUmiw
4GZKvJbOAxnPDLOZ3G4M75Se2FijgR1VstnpnNCUvN6HvI1lgoUiFhOdr5kTZqL+jDw2jFEMtcbZ
sxnTQVCZx2yxU4VIS1P8Qr6UswP6yYxzmE95XUF/MAktISSKWukjYT7lutCpHaxrE7tTew8hhyCE
H7qzRm30Iz9l04HmsDZ5PUGCgl6EKC5yVDbwN2JOWXLVrrUY04fM9zMLfxMax78JXyUQOwbYq7t9
pZIHGKof8K2ehaEgJMUA5cR7214chEbg2Tu6SN7WP2W7InM6bbagWbE9bIHpErDte+Yn2jH1CtAw
GCaBOu0tRAiJdXk63dJmoE5VtzMKieejoqINhJ2MOIobqEROz+toShoEzczt/CsZo4zcblqdhCLS
nv240Qa4/cXlfNIkaqP/SnNQqgcpl0UDAisUGSqfDK+aUCm1/8FYXjG6m35AflhftBSn4kXQFqMo
hI7mPjbf18iZvnE5btvRNCDNhAKB6TSygCgjN948Tc9EMSz4gFpvbn88MrsW2DmOy95L301Jturv
Om62ZOrOsv58TVKyyCy3cNCrjlwOF0Zhph0Y7hU316V3dwp8OYWGarcITav4f0BEs7qOlgF6zIig
5nsx166EuwVp/iq2xADK8G1+uP4UEl2iTM8gZRVccNXOnv1T//cAUkSsxR08WKt/Hp8UFhQh/Us0
SHGlJAQ+o70jSFTHCG4XV3jBFRtP/AEISwBUBMJeneZa6siQhA3J0OIZso9lM8f+qZqgSuVRQ86z
uoUEshxZN74XZooIp2i98K0jkIlWTe+LAnExvBNyoncUIZnG/SqVmDiLGecRCkj9Hfjm4sK9UUDP
jTh9hcw9bRxCyHbvPfmxss8U52oTIb/srfEN0AvUzpgKx5HoRVNzK66j4qrVHNctcdY+rcI3ENbq
vxh8jFmuxwRrwlqxJqCapmZ2o6iFEH3Oi2y2Fr8HtpUeEYo8ayQ59ICfDH/9vPe80OaZb02RjG9J
KKaLO5EYja2m3bIT9JqC3b5cJCMozyJFDgoOr/pDhDWVCkSR5w1t0ZFCOPWG0jG5eYySmSJmG1hR
qDx1QRK+As+rVBXE9aC7izLaLr15XDl023IrRZEqKYFcEZnkEYVp4blMZcz8+Zb+MlixHKUVNs2O
yHcSeHdZKx22VtrHy12ggycyCZ4kMnSr+/zD465eUTQdxIMN+cvXSfvqrhsGCgJ9U4IW2nq1quAD
OdvHIVrMRsCOd0cGlFnmXPuggfVqc5jPGn/zD3Ru4v1dCfy3m7HP3xwIv2104y6IuA/FIpBIuO/W
19XSNMNJXm3UMDMRAcXqV0Ci3VB1B0IkAk6M6OzOfvUAPX0yRpWkhdSaIBShPO0MozaBmNm+1UWP
V4gCa2Q4MVdWuO8PvvKNxzzTU0uODiTQcNv8ubrT705f1/+I3DDqz0b6P5qInkkiLpFUHOCEGxUs
9jZU8Msuq54VdrcD1o1RKVZUURDeOY/dLpHo0Wt4VXy2FUhgCRCGvk6nNcjVly4FLzrWc0p2GqO1
8oI2c+QvOYiNzFurfHYUKZyUqiCOKT4nELp4yM/XFQM/pi+hRRgtPlRyWCv9uZK69K9d/2bkvu24
UHjTEQ+aEv+X7jiWxzLIR/Lt2O17eCxxHYov9QfaGdrftYNHYBblvpTEUyVkYI6Kl5n0cYXHm30c
NQoQ83+42Vu9DcD3fC1l7E21KZ1cN4L0NVNcec9Lg6ffch5m8GZJSoN8doQPo8Q8r9tLytfZlqXq
gdffu1AZjFSjXeQr/iktQSVl/+/5k82Ugf44qwI8uPFvFWjKOR4rQLARoUjIk4DhfOhOqkVJFwNq
JfOHa1tbDI8bIKzYZGAQpMnwxvYwz19IanWKh5v1ywbv8OsKI284nwZuhz+xAMqsPjuH4pXrbZlL
krgr60gawNvlcOGhL4fS5vWwCBUc7qvxonDn4cbsOJOmjWxO5JzB8R9CvyLN10vINbPS0+sTVC0K
zODCPxIKZQG6Mlp98Tls8PcZ6KsC66escdhpGqk5U/uud+c6iz/dDOINLf51suvTgB7WVG6GUpME
ptV8+SfNp3mlMb5UbIk/ZQ+9p99ruSdyTJGnaeBZrUkPPFtgzjiivXpJ7akUZ0WqUwhh6abmYAM9
KFsPCAeTzS41eokh25PEKQRp6lGs1f5Sm+I2ySUh+bHIAFE/ZX10UCYspx0mRJLQCoytCcH4gZmi
oOUxrj3mLVU/MIVJckpE3WpcRJ4Xcc4ueMRUkE9BkfDfp2RyGZfSLIAfD+JtmU6Woea+NFIWcDzh
IkzmARYdKGOVFZ6oR3F7dJTts0C7OtGWT4cYa9kdomW23LXYiATfnSHzduUq1WaARj7FGmAuIvGo
ljkb4a/0wpJZMUdWJYpfZebe9A3nKzINtDgKDh9YmVAkTWf7JRPVFZGy2wSH7TV+W4EyJbmko1mE
mE+u2ojdorETl/brQJ8YXLx8JNIW6jEPLHdCo3U1LgO8Kmu4wtO/LTcnCbL4ue3PjulTNieFjPum
9AiHfoqCRMChK+eEG8bQvut/QEziOp0ctM21DiETbBDtvOxTFrbci1hb8HcgS2tuqJQ+Rg71elX4
rYjwXHkcxVSycQZDknrLY7DzVsanrhI9iuesD2uRiak8ZndCLeekMnREkrPqrIG7UmjVmwBZsfz2
hIUsaigVj3T9Pjwdq5AX3HQVxX6VqXTmiHe6h+5etjM019txqEvo7l3wseLAtNNeAq65PGk/rzze
jW3pSioEZ5+OLyjgJYPWLEjsQjhhWVxmshvmwEr54K0YV6hKduyKPDcOjmz860iyJXjG50hhxF0z
yKaPfXJN9O0BJju0ty6ogObNmSd2KzUEqYxphgay19M6Er3zKjfGOZ1PC/hb3Cqb0XDYf6yHM7ce
RxsWRCQ116z4gJ8z5dbLbrPs6bJyJ4qPmXKI5xMyUwhFJGIkzP/u2SlHOof+fDF7+JTIe0SHeC7C
+vAN9o5g4KQzFNNuZ9W9Bw/sh1T45DbNGQZZ8eX6stEgFHHn9AA/3PP6oYFAO3bwyTudEIHc4rbV
56zVTOWr4WanKIXRmOrMWQo5usWhP5I0iCNB4xKhNBYf1jLyilOMkiky8OCU/TTl83L6bZ3wVvTa
YOmoBb6AlM0h/PFKYAuUZjOdB+XDTLhjWnKVSfe0sBSPZLj4P7tNSI1wZ7TMAdDxE2H15TCC2RPP
etLr6tn1onYoVfHkEmL/8wpgaBfgP6l+J7V0Z4b4qF4FiccxPY4P0aDskWlMo7puq+AUCtgruoZx
T8Ux56KNhWi3S2mOVRpSPyTPs90FwxbVxZSZrfkf7q6xiiEB4PeWL680NjZZkc3kqtNS1hscYfzy
FYR5p5493mwtmNTkOYGdU6jCYRivMqhiR9D+0I8mPBveLwoZGZp/eyXEByrVSXeXDCbhhho0EdiQ
9diKf60SCyopLoad18H7YAuclcO8QZ9wNoBw6KvApoJCAvD7nqMJKamZ39KaG9MsCw+1aAMtinTv
2nh8lpZad9SNvopXqZR+j4q+rdagGD4pMguVq2Hsi+6Rp/qXrtK07cx+da6I6VwQRLBrjrz9CCzw
DtVKolhdMnbQ/3lzgIqncWIHjy4gNb1vhaDLfr+GsCmSjKp4K+thl6P5siFWWc8rSYWUqdVIUL+3
8DBntMTUdIWZG2dOg5sRBp98y84t61smxAiP6l6xH+NJ3vqmhvDQoFKVIdsxtnBIagVnIivrlZfc
qGuLZ+Q2QmnXlm0vABM/JzxJuc4BcUQzk4b+nu4HAY0WsLdye1+fkhSbgQqiGQ5zs9oh6U1SoQkc
WW9tRD3I78j5bbRZTER9YkN3bajToq98ZGbfJzHaoN5lbQF79ayg8PKuDtHvP9ysU0vR4UmR1eay
rtudcBkMeolObi6eYkR58VE5aFQsKc01niykXaEaEAHZ8vwkjygcIlNaMXO1eH4l0gSIhGrRZpNa
fL/RjM5lEzCnLZY68paom+XnqgaqLnZb469dzTy/OmPmiefhH09TgviZko+uMKgWabtsSZ6OJtrh
XZg4OVC0Z3xsD+37kqG3hKJM5D81BAKiYBIw8I/PnaM80VABT+ky14xrtsPMHJvXWikNTZaAwihK
vJbvo39+Sgbo0nmRNgxwbLMt/Tplz5Yy7cAmmfbHgJeOhiaC6e6wfqe/wlihYVVNMXRBtLwmkxnx
cqSEzJ+Awzcps+CF21ffCPllRPVYDuXK2n0KmDq+EXz6Lp1kWXg7CCod2xfnFL1pIjKt31SXC3v0
N4vTnKNIU9+VXQRPGvMkTVLzlfMT9uVj5ZBPFQFFmEykCzyTohkVFbomFxT6FM7PfhHObKKEbdj4
lELtSxqHoBXuqX0LcPoY1c3DnILobMHcUCdYPOy44oClVwMuzTQ8YVQBHC5PWgPmUMFPqZesIXBQ
CMg7lQKvGS3D5TUnD0WOIImDo6KzGf8uxMW0x2jAWMD/AKorvFaMcFWFy5wVUmdAxzq70TY382ZE
7y85IKp9MiQLVAzW6t0kUi9HrmB3Qt7A4iodgqL4/RZ61yiBVviucIcMbz1NRaX+Sk1wfES5Iib7
+U1BZ4IwtAqpZHK+UNk26PcNcSCg8swkLNuQ7T9vSLtW1XXQZq1budYuJO3zKNO6u3CW6KnaJ1Da
WqzPnaMZGiIkL4RGrLHbvdKKc8yteIyBVTzukR2F6YZd1TG71fnbmJPAh1VOtTed2yRrRc51twDD
JQYVR8deVC8KY6uoPZagteS5WOYN+SfQiuMU4Bl1/2AYNzCTxrQM0n2HthFoa3W7MHQynzVTrdPg
x9hOJccNnzNUSd83gFzw8TBNG9Pv5l6SnvBvYngDDEt2bj675VkgVrrpw1ZyqTFN5O/Y1RWSaDfO
ZC+X60bmN1hvTVxf+23MPr7BtkGtAB58nThKG72VH3d+xS7OLu+93jSHs4XIkodb89Au0IwbsCxt
I7Y6MqDBY1qA3/KlAipEYaNsCXrve1F77x+UQNSrjXg1/FzgZasdSrj+HbCE1h4xhQbzXg57D3Qz
gF1BIS2MGymagU/pzam+2XqxwV5EvyXUYyGiDHQZV3tjbasWwJR3zrZfAYd34VghPXIG9iGrK8hT
BnfQde71OwP8SjWT6RJeepbDY3ssviyXNkwuWkI6hOmAh2xqYunjB1+rWeQkHsX3Gg/o9LIHGVja
tCNiwsLVbg8GJdHEV5337zdq9ciWoCXUiJWfvFbzIsQssh5MxlSq1SQiyWSMDQPHwmuZ0FkMH9jj
u58CzL4SoNjuGEUDbn8FgJnggw48ywk2kGSdvWPz1hL4dLtxpC4ppujPukqWl0RMxVofmqZcg0Ff
eHQpk8Ngub0l6TY50ACgbSdpSOmMgoGFnR1QcSHpyd8zcCOu0uPoGyoBb3pQSYu39S9XBJEuszlB
AMxJ2IRp7LUsX8ygPAnQRi0GrvGaZxL+nYeUAmurtIMn157nn+HSN9DLvt/c+OT13oXWL8HfQN4d
IPkEgLIl/7scbv+FQ4dsiNOqPlcNS7+DseiQYaZJSh3KVO+9qks3p8IOjYv+pkccqk0YUc4sYXQA
GUkax/vOLoie3m3DemMD7bCcXZosvnrldYro7KboOk+b59UzwzI/HeVm5AW9rXrSPsXqu2TCE/x7
SOBDIvDy2/LBMNbo5U35cho7kJyIwdFxoywKccvaCgi6gabYvtNYd5XygXGBRs55+EfBGk2wOzbM
pmM9BgxnWdvGe6UaOx+oEr9wbdKn/3frG/VFWoVq+DbnCAQ7ioXpbTESuK3+BFxqmnwa2axIkAmP
1E7pCLIX8PMkdUjpQBoPQEHyR1JTFA3ocr8uiea+OylcfF1FwKKX++xEQ5XM4n0xfz/1D78Tsyue
PpTWLkwtgdC+tX16Q3yj+EW61Y/B+wtMREMh+Aqrj4L1QWgM1lE8gg9SauNV5iYEfLy8FS58wh6l
CaBHJgtUN9fCYumAwN8GIu5RKC+baCSA9y2m/njeuXHsghzEWIA9YcRONxK2705VbPazuJaIfzsF
RNjR23Z4pIyGacFQy7kzP5pdp8CdhW7Lc9eVSJ47bPj9TQ4OribiLiPsgH1SGoDToNWFrenbfYCN
Ig0cW6hZOhHvdxe3BE8wFqStWdgN06wPTaAkKGKeFla9lz1z+NZ1YRzvisTXm3C5PN7i02XoMSmC
LnENhMkR7iaKrz7Ftms/ez/bPS91JTzWowQO3DRdpVm9pAJkY/ljiwaQwrhJd1Ht3YblCq18PTLl
JmYvDQgbL+4EmybSyebDfesGJ3OdIrMV5LgGnVkZw2yNjmVTiOKNNKSoemWMmY0df9+2GWs+GZCB
YxCawqxrBKbQP+kVlwwDtj22w+wObf3BwTOeIumRQijBaG22KpOYGuXhvLzlSlQFG+VAmaNxAcH3
qcvsJ52k3O3hQ29c/mRWZ3WF8ZisVxTlj603Ts/r12DvMGlJtmJxIBSW84QZWN0wDgQHMZx5ot6H
6OQcUWsuJVIB1MN0hiJDwXTJCSIdg+sw7i8ytPdRLAZHiCyR46vOn/8B4k20mDQEDWWMg5uNzbdq
iVVE4jH+DrIZzW2J58gTc7nzXMRJAHeQxjlneHdz/jZU8JURdJlOJOheBl4wSLpSI0C5c9jvq8p/
iq0GV06aTUTW+pGZEifJdHU61fsl+iOtlM+sIcn16rrXxFz78ASKXuuSvcLkO9KXc7cn423ONwMA
AvIxsvG+9qqyn9WYKEnrwuMAYhnsGQcQ5uO76bIy7rPW7hxx80QpeNFYCxEV92XBoaByd6w1CXfF
xKfaZrM3q5mXGu0z5LMdXVVY3bjgz4DoAQhY4IvU+inElcrnw3MsiXsjcof7OjO+R5i1Mq0mu8nj
ZKk2wmMeblb7POHuYyhTfJGQ9vcOQulnLM0uc8z/ayYsM4of1tOnmtUBq4Dw6Qd/8gww9TbDObi1
3zqv8zYb41c0Paaco/s8y9hJeAPTYPaU0tCPBIBMOCgzms8jdZDMqppHO6WoJspe66FzB+JJzya+
B1UEVu6FubBX701YR6QqHStI4yN7Qo3ZMMO4Sxc26hTRgg+aB5TwLsuaDgRjv1domoCJWsrJ8tQ0
FEzhErXggmdMpZnMQJsZfsf2HTHUDxOFQs4Aeb2lKGR6JPoNgYh5QSEpPYz6kUTcHnxCywSMmsq6
BArPIo45rqNhs4EZhThNixuSvtpzfr+OVxUky7GfhmpgUdSDkUNG9S/rzAhHZpBwS7uVllBXSQh6
bzqPNXOVZkqoLK5NNx/bjnc8H+h65MKjlhJ3LSqF/YarXpHuQ/vq1j2COk2qDBgIL4PjPJaOfDPx
A+/3qocig7+UemfMX8xcH1cq/78IFSH78wVRitCDkX7D5V/XqRnpuIFMaaW2T6sqyIBtffBhTslC
7XotPn/htPalrWsR0ek818+fkAr+VrdKZARz0e6WkUIZhPNDV26DGRElPZ/QrggoSNqQJTqcWDCv
Fj3TvnUS4rJXlhQlqusHeL49oyL5DZZdyAinQQroKr56EbZG7S7r99pTieQZBDHODbGQ7fdOpbCw
E3GwKAgZ2pDTUYxtECKkIuvZ2+IQZs2+b+DYUhKp4quMmRLVD96CKm9Q71OjZR/GTYuNKQCvIREB
TX/0rCSk//oBrkO3lIKzt1zyxh6BCqAIK+72zkYbd6q49z5ua64byYDwZT8RPTu/JX3tAPDzG2NX
RkvkzLhKQi34dCo7kGlteKyHByqlaVfqZU73odrLxbm25v/1g5l+DlkV0FjYpKhU/M9slbBRRX2d
fLMhovNcdTNLuMj3zkSkj0nXOQTD4xiEQ5y7OSFvNywGRgcy3XGn5TrqRCk1ZbH8bLerBypqmAiP
GkgqSesiGiUJEZBn5EFfqF/cuQ/bNm1dEltbzzwWvQ08PUOfZovWKHujKzTdQCbsdLzCHQmsc+9t
WN/KZGFx6bCR0xEDL0xY0s2Rrss9Qa+fMrBDHxPTj7zmdm5WOZB6KWzYPjVbguMjYgv+EX9hNXYN
7TjtuFjRCVOSUqzJAygNNNBXZLE3EobikKJlX7anGT06uKTlQfLuxGuwNf8tUFQ5b/FnSUPjehom
fS7MfrlJYHLWjq/D9c0jp5OxhQMSbl8jlCrscQYVw5BLnyne+UTHlQAA+wvnyIdPYWdWEUfbLXQW
0YrR1gzJtPQq2ZJ/jnLYzaqabV+9qdsFth2cPwQKDt4+RUCpRHr/pB2SQAeYaFV+HoxdQpVCeeLn
gmOnCkC3ICm6iTzlMCrc3t/xWytj7SituqZffqRqeimVGyRHCZignl3hxd/2sscojeRqXHyjKtf7
QhfQ5WUVKg+Xu0Hec1pp1TFGdEzwqOSczEV2nUVt5bqSc074gR7srQVJVwSfw3+8S6gdcchf0XtI
lQGvFsXjCLSIyEw1UKs3lt7be8R2vtPkMPY2npkOdkCMKLY+9tRLzubFyr22P6pAr0fhSZIk6QgA
ZakzzEoyM55qxox7gMhzBXAp4fYJKe1iRaCG9OfovKO+T3J7k1Z350erEIdJouF65pRJKGQnr/uq
jlJSZxuCo+QmWDaxaomH5NHxm4ePVogsZY18G3E1J/csLT8hwA8vBJx9cRCvklz/VbHlbAlGNBsP
NjPZ7YH7ydXfJkEmzeoKfn71W+t7oGPTUJCtCwS7Z2Qa75eQqU4F/2CEnLPX7vqbXavEZQmxF/1d
FDN4ZmON/DuBMjw+t1p2YtCgik6vrdLOkJQc0HKXTyTjC6ncSA0j+THhyESNN95CFs4/8Uyk9n2L
qPvZ6GBhq8Wz8DRVgDqVf7b9J9oCMHJSPEsZ4J2VmWk+HGG8PP6jMdEdvpVeZR2ic4qRcJgPdv+5
7oZPVNcWDU0HpInpjg5kXXOoUNnPFaIID4upWpbN4nk9uHioT7Ha9icEYvn05GsOSkf7SgmoWGYs
Sm2rV+uekUAuacJ3NYEy9zjavJcuwiLt/3B520LyW/za2KHmqX4Sxzf4wpZcHu1frSdA/NK4JDSx
yrYK14G6YjFn2qLhkkXlijtaGx+ncS3kv0qXjVvONwalb1BlFYlVybbui/W8K8INkXpi0ePlCTU8
1dORm1hMnAT1Pm4DEW87Ypeinr/S4VViyQBkmnt3SD8pBg+/WLKlzh3l206Aen+y2Ezy917SVCqZ
b4+GRxvAFVTvzlhIYL8VdM8V4zKLemOErXA3OhExuy7s83snybE2GJd47UjmG0iFRErbo7Jq2P3m
w2p6HThpc3tjWUsHTZIVp8gcAa6BKNr75AEp4yJSowA48OAOqXqEjMxd+PNjOYuWxl87aH8AXE+Z
SV+nIMuU/Bwj12JT9RzkdAJy8gD4hKqElk3dDl5beIACrHRCfdIJ6XfZaEeaGQqi8CAyqA1jcRgZ
kzSmdP0efX0N66VX4uTYVralgzUyWm1hsq2D/QppmSGaQe65/VJLB4/VuppVo+IfrEVt+VRhIx03
p7Hfb0p0d3eJn0kyBxZe21EVmn/kF7Fm7hm1fPhUvYnVG8H8Kes1LDUrciH35lFXKbSSQUVizy6j
Km6uc12nREmOXgrqYwJnrtiYvxknXHoYgu61JlS1KL+4J6hGXBynMH4V94sK7tTJcciaSCUxmTP7
X2IO4rJRtWmdL26TXnp8OiQeWsztaLItUB9G85NaN7+M1TmYIxurDqs+gbauZXZEWaIPqfLQCZG7
H+ztWRg3Aev1TeXVF8SItOCdZCMk1Igoflnn0PUnB8xxEGeUtQ/as6wYmTN2xZqoNRAI0yTPCeT1
0WRHz/CNmFo/6OJe+37JJO6UOWCwj58t8nIJY2Kt4UHY676tikgCze9YxWVVegMpIlGmR/LFrxdo
72bv+QXoV449+8JKgW2u795J5PqnSlr1GEnWzjkJt8nE96+BM4nyCSWvPw+i7MWDzJkZmxM/VNLl
ZcCPYePivyoru5Oiuh7rLguH5z+3jKngWbCwhul4Lz+xqWqB6pbdzp18LaMlqwg4uUlesnBTbnd2
adFb1XBJ9AVb0eSJlYIU2/trhK0Z00cjxcIYKSP0uafNS/GuMbRmvwgbeokhxBbJgG2qiVU7pFS6
HEQ3ecEZAywgawfMAdDbijg56DU73cVow+UQMnO3r95B5eILZaGLC7e8MYiPzemrNAGVwVN3YfgH
HpSMBJUX4RXj7f5VHmIlpu55nXl+uGMYVrPdktYTuO7m0ZlZap6ED9N0+yPTymgMkf3I9pXVEJeN
HVzitklowGgLmdEl2WQ+A1vNVYvC3zvdNcRuxKAxcn1OQlI8qpzI7A/xlWwIjd9qBAxbOhPyndKv
wJd4+3rN+jn8kjexp27s9j9WTrZ/PsqQv5PWna6WxnXN3yykHJh7rfuWtABunaqtorFrI5UUOnXh
JBBLtlG1pgt4EcVY/oLobAThxeB/W3whUreYAK9hcDbKeRSDqaI/JDjfzEGhDjJnl4tbCAvr3dfZ
xxnI1kQam1QKg+IqNNutGUt1fgNDdASNHEWFTADkp5SFKQpFlLO1FOgRBaCy1CeLfJ8P1BjV9b4Z
kPQZdJGrFI5r06rB/7KxvVAnugGn61+7omDYzgKES3Kw98dTbo/jvNOZwHerLrf3LrACRBW6DuhQ
pbVbms6XNbb6IcvqEq3X1qfAlN6OHCgPlG7tnGqzcY8sU9kSOrj5RpeBlMXWm9jDOIO/osUh0iAJ
84BOGxYo/8mYCe6/k8l3RCokP3eXoKT5nEt13V2dCpG+xCoxIgDB5OFY6Z9tOCRDaBJPFciAULhe
st3Vabzcxa1Xap3QoAccJ2VqomW61m6EvMxhh8rKYVuYhWoiZ9DqEdaqXcdz4XD9fY4bBbu7p1My
2BP/XEBIOhAcTrQJgff6vCgY9IQxXe4DF+RqjnqLnNV7MDYlo3HRPuet8QoUa5OgVoAlMN9o+kOw
qKowM4qHOF+WUUtfgrv1V7ydEXGVgTHUcj0BAY9MW+vQP1gVsU2vf9cEZZ+CIOwpnKngg8NUvedv
pNWj3GarQvskeroxD+KlOMZVK651mdT/kQEnPk7GH6Ud/xG5wmyDhq91VIRGtd2YulveuQW5Ev5r
4yHkqyQzFSGujTyDaaPZWzrYx7TwbaU7/cWEuZeIngm8nZ3hnGy4bK2eVQb1MadeE0prZFQHaPoy
+dpxV/iyRZ/DQEgFd0lI1It1wpdFqBhQRnECEvMsd0R7lWGazP6uOAu4Z2zsM+lxzjQYNTz9ZOTM
AjAW5GsdsTg6jCUP0mDetyPFRilUQFl3yIcFo2PWCVnmnB6mcVGmbHdyIUJ1OFa956/qiAtgFULg
bqFA5E1bkOeF0AgSv47zRrQ7y3oP/OaroLOuOtLtsY/8lW/Kt76b0puGwrFOjO07ZVkWlwyiQC6l
4gVSCBEmz/NzPTkUHofq0fOesrGI8gQ7wXHLGVEa0uTQmDZdrGrhnF164rSpq9IkBmkjnOarbLxk
DsHSE3dmz4Mkr3OSIlpffo28zWyUZEMLSQ97j/mW5yYngWy+w1dIcPp+T1iXPFuQ7YHYI7u0PQWd
RchUqsrsSdiFWT3A3IOnruGtmIkTpa8kuh01fXprQktT7m53q/StRNrJmaRQnQ24wtyiQ8OasjAd
vtPHFk8189bIzbwROABqhWjA4bvyLuEGaw+b9OAHmu4KP1UFoRwkf233WYfqJHufAGeseGHVKXZW
IG0kw8LZnv3hjKabsDBqmZedb4T43xr6I7PX39Ma1sukChYnzPQxh+5LQfO5kIqytxl4/Vt4KLua
g7n+JJU8Gf1jr8Ig7iAcjbcrydOkIg+ys5N+Q4EE1p+gqNYKMqleygQDzuYDPJYGoTTNY6na3aab
/4KYW1KQKMgIgxX0zCi1lbAv8eD67iJKgPdQo18YeRg/j+NmwDVVTEdtE2bDe1uQ21cmXQ/ZK69K
fnBsyz7m7Ibg68zesTaYGDMZ5I8BZVlTDxdyVn1p/ltdD2gqZVB1UeFVAEnB+mCbHuPebz0VxdGp
V6lAF/rLr/01DiZGCInaQ12N11ZolFAyjS39tbveK/CeX+dVDT+kdJO9S2nmBtMQgH1OIQezl07A
bOow/lTSSL2S5yp1GebLkPIOZh3Gq8+tn3TLs9/105JazE//XdTvXVmRkgSfc05TNDkNkni91xNw
LH8hkbrIIx2gandMPzSBMZVL27d7t4XuXdrs/AdNo+Mnqs2dFXx/+Aiu1+HmNmVZ5vmjDKhUYTeJ
UJk615h+oDjdOQuOKj98JKnD3vKhU4QMkAhJXviY3fLTwjPlqTfy4KzO3YDi1sb1sdLa5uekH8y6
6J1jChGu3m4KGXvEDQvDZZYpE1sGLfUFmlF5slbSaESpf3GZzJBwdANz8mxaxvTS2lL81sXHMsQ/
HH5t/9eqhW7OHu2mR6L7MIJp8fEkPGcWUVc1V4VafK+ZDwRHMe2ZpVlgpYBFApnh7ZJChCSpChN9
RBT1/j5Fl9vqdPCZytLb5HRT4L1SLij+KngvdY/Rmn72U5S1kuA+jOMgLV0XB7BIQPmWS/BXmAPf
9jQr7LnaTC0qS4Af2f56gX1VfGk11s+5kbtOvLtiX9Br3HKJCNtSgPvaDm0IeGsUkBDFIP9sIXlh
iuekFrTUJw37yf95DmmmKbRXGbStsTd/8qsOIs0vJb+r48LOY5xEXyiYMPB9/okpahF/IY+oP/Zw
86YNLLqtrhtcNN9RmzmVP5quYVrzWRIdAeVYkEdqOg+GSnXhrZX/aTwxN3iqQjrD8IyxbqJtVMfe
78hTE/TvDtnSu4p9f94T1T2fwPCwXmY83TeWaasLo8C14EUJpIjdSU1ZaKqGOMYC8/rP+7+7sb9H
dn3a7NQyMhertAffM3cliS1Vc9SSMwydZgytGqScEKL0Vl49iR8N7dFUZ1ayrDrvge/klPkqMHAS
gckBpRKx52ddv+Vk+ZZEvc3+KTVUfGigy+Eaxh3s09EFyfAuEseS1rN1VZHy78+I8g9Epq2Jq6iI
2TKaxIx7Z2kDLxu0pchYi/OaEeIjAsG5CmBZbLiLwRUQSfYmy484tVWm6ekwnm83OGxTIvprKHLM
w3UJbKrH+cEInRxoGqLvQr16nHu5K/HMAGnWdIHd3R6ya6VQBwfNtBqr31l2M3ymbDEJZNdPLKJJ
bbJqHLuPEzS9O8NsNNMh7NVCTKgW5sadHh0JMsOc9kGi4S9MsjSWvvConbC4XFgLyGDCDqbVvWMW
tT+M5gf0ITbZbFsk0dXw0zXmP+NXf/519Fn5MvUK42WR8NqJXj8Xhd/xvAVKpek0a/v/GrUlJ386
5GBeQhmO984Gj0BebE3B2p24BbGI0iLeQPk6kZhpDxVsNNtDq0kGGdEhwVvOapZA4RfJPnuoGRsP
NfXAofez5M4mNrtWZtbNx4qeYBvnbKbQGguLL6iTi1CZ20eXpQX0vGW5zqFKkPPKD37/jN/weD4r
A24rdxbPFaaQuhpIz3crXhpT+HEr1qiCfbcc3YM6uvEVgU6EeiXdQk/I97Ha2/4yZW3IuhDA289S
iwLE+a21AqNPmYGdD9VdyetWr/bReH2ATHzLZCzz+UyYMNtvcSAjyhlQOEbJ6OcmhYSjgRHbtVQC
8KWAkukvSNR7K9I+xlKDrzbZF/QtGWmh+pBq9USjiZs/pzQSzKSeeEPBpDZJumCcDLMsx9TM+4H2
jI4MAgwbwO+2Kzh7fsPzQ2KE2hrMPX2RbBWEg/6Usvj6D0CKTk2UmYM4wq1CbkIQuyD+ofa0nGi1
EKDmuAti6WOF2orMTKC7NAZyTGbzDwBAplZDl/1muaj4tN+S0umuFLCkFPy2EBVJmfaTLeaOaViV
3st9yV4FV2vdhNJSasAu/eiwSmVpMvcEVzuwGPTyxlrxuZFIRpHyYSnya8gczmYdh9j/e4oISkjk
QW4kXNRIyeKVk8na/ToCrtnL+oJP6p+SU1DMHlgLF3LyFgEquDYV1SHQp0h62pwu+4YzGWdVwNB0
19mpHU1lGsDXXT2Rq1tATy4IjaD90U/Bl54ow1Cx2gFGEZ7lGIV69fldZEhpd60FvV3ZL6Hxip5P
VcjNWoY5tyTc7OIbu4mFqd0erA4axc9l0ohcHarmHPqxP658sdROEu2NGLgN4mkF6PU95PXAM/dL
hPxHn7avXI43eyCGM/yPsedOtxfLYBkmeXIrCS9pAONr/qPe//avlrmP8p8ue66PwJO3IA84E4z9
BeM5QNd/Rg0qOTxI+nGankoJ8z/b9GDrYy76cK+igJkWEqNebPmsGoyFNBDrdUFHIskjbi1iCwvE
Wf7B03ymOYdM8PJz3OYyP+nMgmoB1DXRsyEjqTD80EcWJ7hCBQVDQiUOU9x7ZJsZD+UBl6bzmSSU
TOBx4EzZ5URdELOMl5NRf7O4NdxIoxOOeTR0ezB7Lhsr9cc+I07OTsD2KbCEhu14b1ixUs9qyjwH
iNlu0xDFuXE0jnEvCywOhyOcbFyBopqJLmYPklfNOg1xyLcUHtYjej0bdMoXly+KEQgL6s8R7laX
R6O51Ozdrx++Lp8Ens+IeVk0aG4T3lXQ4FsxIYmFZ/WbXJvsy0hqEAp2iVLrm4fePIqhKlgfQJHf
tMEEomvAJr/uvQHuOZTP11DwNwJigp3QyggW7nfrizZPjkxdKRXw6qjO4SYJBbJar3a/rdrb3KHa
BMQE/HKkhy3u98MxcD0HKk0eMnrqy6QDJJVBi5Pn4c6grf0hakjURAbjdVSLgMdXtw+LnJpkjJUQ
rhyLzjgCCnyDR/7YtXF7cqjIV/A/gPNukeLljBiQzq8CcJ6taI12MUF6bVSsXXWJ1YU7tMW37Ipf
LXoyxYq8mdDZD+cKbB50aAtGkOALYgMQQfAqq3X4yAMbKsHjjNQeHgMC8SvscfHyT6rNxWzipwdR
f21HOgzBrwSeWXfEmUYVxSUBVmIkNxPOIaIc56AKb55ls/Z6DNQOnT1rH+u09BA4boFiZxVIhLdD
0Jt4imlIjysKxen0gnOWBKY9RZVTcDq2cKlUm3MIEV5ZwZ2WSSM7Qjtwp9EL6ZDTugbL0nWWy/6m
Sr2h07C6MPY8UbLPcWYUdxQfLjHJQMjxvzydTCzFG4GVSMRBRSSYbRto0X6WjPA2odIcfPTDwwDl
2q+xt3chPfo0dRsWmGWX1uNaqHPYAaoLQtuXTl2C8Gwd7sg5k685Gww4LWVsLTQ5vYfpfj91ZYXB
e2IuW0wbrc8odC5HqDR6EruELxYcZasPFYpRO9xBJedmZFnZ31GZ9RU4qd8Q/5xlFBs5mlpFGUWJ
kxOhU3kis4RT7qnnVe9K6/jQBn0jQmRgtimTYcABc9WIapdP2i53j54aj4YOgaj0Le1AvOff8Kn5
WyNGEFB5nGwQsaKHNUjGPRU9cxPtd68pLdEbB6lnl4g6XU7+Im8IVqQm1UDSUOstVpHwrkEIdqJp
0zEeMA7/EgPX5zN01l2T1uvu0ERYryaUCBdGQ+ZefaOXVdsh5UHdE5eLzqDu+o9zd1STIwd7CQUa
y9GbunSdq1gDJ4cwSGMPTR7m1O4dtGQ1gU6MM5gCGZN5o37xGinYrHkUiAjFtmv4ZVdpKnoUs7Hy
WwPjhRSxtWV/+RTMIgh+a4XFC7DUsLixlpVRa/oJLaDcv7iLjqzQUr87aw5VSVbSvUebM+SPxqWN
NMpD+iw60FutTAdlPuSo1TRGqedYEAdWuINBuNnMoZoepD241oxu/s3+0f3k/0x7ZDlAsE8ixar0
XkiMl8S+RhtLaHxIJ/4ra+bnfjjTUw2ZguzPIvGZmazvJEpP4WkZxPh+lpZloB1LEHTC3O73RY/S
dfQ35huGj2zMfzvi0fLITUdAcF0UGj3/6oiEq4gyf6+KZinK1nEKiOuwRWaK5GpqYvjrgeP0ZfhY
IrUuT7I6+3M8mMUQYdKcFeUVc40kHyi+fg34uXMYXjfBfmPYXvOZbhPNbQb1Hgd9SBX4M4cqpItU
8vtufakv15u+a5jTLahJOjPovRc2OhdZ6++6Cy7r8kqOwAsEzUcpK8FdVnsB/6d5Fv/Ys3emNcmx
K3CleDOSiIilJ+4O46UakfCUADXrt2q2+GqOAusil26MymCILDjSLfr/D5tD9KQod2PmKAyrKUz9
JGKDpmLiuy3qtJj3KHFlclDJ0v+KKLPimJuzgTGz4R00DZjE7b5jAALChReqvqKiQ+K+kUac5rf4
EPNnnScesJZq9iZQFD654LSDjgcNcwYpMuTmxqFr5MsJpnGErWwyoByzRTehA8jqQpA8spxb3j1i
PRDZMs+A/CJa3TR7n0WDPYJsTy7ZKPspKwxJ6Uq3l6BBKmEUWuwa6pBxhdlPuVJHjMUbUlTWITjn
Gpbp6zGs1ORh3kRhc9DEhSFGeJGiA7rzBmr4jvqLmNNuo6NsGwn/18cfgTTd6cswl9zMLJPwTkOw
XnW+VpEtbgb8XCFrQfls9KBVh/KA13T+bDBUTHknR6CB9x9TzMToGcc5TP+y9DA17gPGVwsKvcdq
y/K3bWR0ZcwZSO03HMwbt3wH6/EbEz3X5aZLmgCcOATKQ4g3v4S/KYvIkMnqaz5y1XSVP3pBreWd
U7KRai263s/+o7lhYZ6kQbdt4m9vjb8Ey1W5G3kHoF9d7HN6xXECPmbW2S0Yx6ZF5x4aOuVEfq6v
8iehYPyhkwRE/l/vnodusSORx5peL+JphOszps+6C9FdH5bXa7jJCUy7k8K1u5YZyZN5pJ3J13Ej
bgTlQtykCcES58WdwLj0tgR/OMlISL2BQwaoAYrUjYKxMM1ruFfuw98uZhUGir76LDREDJITFywH
F92vE7x/NZm7fGuPgu3aj8OR6Ln93v70r0qKo9g0it3g1t1tIHbTt43GAz+Zmv8RagUNlAj0T+zF
RND5rbqPkf4S5YvzLRG98BRFAYXCSQ5VelIzPt84zLBpahf+ywS8JQEENH3Ivk3bpeIeS39lyRdI
/SB2nuo+vgwiBERnYMG37Apcy6JrvunDZ+1UYr3NETdLVHGM/vas01/B/K3kazp+WAjqsHleExV4
9WPo2t2Okjg9cbvyu4wkpD4qnndug3QMKRAqhhcBh4dH1CCXH81fsNtQoQZeCmh9RpbWdqzDCKSU
uBGQTJo3a8IuN9A9PjCVrDrpaltVzzcy0CL9u3M95BbQzAFXQlLh+ZxySKi26CHcOVZ4Oyrd7nnP
UVmqPDjfyrw3CjcWAed0JFXFSQB72VIdBRnVZl5L8B3+YA80UE+fd08UEvwMKarJU18yHqJuSzsT
1hdpJUjWctUx0mNQmUjlaPHyR/ZooZdx6JH0RU306BhurNkF8JnTjFR3UbRcvYnHlPsZv14ErgVO
umM5MoLOyxLi6FaFZIsKPVG+8M/fZjPNdb/jmnObDXqt6Vz9dfVGA5EiPjzItcwPN9hwHOOxpsc+
tN/vh1/z482boII0ERfwEYGq49ZVpzuy0uAYG4rlHnxYPmtWt8DMJVdGerYpgGmgV+94r8lROMIJ
8mBX1bwGUrbV6Ol/7QQDa+5jbIG9N1weRn1ik3ZP4T+AgSEcMLuB8RX6/PATTITX2rAG/56rltLo
jlcmzQTH0whMBG/WUBIIMKjrCZ5BPKfjQlNkP6zSS+1Hxw34HP8D57HIYf/jq2R9445tyBPYFaMS
POOJOUE7LR2dWHdfkskcPR+m78HYKUYWFqc++Fw1AFO8gtJLH/XO62BVpxxRwvIcn/REdebT8iG7
/ZknlCiy4X+5KvmQw403G97RrXIAh8+KBqEtu5pT7b5WNL1hyq396xB2wvUKKUxvhzc1oE8vXtn5
BQ7ddXRsvBY3FLo+r3XRVkuvUiTMKNtNqIfKrqPQlalEHPHq6PvYu15PsMcWyYyrd0GVtV2s/UGa
1CKLJknE2GgAvjCqcPahVTqeFBEQ0PBd0m0tzJyNKb6nLOgaB3Qh3x+reyJFri5a28uBsN8sgCnR
NBxA/CmA1yBJUeTtj0jgVz5PRz0JTv5q9l9do0MuW4ValoemWi8xAduihmESnPfthQCjgFxzTUMb
4ecRAWUhikrJqPv6bLyifWIozk9UdO4Z64uOlc2ttm46+AZr7VSnCD0JHQc/zxWMHtg/xs2j9wKP
nD4vNz10rjfosib+WVUtdaKpB3rkZsX2pF9OAkcZfY3bgRjFFZplHH/9UByB45IcvKbbeD+EFeQo
2Mz40CnsOQ02/J5DTD3mTmZaqWBWwH/QO011CjFiYq3ctdufDW7LebWmcF4o3KJT01WeaCR8geFF
OkDL2FsDwM/UD/ksUcDA+5xY1cKQdUHlL8B0Rr45xkGzGWs2NS1pHDuJ2h9PGhpReCml8vInQPux
vBOa7UVmzI1VIUweXoQlCll1OABqOx6sKPfbOfaHTgc0CpGWm2nMnv/779kQGsmRG0BhQ60mhLn/
wbhmYi94llO2shAlQ5fxQ+YazjHQWnft/t1Fgl2lCwWynIeKWqKPt61+L9Mki5QwWnXgbhGMSHGt
cy+X9O4bR8ZIAWST0bQJUjhcXNZWYAhfEPI7XJsnii+4SvBqWZy+qZqAXyDduIwHJvKlUjyw03ee
7vVgPaz0T7tvckrf4XrSEayzWmuQlqR/zBhd39adzCl4z12ypibjFCbH0/KNxmenZpBoZHy9LKWe
iVO0wMu7zSLZBqynczFeSB0w8QRswOvZRIm4jNvdzgHLZVRwot2oVynXxxenYGGpS7xtVi/4/zyI
m5NsaX2jM8Z8MlTu9uY7eLsae1kXdc12XSObInRWCZsvZjX+JIWCJ4AwnvYMSVvhMIqWXVkdHDF0
53jfuJu+kdpBeLM0Lw8V/Kz0/Y8+TzlV7afF7WrCcgQkdvxrUFAhaxNVTOd7HJcVWqHoS9B5ZH/P
Jj+ghTJBoTLLuoiWMxvaswFRUX8YW2zwi2+ILCQuX9IaCxdqOljYWpQUMJPCbPh5rORiYqBg5/QP
FtO11DXyzfSWV5LLX5J0pgbhw0TR3LRb9zr5+gsdXmZs2I/YmvUr/9QESWdrxM4UG70JQ++XWJFG
8tR4t4U2T7v8krCdqousl1nHi3vc42f4BwWa/88IH21g+MqoNfVUz9GgCwZKxmsVIK8fy5ApLmBS
L1hmyYrASfmYvO6izaGnF92z5pYIKO03aAjG3mfpVTd8TaCcfeDU6havHya3mV1nn0UQcqRLXlkV
uiMxQt1sYnWKuYUHiPKgmMUI6wBfsfATcpo007LdLmRs6gjvWV/7mt0nCg5T1UaABKPxxK4yzvm0
HJ9Fg+mu/EEodmEkT/PhtGohp7BzUpp7/2KCOwRo4kth+eIlr8xkBlfwlODAMLlqOiVudPRIga75
W7PLFMI6pTfht61a1OH6wEF7ZXa3IuDosoUutiT4Vj0223SS41nky+JCFwJsZPmn+8LPN/PpWMi3
vG5qr3K/beMDLErsmJMqTbAbNrWm42CdVIPWTmL2PqIiFUyAuJ/w86Ky3FKqm59nEDDOm086wIq5
87txXX5TEXiPkDbOTFycJfx7LK5ZToo7C1DvTA7otDZavl+n+XY701lBwpp9md048qU4BpA2YbWR
4gW8SSwDTuIng/FuvGBYElMoZ5cVQ54t4gko/PRhYnah3wStybQW4PdR1RYu3Z+3f5aqRp6krwHN
TDe7qxlAXUmDRmB2RJyd6FQUwswt50WDPeoCl0vbseEdswS2Se+e26rJuy9bmZad2Q9orgL0pHTj
psB2zVf2W9cvZUi8W7Z4MR4G0ia7bol1cUTOK3vUWwje62xZs5Xl8aRWTMw02iPQY1qUqmP36keb
+zIIe7BvIFoHcb0mHJ3aRTbtcok/zudPo7BepHvLiFC7j7Z6i3cmOuDP1zrKgpKXy0F7DPaKZgFY
Fzs5n9C8Ya9EnhtuRseU3wrxDyIFWv+75p3QuSBz60MkCWDvxCvaKriRiQvOzExDifoYHHuAQmc9
de7fR2ANSPM9s34H+/3zpLGQR9qopA7LUKz4bg8R4YgEelmDLShXgmoE1dSuCBWShd1R5WbKnR04
Fgm0UWTyjBeE6GQ2P/TkUoSIZeIAjy0QHZZgZaeFsPzPUrdh1BRtOcGf23tGufeEHLCzmkOx0y4b
9NCpvw15WcH04OfkicNRsreDAk8wDbowe+bIJkXJN7PrITQLcwDAluns5VCGgOwb1KJdlIFB23eQ
fhMNfn2wno2gE+fikRqsSWZP7/nZmXrYKDJ2nD6rTgz5R79Y2q/2MG3BNq/cIu5OXlXoO0I/TIOJ
XCqXWohCvKfbYyqtXCX3bQmwolS2yM0WcUf3K2AMbs+dyIz3hKOATmU61gQsJHdPaxA3UJ0o/2ri
x6aN83qgEDZ4nxRkhJi2dxkBsGzH0xx0urviQ7NsA/Aur1n/y4etUe1cosmu6dyG1hFuom6qN5W3
lH37HZJTVCwADRSh3loxallpPRC1y5TlPVEMkF6SqF/un1axR3vwMA7eY2RBHz00O9yX3urgnnQO
QeuXPGkbsc5nttEQC2+nqwo5GAKWE6URzGrYDBplKAd6uj4FRMhiBsqVxWDMxK+PFl3uWQ4/O338
l1OXAZwHyUOyzkpcfqvGkBfsISkgSgpWHnJtfMOSWcjCjOnB9WGT/ObQuZ6adrZ0UIc+qOmkKEHX
vW1wDErBFsFm4r/AMkMhefZUwRa4Z/0BNOEZmGyHsFxLWxeNVXr4OyXZRH7qnyZhVt0r+Q8xy3Mm
7z48ouZzy72hBup07EPtoc6ayKv34qPoM9ikfZuaaGjA+1AfIN8gkHPhv6LREZ0Qz5D8Lac1ve5K
fAd1wJQEcZGA4D8RotZU6nq3uVivY1oAl1fxHtEZT0x4wqj87VGw9lvux3JH3q5fgIEP9em5zaOd
ZP7IMvd/gDqM2qNqME/xahlG6MJJfQorfvN71bKc7e/3XgppVpSBvB7Vbs8laVIcn25nm8AHSpcL
k2rxqMbyHf1zK5ohaavyKkAFuz6ViNK03yjN5AtEJXcvWEIrrK3sKrGix6EhbnjUkx2P04sbakCU
jape4uRPelLUtV3wC3YOIUk/uKV7UOTWvNzlkrn3Ypl7RhNUn6gqFTY63Oop32NQxIiSpnRuHUiz
WjaZ+CywVvv/i3FML7ZKrPDszcPKiZ2yx07J6MLvy07AOhCv8Ng0GrB7o+T/foXe4onZFJpSP0BS
vtKo+nN7kcI9lmpznNUUe1pxRttELe+Ah8oZFx+sZp5a7wJkP26DDdSEKbe4dH7fIrYGLvvOEYSN
TuNE1lt4EWhPHsgpZJXK/EKWD7YNyi1kcLPcXdaw+ljEk3RtIAaDt5YTJEkGRelfZHgMUxLWCRPu
Cw35QE0VYsVLuj1l3Rs0kfht6MMndsIu8oXe7MPY7lyAbPLslkL2FGsUTzFzm3KEbVxtYV5CWdrL
IgV0Tm18Wvmde6OVABh4u9LabIl/9FVZH0ZME+QbrewThbNON1ebXien152hjMqsonkbzpnv6R1F
NdXhV/5r/OpUk9yWrOfr77xNIUKPeUKxGVHyZn/TmW28zqzo0Hklr0VWJ6OqnbGwy3PXvUZGdp+u
hoaHJ/1bEf4Mlm/GjOl/BoywH1+7VXtY3JKWS7WbFrkCSoeZlBKnudthQsiMZW96yevrgAs5/uzd
dO4HzFLMUe0BR2ttwJp6Fz4WvT37ukjmUDsls5usrpLkDyrxoWdgD9DdVjZVu6ClhzvdXvO13X7Y
4dcMssI9JtKzeF70JmgVFLt4mpBSef4mOmnDDINHtIv9l9gWUBckzml9HKCR6Qh9bXxTG5sbbCdA
hJ6uY+xH1EHH0uk+AnmMRGyqhk1mBy9NVZasB+jGJ/QfBUKwEbRpDQTa58qfhpFY2djnqCH4egXe
NPg+ijZ+4qqc2QQhjbyHyJs55YcIAVwR4MRr8j+QJjey9f00dkiyJUFjY4RbgeUM8ucE5L8N87hE
aYFG+d7RRpOP8Aoed0vjD2SGmPMp7UNaWvbt3VgEiOrFtylhH6fncFHehrKvfddk3yY19nv0hLyv
gjn8mOX7bYPZi2aa3rZx2+olMDA/rIxzDk6CT4QGgYxMLmBXp3xidW34vljaWxzOsTwQkTQz4EkU
ttZpspDqQRdKfYPxR+29A+/gKZN7ous8pMJlRrSzjTrYSR3Jh1x66AdCzpnlmxPy9BqR62VUjHTQ
mdNBumkIgVtEtIx+Bt1lP50DkowsV2IFP3lgzWPVHO9A6D72w3iYMr4dlawdVHnZ1FRE/yDCXbq3
PaI15hnlNumBYug2g58YbBO0N2ghfBEgx1EwpFo/zNVHa6PEn9CtrxVE4LsUAPVENrJzywsFrM3V
OxCS36aLienLgbKNmLJ5YdSW5Pyuhr8MqRTn5pvMRonHo16f32AhZ1FUB4JLoJ7hg9cpllw2mxYk
wXqYpAUW5d163Qpi/cttsGzIG6YKOpo4pGRAFtuHszan0rm0bmA53/q6d+P3Cud+OhQF0b/BzkdK
ZS8r0XtliwteYd1NUN5w3CIiNxh2LRts6HaNz/e71kbs6Pk4v++ntobz6ac0hmMVabrpK0toyzW9
Ey9zLXSVxCh7NLdtBJTrMuhoRHqUeBvoun3XnwNqkrFJAFySCjkciv9Gp/Dh/+HgHHwEG2kdBfwj
qbbfGsvkI0cH5wDnu6P5jhHWeXhlrHbtf6n2JHqP2zG3FawykzQ6kdjkvkLN+HJg+Jm+7RMMkacL
qUrLgg9z4bgMvXN0rUGEOF5O5kntaoC7ChfRW3waPTqHC1gUssh2brifTyXzW5pYaOszy5Zsls9x
LCOvTPjtmLIiic+WUVJ7OimTevd1Cx/nwraSg9NmONDOhObGZqfuEfdRvJrJ4eUu4XQmMs2FxU18
co5vVGSalkXWI9Qg33DsQl3HwvAPU8xH8dqaYPWCj3miWF7X2JpUPLvqFi3km2BqLuyfrEUH+i+B
6p8AleqNTz57lfdZMiRkzCOA7TOvsdErIUExVY7h9RKSnzIAxDaC9vLKzdsPLZ3VdiOswXxWn4pX
++HzyPz2cRNnqQnLYTMJBpM6LUP21m/U86a2LkA1VyoBtSEEVk9GyYpjN9MVJBMyeIXJcfkzlnZX
7rdnPCiFaVu7Gj4+Tfj326PTgmxFpy3sp6qt+a89sYDvgNMIS+dIKIb7ssjDaXxIDdzCR4DtxGMv
sTrpQujzTlNuOjPcNF8aLJiR9hSwuZChpekrUtG90bkIiFO8MwxyOL2ycwpQKtHN5f3rliVPj6Nz
FUQiahptF9LIsj43UxK1DpuIWnEoZaT3nvY0tZczbOCEAbIdCUWfUrJoJBBqMD0WhcVOUtRSqfgM
FwaP8WFvUKqrm0s8AipO9DBWnKWKQgVW4xgqXJ6CORuwwcnvnoA2q2K2irFuZRlIm+FLl5bolcEm
zP8ptfmnSnVlEMSZ2Yb2r2JLiybXTlR9IRbvcmnT/+trgI0o+zy4tzfdr0sJuqdVS1T0QG9yiTg7
ZXq/V33U0fUNNZ144pTiEN+ZcICY6MLeWkUcEjhfxUIHKxvEiNrhStyobPhOXwNIFe9iVhQLpTLp
YO+T6qoZmn8m7lWSO5/2nkC5whfpGqc76hSDAZvaMlzYgKlICP94NUw96wi5KFVzXaLYTpL0Ix/r
+bDd+BEWScSDz9kIF/R90XJbKeJUGLiYTrpm+TuXtz2O8JQM6eMkT7HGvqIKAVvL7U1AX4E0+hIu
q0yIrKL+gov6w1s92BUErLR+5Gd1WgkrBzBZuit5R2XJziC+Dley7iPgF0rRd+ErgNQldbY8Ff7n
GaLTEmB/ur71sCP3wo9qsxQAxENmUAnBayHvZ2SBTSTRNvBvE0NzeBVjFI1V84ChS1eVC9TnF5lm
P7n5CXR4v5fX1JBWcnfv+1KG1uvgMOMPYlMaU6uF76J0+2EyqY1s9ILY//gl4oYo5usfRaw1WtKn
VmGgofuZmU6Wb7mLhrn6TFIaGmGcRV+Am/NdA3OAa0Bs5uM3sTMXw4KQVYo2XrAB6SL9ZOdhC2na
1Ln5LeGyWDrdXPVJksM6W75L8ozCLGCyzOta4kPcRKYS8IyPs4MTcP6PWdmZSmXWEQX2IjsgH2Qv
Rj8O1cBwp7cqhV8yCHJbwgXuJ52zolqw84+QSMxK0tfSGmTO8cxF6+ThcXuEd7U4wZV0WJc/0r3B
QCXuWEmgpILlLIKBKJEJyE29x2uKpv36/rK6YOlBH7wtooZTFZ2Mv18bIe2KzsOeCnS/vcRyRWmZ
VOtPNzNp8RiCU2roN2WL6e9w7/LXWRFG0JrcgmP8/9ufJWlBdoftfi7yszuvuqNcGjiufweM2f+M
pcCI/llY4gGL3ebC829VkrKtghIz8P/nSp+HQ7CFoSIUgnZed+Sb8E7q0DWLsaBiSUbdTAbheKdX
A1DF2mLlbHqdX8DEafblSwEiT18GKMj0IWcOPfV/23e9ZXHePH2rLME0J34hNyoSAHzZinXx4iJr
zc2Gvd3B7xltBixhzWhERS5+5N9mm1tDAYPIxczyFzd6oc4cIBxqLeXIZ50GvO8N2EpUlh92wYsm
uXnUpfI1cAnvNw7xOJcIq0APMnyRd3Ab+IeFPnPu35hDcZtRspY2Im1um3KhnJ0peE5w1A/gfwJR
q9/AgtxW2s5ubOzrs05u29C2TC6gaRBK07PUGLUVSrcrkr8+UGZ0dAB14yEJAXJkf79nO1eG/tZH
5SSTPNq20ESk0Qj2NsyAaaVVx5/vDzRJ+yQCwKN0OjYj42DgEWHKQADTUtZdl+xrgMZE/Zr63lv/
PG6BkMGDjjdf8YWpJYmETYYdtKl72Tvja9TbGKBiCSX4N07q21+3LZWgaFWT0Aq2l3hwxuB5a+BK
/Fwqpv3rRI323zWe0u9cVGu3In/jswn+K+PVXlR5jKPdiguFAqtE7w/f4M5gXbVvyDXYSeDf99go
cUCJEOmilAcEZK2nwi7I8kN38VcDPFesxckaPrgIAcEQsunrk5jqe41NL560S8id9X1Sbi+693gs
ti0ngIBJwIszQbNqOG/jSG9ai+S0NZ0RkT8Z2pST4MgXS/KDc16Ts9Ey7SgszTDal29fdZaCtRsx
6tqjrkN5GaVnWMrQgKq+libvh5q1ISjC8pSyWLw22xMI8O5jvjS0ywfLBz412E7gQ6rBFyrQwE8q
WItdylFtDNoBFb7CreHxSHTJAhD/NPngxTJ+a3mnVYsiyeg7xsuYorgzxqjuhu+W6kwEfvLKIGAY
bymm8IFh8lhsmiBhbXfrrzQ+lXhFjtbeRoVhXSObTWr56MOKLA8XeCwnryDU9iJl4mWWq8Cy+AWV
sN4ws6eJmn/M/pq1b0Kyvwtwh0vl4RJmxWtapt3RnOjcGIomGtnGWjQYMO1jd61Ap/g/SzeewOId
uU6YLK6oA94V5AJCcrTGNQa8OTYRHu01apjNS+XlyoXV1gAksMwz23ffEvpUd/QxqvdyFjTBJaRs
i8sC/nWTqmEFOeQ2AgRPdXg0Rveacae5HFoge6YcgqcftGj08nWkgDcXxGD9pCSUwpwPtSaSuf2p
5nLA5VMHb+mnOUW3SN/AjWW0LlHYFQyDMHhUyrrTlGYufyIdgLnu0ryflA4v46u911BbXbG9K8Yw
k4+nwjttFqU05hCXqP1hgj3akUdkx3ChxbivrgltK850vOWRgehckIlahqvqvCCiwYzdZVSeI95C
FXB4cJQNrdUhjKsnOiBtaORFKKRgGsbFyEiGakwm1ARckU4vklmrQ1nA7VwYc/rVGUk8+8WonkXu
a48656BeWVXH+LbTOYE+cOi4NOpp+oaiMq84FwnyCHBM7l99uEf9NLUGGzmAGkfM0KV3n6VUkjYK
NI0xksUQaldbHZ/zjA+F3nAmiiIoCPuF7UhaWjygvzlIabQIU8HZTlHorifAHRwA7owGut8TVKp/
OlVbO5bxXX01HU3c243swQa21VRQ/smGtZ0bypsZ6t0Zqv9nmQG5YYmDXW+6wUSXz0Ml2/cLfuTC
6p/ng3U3kCSgh+dnG1ROuOkA+2MFZSEkofQu1YHNFhrg1XQbTshHZzdU6rbW07ykTajtDZAEmU4w
a3ptXkHupj4xLBeKkfkYWMhlJ2TB/+pRBtznyaBql5XrbYZM83p1fwHIC9wLLrag6cfIxyXq7mJQ
Gh2zD4O+wu8ScltPKHUui/MRHanwx34nMeup8lVqd3j2dj4ve6X+bbd4ssCam21Bl2phWLlWnfR4
s3S4wiCJPaWkzw8SWKeP8eXBsqGWitQqDZ9s9J55bcZLZjrHre/1Pj6nEIalJLMO96rSvA5zPZN0
Vk6akj1qoK/hTQWL5hN/6lfDeamjtBsWLxT47Kf0Vnwbw2gEpWu/LhPVLvDn3O3+4juRJNYBxdIG
1Ar4+p2eBDsGzRTNKYtWye35rghzFnp950Y3H5vqOEf25o0XkVQjgiF32eMraeFUgB3OPisSI817
TbmtWIsBy3qsYy/GFDIfKJaR6UU31HXu9nkjfrtk3ZSqmMXmA4qoQimyk0XxAF8LJtVEgwpQEqOX
IwydlANz1cxakkNfUbsX6si8K6z3gGrShZW1TMKF5ZpwCAa/FYBAo/gNlM4dJtvwfqksinJOulFK
qICMZb/WwezwPmVQZgJuNzc2cYBkAAaTV97gyItTjGAdXPRQ87Jkbq/4PLY+pF3sxoysBxBlngJc
/rMx8IXX0i5XFwvdSyOnP1kgAhA2QtE90uPdtQJSXL5YyMRWYQ6eJ+/GCj6+LzlOHgDxEk3UtT6y
cCLoTcJ5jJ8xpil4SFqcaZcGmB0M65FRqj/q8IH5w7pvfdprfS0Yrxv1CcCZmX7ganhV3mDAeCYz
lOd5Xpq3/nHZlObojcDioI+XOMJZPhKKFV4qsYdgsMbPBysdpfyS+scTMi32abgJ+ZNPcCEtKECk
oKWHmZ1Ikk+OOYw5V4caNwJR8bZGSxVadRjS8YzHC2cfYPHn111ubEkRgMvapO+sUDuraZDYt+Tl
OLslVB0yyYq0vOnr36VJhIaXsndgcBxsK7np86oAvrRoB2sZsnGrFxlyrvzFW/cgs9wWvZL5YrJM
byC3zedpzXCrU8ExJjyX75aUhJ+vQNnaBovIypQ01f7gbri9ACWDhoBYpSAmrowSpto38XG2DqM/
UAHL39VDRja9/6Godf+u+HDpk6UdaPRQCPLsBfmdSf3X1cSXjva4oR3U4ndEil13acbwFUVAD7dN
SOfjw5AF6S+ryUJKcsLIXFbCk5ZMQstF4lCR7QIKaou8sraxFCN7pAncWxVu+zk3ICQl9HPct27x
whiVbULccuYizmR1VaQlh4tjwK82OFvT6TsnIo8GBzyZ6WdsYsmKYueh4Wa0KNK1AzVjuv83U1NF
i6fBYi/n3UtasCC6eZUMUifGch+cd4NBG5OhE0j+xFeP5GBmjOuDCVpzOKnmozcGs0trM1S85NDR
5UV/uY+HNoKf92GVMi/0H8GFJa1oKNQz4NCFiVgGUB7DRJT0opGybiKCtmj4Pp/Qd3SQ8gsFcpMm
yHtPqR8va8wHUAP+nhXx985R/tCVHMBFCn1kXKBjhWYs5AuAysQKBiGy9j8VS8zhfsr+Zb4J3KI2
dR49RR4L+RM5tPvar/Rx2fnjGlDPCo5U0cRuDXVnJByKZTksUOfIW9WCf+hhYEGXbPhjHaG9wGRZ
c9p+5NP/TXouZ2I53Vk+c9V+y0EyCze3Q9KUIj1DCCnc62AyVmILwWY/erqwDNcN08P5wd4Ii+oS
YDBUjvnOA/Q568oFZforf0sT9LTWIR+CCVq3SKCSGkIUlS6g7S731hxzVjoSjnKpDNsx8GdH9YSw
jMtmfRSMu215UA8agu52fo7jdwSJfVi1fpwekKhew3z7Pgf7vc7IV9Rk7/UGVFPlDBohD9AkJePC
hORFBThviq/Vvw/zFG1JFCGTrmRrYwEQUSlD653lvptehsivsEdqWM8htOu/7TxZdrvM9qQarIke
WBn9/3ctexrmta1x33cKJUA/afy3V93g1NolFsFW8d1fe5BpBgBqYHV2+Z9/PUr8tYD5OqilEj5E
iAB1ue4yYzNptHPKzElqnuoON92T0ja5tGz7islSrU+zI+Q2Fj3AkLJxrbOoplxEJhE8rCES1ZsY
zB+sXjo/sLxOcv109BT4gwrWgyXxgwfta8Z24p0lrjwADx4cGlOsmWci2oBhhQB20m/oEkgn82jE
eCj3YE85V4G++868tkx6nccr82De0i/eqdEl1CtBiGNtLwL+2w41R2cy7tyhMUMW/2isCZ1wQjn6
51E4jD1qQgjZYMdF3X0qvAz04K6thZLq1DMDXMEPr5HPIjnLzcf+nAJZOJJFj0GvqNOu9+O5+ekG
n31LvZfcDbWFsFEzvpHXuAmszdV2NTcNqn/gQVW260nHRvcX2QLevAVR+qPopp6L2K1NoKZAXspk
ZRHRhF9BjDZ9Bn9jUMy3sXMw4TS1s8W+MTEBnH2FAY8QfdKp5skLMZf8pDKXYWG+2Elb7+GmvIZu
nntzdIhr0P6YEEAtPmPINbmRRgk8jOwtq5PjWdQ/svhzQYxyifCKLI5OaLR3VDwmuxgDFojDAq09
iR2PvQ0JV7LbDd1xMW+j4THuzztfgcm4BM3iRPAfWOlpbaSvBSPRTBF3SZ1VKmJC6hTe7EOJX5VW
sLitxQDbLO9AR4cy3XVrAk7wlmQnbIPdqF+yOUX2t4HDt78uc77gUtI4A91qtt+K8I7W33Ig6HVa
VJXLcRgB1drUIQ3EDl4oEwHNyklWqqpvZIIB0qDcqoUPGKuFfotByJAOTVfMrtySXRKA0rnGRI/2
/xEQA5W/P8hvOticd2upJ6XEl+SDFvIcbFWAbGEbHfOM/65gJGZV7fmW9sS+H7v4k63MXZjLK2bN
LoqzWgC0evoulRbN/OPnGAdzMZot8Cj30noVTY0YeKmcjWLf8aLs7Y6Oi+qlnXhwv0o8Fl0Lls6y
Wz68PwoQaRcK0jpUzHvPSYDprLZkF2dISjLzfqGXLRpVoHBqSewwJ9ouLYeKncPqJg2Mu9An1mnf
FQT5AWu8CiNtNQspz/7O1mxMap9feIn0ZskFzVtjrmAvA8nWKoJa9DAKCNdPdMkkFMsdc/ZU5H46
OqO0btqV2yi8OnLYjbOKIiTk7aKyX5yG+g/ZYlhAWrU7RGK85Be/n9pQMXfvEyBPJakH6+dIxdvT
c05h/h9QtKplOuLVYcEb4t2zLRmdeiBFdR5yqfa1q7sUkwSs6lnOU2otxw5+kU2sI2tZvF2lOAgu
ZhxZARE0DYS07HYJKMmI+DI6wBCrPSOco3imbSDoxo1I5TqcOCxwsmcIOjkJZRn4ZKaKznfiOR0o
CuUsh1URYq1CDDeRPAR3Xj1sExqWndYfrBBAIaTbzCSY7XxJTeFlUfIv9mLJhddA9eNjp3Bc1Vke
kOnq/DNRXn3hKmOXIHcsKleoHI8IP1nC/LOr94ub2fNI3mBKw2TZTANEc6QMJIZuntlOrDA3c/Sl
fXAve4IXu/P0XT8+OhZoj0Ggo0930WaiOVhmBM1+fYPHBFRIXCHuTpxkCURCNPMa+sWSYglW2rQC
XiqFB5BcKfdp+wZaJNnLeDJphX1cy86d2qJO9LYFqEyQfKUGpcsZ5zoaZ2tqbuMQkdot066RseaS
k7b75abTTYOM50ohSAMYXWqF5ZO9im6//FejPidHjXRCa/3rvWymQj01+IkL2NC5QrP7js5dzozP
dUtUQU/H7Sl4gnMGH0wSr5rS0Y0w28+/sv8gSHJYQ97yf17oK8WCUjg/OSDGL3nPsGhV83ocA3hB
lI8atRrNMI7gY0UaQHFILrgc6bcCGZ5fJSG1WFLZZ2lzvBPlYicxYQHqh+cwzU9PIoodW6aBzLNz
fNXIx2cX4Inui1JPSZ4Vy2Bf7y552Qa3Y12XaDalnNjfOx1OCiGPMVbbuSdmkxtUy2mRgHDOCCoe
ocNli4Rv+Z4zzg3evOa4tgKl9aC+rSvTn2MJhp9qXL1Cbhy/Rbx7pKl62zUX3gnhO9Y6/Y1/kqut
7Q/pdDhefbwHZnnZ+t4Xl6/nDUrg+Z+fPkCEvEPUNgRfFFQqTtjoy4tih4uqgn009CBbDoM+Fr6B
0ynwxhKFFoeSL1doHRXCJkCEhO/2PVH9CGom6a6ExsTGHiZzDsqajQIoWrxV874QXtWgj0GnztGB
HqK6LnZm3ZgVepmO3VZZCHAsyTwuIzmtr2LtGi6GMNji7O6+75C2J0z/G+pYu6o+z7a0CdOSsY5+
xeaW2b+XxGAcBqHbB9WzDqujDB6PM9GiDcxDFM9Jos6aKBhjXJZKd7GmZHzH2cnidx8dGGxN57Ke
OP1oGy6BKSZhCUitxscQXN2HLFm+YGlcTsIcKaTn6Wt6sTf6mMNNi8sIHgS2Ql/WIw0BUBrEOtBb
yGTzinbIGtmLKbJY+Tg0VsSdyb8DQPKBeg+operWmoDEfQDf+vsPfSBLEUuBAmkjw1VujvJtCeAu
/C+OaXscwXyMJ3Tr9yfDhS0xyTR/OdGMMtNmlKgAJPSSV+ADC5HdBV3L5RIUtrSijHXLDckwORGl
hpGmcxi+Fzv38MNA/DPa/8BD1Q48O9ZzEHKSvP7tm3zA1KaB+EOhDuvk1YF+XVeiPjMd9PCu0kyU
seKIH+aLJa5iWFQFGFoxYtaRKcPIEx/EjVoupOtP4RUAJbXN5hLEwpPOH7Fez/q7sqNcO4NHFHyi
Cc1tsv0vmLoosBMvO7cNgInpHnEKTWW0QRTPK62xMi/YpzWGtPn31ZGaQCD8oujQW2gCE4tS8sm4
asl5f5OlnYkLyaukjWPIHWc6rcK/xVK9M1G0fcAMLiR+XVyPqBiVr5e5qMkhSR7LJQWeP+fsnX9t
GWfkKPoymzXwsTcrIKjV0g+5QQBvXeJf/U5zvYEl51IgNrDHXdGh4RxNts3zM0/s/WpVJuhQOyDa
tAcql7AHufELl/9VOSL/iG7lIBrUeYmNyqcXYf6/BZaYilopd0Hk52R/m193Sg2gkMlITLdyOCnO
Rxo09DnsI+q2lIAuD8SN9MDCVtH/Glwy0F0Yk4bE9QnQo6ZI09VEJGlwqrLs8VZSaMWeuBu6N4jY
NCZef8mTjsJecpfxCduNpTlVHk+htr5PcDgBUHB/PCLrctt7oB6QVidk2uFuw3CdRqBy54RYZQdz
WHBY3FRukBa3IDxX+w51XDl/ja78iPnJgn/3Sb9ZWtPpMrGpXMsHI0NhyVmGqVuTHHIgdDCW9Yis
iSikj6DfwTlFFTUF3PfD7agAq1sQ3ALcxOnp1xO23xS161uTv+8+pLmiQ1BsKxEihcl8PaPuo5mx
lWJOWTF//YpDT3+ANWdKwPeL151K1n9EkEaNilRNpDLghCVKiL4EHQCob7JvS3axaEbGm5vIwC/0
tbJhXJsZv0OdwbAwtpSXBEXlec5qbrPDJu8fqHzUfKL+9yMnyxIwrUOZPKdnLhulp1gzOze2s2ni
pxy359f2r3u8IF75Kqhs62BjyV3ptBnhiRq6AcauIKsf9D0MscJzgAgpQt9htH2zcLVTCm5/ArKk
gUtHD8uONXxiHKdu1Bz/823gIwEaxk5phdB43U8ZF9f4ma4Wugq+DRsWcxgenrOtUQ6IDVrX/tuo
080zgJm4nU6JipWSSlj4LcT7AOSWeVbQOSZzQgEWyWlIi83EC+bhGQU64IzokObPmZt+RnYeGOQi
CyXhnR7LIlwJrysRpY9ZUiAhKBa2/9m+/8r29jXt0phMNDuCEJMUYnBBzc47kdmmgpaWogZbG0vr
mnZSWhtQVEpFlbTY31KB+UfdqlLDmFl7NP5OlEr8gqiC1kRjjdsjFMlDdhW8qiiL81atScrSV/zh
PgDJffTifOjaNNhlo19uIaWNU4CfZCkZe2Bdg3sPraHJKF4otn1FJNNosa3nevPgY4LSTmd17zNR
hoxf067PxKJFi3WHLUys2t2af1qGikM5lC6ukGJlbOWH/JfP0t08CPC9I46XcWxqEwjt2iCbATQO
prpGAKj19/3WuEYTO7uqNAR1QpIGHZqxAMgVCoWOSaVThxPF07kqTHCkFMCDiYDhckBt3bCrdced
xT/dafxQhXe2gra9sfasAaPRwvl8rJ8+0V7WMNbJ1db0UtOyC+Tv8wI2GWCFav6V1Y9lDcOrKL6w
zw7hNVs9mWFL7XbCmjFVaKB2nkwbnrODpTP1zOYd/zHkR1g7tsTZS87G0Wa3qfRPiy85VXeC6ywQ
G0C2UgticrQRjhPyofEdjVAAmVptaplxhaKmSkE7RhUcLAXT2HKASx+QCXOXyLTmaHQMkY6+4n2g
oV+fsBljDuoYv7N8pPRRDjeQfLsb3KULR0K6dHxndC0BdWfZBWEeY3iXTx3ljzdn3dW3RhAtBbgW
9VK0Mn/f7Avm/lRN+7Lmy12iaWf8NGYwZ8rqrK0QfoDscZtvcW1koQspAk95pNhmwzXDrtmnYNdk
76DKnUEf+CEW4CbjloFuSnq5F23YpECKIE9dNMMFqzp3v9SHeKkiQ/VGjBSeMAf5JCOo/k+8vF4g
SfGyR+n+eCrBWGePL7mcL+2omFhPsLStM8pietx2yMwAxvoc3uJLYz4Dr8qr30b/XbdcovkbmhbF
vWsuPdioE59fA/tQrMnkphKSef5qnAJDLhMnTIbIolBMxEo6806AogOlkf+cigGMlDbFaE00n0en
kijvzhpDKNBnxBDuSJ9nQ8zs4z0YIgIie4xBU3lUNJh902YFnzpLJoyBAxXpSnPQGgEaIwAHHM16
6X2kNR24t3516rB9CUpiD2w/3bergEOhT0RabJflPHPKcjeW6mkVMnCAU4vHmAbSOsLlH1N3Onek
smRtluSyIzQlZr99fbnJO0lXE/ACwGgvhz4/2nK/2tw1PtCmXH8VXu0VBWmVOMoTp1wOaW73e9lR
XdYe+qKpaB8qPOulAV9OYoIJ5wBoHXnFkzS5jb3JvamrPg8A5ALdPmKolDT+M0hFK+qtwZ5CDpfb
rkD34zSZ6PD0OwNPdBr0yYTVXOETXnSgTK/lFmyw+ehPqQcUZa+Z+UbqC6/CJ3C8o15Ew3YQfth4
f03vFh6CS4+5H/BA6cpuuvX3KFnqYX+Ix1wrKw8U11qL+V4ASZGmQJsvPfeHKY7h1itLoWG3uVPW
2B3a4UxjklJxVSje5QLr9ZmN8bvR+Rk+l/9G6Lri1j37W3fK097qnw+HrsLG6KvG2p7hgl7Od3Qk
0/zlggsGEfscv1K+Us24pAR+Q9AWTiVB0vwFajP1fYmiJRWm0+DLDUImcVlA9QhCOthAw7XYa6xu
nJvUCHOLWW/v2zxKCJl/thYdptDOUB2OO89s5FqKcYl0W2DgjBMnh3siI9NtmeLgCF7VdYU3V1OT
SzvsY+e+1IeEBTQlARie4Vh7UW0TAfhyd9zu+AEzPZRsVjJBWQSbcxZt3njyHLr2x3fQ8wrEqM0o
/0Y0r5vmlHTp7Nv1yP3LwEx9vFC2HzOI5tbeG5fJkHxqOQpdgd0SQR906rHN5ALYhXkAQLu+k6Yd
l/cRHy+u07vnER1sdsgFNKXIKQPyYppXEcVe2NQAn4rAqMZMsefmHaPONK7vDmp60GqJemzUnRYy
eBeV0vhFvqZqDuJuTmVUHNv8Z7uqhIpxZ6PNOtR1hViuE83rkcEdYJ8t5T/vxuQ9PO8yV/gwxNwM
A9ZcpoXBprIUIPO/cXQ7vOoIhJXgokZREyJwa06A66AA6T+l4L9Sejp0EkoA6P4TAo3Q4vdI9q0i
RtYxNRqA5d11vge4gYjfxkFVZaGcCZr6jYVaAALdgYRETTrz+BN35m0kUCiPXXWxmwaH1A+RezBQ
aDPdKbKqSJN9Kx5QoGUg8oSFd5WaoBLYY2ZFzY6szhbyKzagQlkrPs7xhNSZVXB+l0/Tec6NjuXn
XIf4OVUrxfa+ywIB6460ViSkJ/DaSRLQ1PkPpMA0K7wudzikXqNGYaX+a6nFYCAk5Mf1bO1cg9B5
/aRyHE9NI5xKjG9DuvmnF36OLi5DB48PqWOTV0TxnA2ApPv/gIdZ77Wwkb8K+tMs9n4T5wcy3VHM
c+Lfm8MCizKRpVZbzzvE6QYkXXRjxPSaVeOeZJZw3BaOthRr4WT3+djT//uLIxI7TPr+32+zBuu3
Wvbun9qEy6kRPQFcOrYJb26hXbys241nutj3wznlxsp/DC5hD4O2bMpiiDpt9mMIdvJkwJFeelPd
msmh8+Eoq2At/4/lZRcMW8ipZtKoyccA44nAnJSel6QK09X7M5qsl+9GdC8JxgW5uLQOlLOLm8eL
tUTf+kXog6kP+EgXIJyyG4erhJu0Bnohm8kYMQSMzxTIFGCf6oM11EYnkLXjFtB/9Nmanhp2juth
vVkEUhojPqKY7lf5Kjn3WBfZ8o6bnuep4vGrR6QpTSQwV2iBYKc7PFq4h9TYolhjPpZ4N3NDlAkV
KMviGyCwCehlbFz+SLgTAe7XVjSSlcb4LnE0jPrHuS49QSi4GMf7zdEZt1JUSoQAP3XBIj4AG6ri
jvGX+OcVApGNbBoPJz4j9miCwbH4vj8nrK4W/j7JC36HKMyxGB9wNuQyhdtEEAVfuDpLXPYfwUnK
x5QyfiaSMCLZjA1ueoru8vkEpBjZAtlwFbmg8jsv1AkYNmKatkSzGKVzHm8cSkWt5LB94dp8CSOj
rOwJR2+UZYc9VHyUIfF/rVA78mhSG9qM/yercNVYW6DrwKeLkZgvF6yebILw0q62xaaRAXqFen1g
WaJ0Z7NOZd3434y2OqCnKj4oW+2X/0bL+CrieRblb1ua1vzXGlIgIRUPevKBOG7APEm8BYzrtdQp
zpQhx8qWgUXtizC6ZhB/vuIixZED2uZTUIArWVeyYNIBUErZZU+zLPVfn9Jt0exmWcT+67sFYaOt
L831I4KDdeiRFvlbXadEUw2CAn3WXbzvxflywpngmcnLsSte+9i51zfJO5YcnEg329dXHnQjPX3q
mjB0Jt3aFvOY8lbDc3I5H/hTsLaTPFqf7rF21Cs4J8Ipz8jX5+YAGSnQG39+MA9WsYNTPXT8HRtZ
EChLvkqLFBzk2szyZNQ2YVU2DVNnbmtxh4QidvrAR0k2afwLpy6oK3c/gSs/YWrYiyLueVSo7PDl
JwguGbZU+ZJSxcSzl/fcLqQjTE6js1up6xKWXzX84vJTT9rwwAmSMFPTJ8V60T95UW789Af95lC9
sCeGcO140iAsiVL08XkppfJ8szcCcLENFuApyEusObgP5WmBMQAz0TplP6nZuXmjRtFfX2eWWmML
5PHTNjhxfghmaqMx/TEs0yp4RCef02R86GUinPJYwLQE/zJz7AtgjOBjBVatD/PxJVUVIf5Zy/3F
YxSpUXDMmld1yia8k+DeLgFHAl089S/cfRG3e2pTl2rXJ62DgF6iNO71HfiFH/kk70bbx13CRgdT
Cu8T7SLUcv3tzIA5R6xgDNQT0OSLtBPwiSvsslXu80Z7L1J1p12AtVl6aUD8Y6vSmxSMQYo4cAUK
FQGfgrqad0E3qFY6k48n0qNPgnDpu2Vspy0+L82WH983KjJmMcYwfWa3/ghVvtbpud2F/ntWert3
GeGZOWuH/KWClb9Gb04nPN9DtzaNkpH/inbVAYFoKjUaWQDGlO9UTyq7CEZSgyeAntTOAxdajv6O
3HBsd1Io6PL2NUgnm+BG0+dD2iZwlhL79Yzu/s4jXM9whGU/Y2FeYh3dnzFvXE+vdB1BT8e086Xw
AsMrDB68gO1MlnYKzFstwiizHdYVPyg/7u8bqxOmaQxfjGPcI909IdPyntsCN5rqKCYJ1B6bxq0M
BjJlyH/XIX6YQwYt9Xs3aKSTC5diMLUwM58AMeQJ6rIghYsH8VK3eMFrOIFdPhj0equixOr3MB8A
Xo2Pwng5BoXIkAM43+3q+ll+Yra+eTJfSv3/FPcsqWBJewSWqn6YsqR4btwFAB2Jz+Rc/A2FVpr+
fp8zBBQ2VkOPsbVd7hRA+xJiUJizKaW+1sEJUOD5b0o9EvfggxV/VvAZfHZNKPmf3LqMlWXax1Ba
/Vi3z+0890z2nQzA+cn4G3KQHvPmXLFXPf3CX4e1ls4zE2oAEEL34gfJKmM2OXtNAmg2pSAbKwml
tasAGcNJzRp4lpvWAWTEhKL0uI3eecVaeLtIRhCziqhMKbwQTy36P1+6+Pj4zwaNu+hMWGpXl9wd
0ji9TRwBru9WOIOViQ2aTIh0cBa0x/Nx0dsIcGaxMTlgKoJ4FC0t5tKParD13KKp14V8MseZSqOj
8mOPhMNkk8W5jXzIqChk2tMqCe5JTt188BmdVwAWUpnSAnSv250sYHijDU3CsdWtjXbbJR0QLaoR
0//e7L1GQXenEYistwsbd6vai/7SS3WNnJPyYYTANzE8B91NRRvnDMzFFJW/AoUAvIoK2ljzjFme
wSAGJ8H4Ve/rhOaBvTlPQebhZuWrrCiMxed19cS99gbqg7W98W2vKCdpJOCPMi3aBQSsY3Z0vi/f
Sihmx+yH79mg3XQZsDFttIdGP+1nMHDWwxpAbB6oLJGpOGWKAUQTQ7Z9SvUr4nawYt1t8sRq3CB4
D0PD//LwTPDgjfb7BLxhZWcW7/roQ0h3076Ie8I1DAszIYCMxFCTYDgrgidSO9lPSnmcSBkqHXPE
7ZydmgqpvF1pIUal5U5nLcLrkqhFHgrzHUx+Cb1B1WyoUN/KYrMmDOrsWSsmbL2lr4avhR7hJA+7
Z96pEud73wefvWBM/K48ObCvkGZtuV44PVtZY8KkbJ1L/90EzvOogpfCEnd7eC38c6w3tf90SA1B
nCdjwsX0h3xE0fKa7vzEMVD4nGulzeEjIUO6UCKVRCI97TuoaWsS4eyhPKgLJigUpofu+bmFrwD2
kiSKK/Vf6yDQQk9ut1niW8SKLD3RCS9dYRlUwitTB+cfbOuknfacggh6NLX/qgcFkX43CTyyJfLi
hInuou7bYS0e62a6/1o6TmcpIMABZmvOM2UHx3KJfnnoQ878fBY30iV0JnWZ2Kqb5+JbQp7JfVJJ
e6j9DuGRbO7kcu5wfJwrYYQIzRABvcAAqpbyojVubf2xy6tS5m09HgpPfpwVsZW6hPRxLXMGvocl
HXYuP1Ex34SQnRqrybANS9tz4h5KbQseOJRcwU1ZMYWKp9p9RZFgpGH2vH8FP98f+ZIcow2WDXGb
WvBgx+wF/Vq9xlgQAP39zIoprnnc367m6knLKE6iM57LFBnN0E23AsLL5M2eONWRkSquOlF4rCoI
4o9+74YAuR7O2VQkBEjIwkvNsVdKOg6Fig5v3DxNjv12nShGb1V99wrPAnetKYly4EhWppWWApsd
AvVe/YVDFJE9PhNRjZx2BOQ9CokW83z7MdbO0XWxYFg1PB6gzHDCeYqezkFzexELuKZMsnsqachy
r0OR0Dr9rgV+lLDjHbv3Ota/2TyTyadCcI51/KqkrtxoNLKuu6Mw47+jR/W7CL8fsm8rr6+wV95q
xuJVh68yxe7kw2e1KXphZ/oGrco4LBZ4Mk+z7wn3suL3nORwH4xA+ODU4wYaXYsRFVsVDA5Tvazh
/BXnvJzWPs285mrDUfjrsCbJu97YA8VW/IeOlZHjznCCFblhKKpHQL7wFkGrnbID8hFtS3B1VoUQ
mhDK73mfqz056Gfqz+DwlKqtanEILfXIQc1DhPpwAnb0q7gf3QBF7bLOrPq0WjUY2NhXa96UeU6l
VLLFb/V/uUwIv75bclEuWJqckYYXXR9KEbQhwX6MWnEcHXNfVt41KpoRZOgXYFcxSx6k22g/Uc5+
k7EyecmXRYe29jeMRUbBix/csid6zh1xJe2LdNgVoE55F4zXeUFZJywMSEQD6TISKvK5d9sozD/x
xqEzYZy7vwjDImW3Tvg17riLq+XGBQWaG8MfHB4bmZdFkXCx49p2KUzcuWjMLBNA/Qa48gfcUF21
lxheXZDS4NtP/fBRCfSi4vuJ0AEoxnVFyVApk4EPoYmXKSOahmjleBhy9q9wR1eFWuGPZ0IRL5c3
4eflgjpAySMMWQ+H8QbBC9Ww/K5Y1rNK9PBDmF44ettUwGcMp+8c76P6umIQHgcLvgjCXTDtnXnV
ISrgB01RcNl32Y29tj1JuzZgoaQLxzsz1ZU2TOBYJN5ibqLBeZ04kTOPMX6lI/9mwPGMSZ6v75tu
8hVDp9nEJWcV1AzMKsa5GA6LYYkc+njfiAAgngUzazBy5bFJO5nxL0mx5lFWokRzPdWQUY8UOlfX
VQ8dzSEkf6uTFaAnw3JP3L9hSyvwp7LEx9kyspahTzmfCMrmiupsHJ8JPa2rfUFxBcgexZSwbrVZ
Hp1GsSGRTy47davYO7MbGrBAmAoUJwKIJyKNW8ArM6RFqvtzHSpiMl91SwQwXRKDdB/79t+lADsD
xSJRgLFmPJoksGfXtsT/GJgXCagukkeEgIAJkyT/E85k20icZK0jwDGLxfa3rVYy4NWaGpJ+n7b4
eKi8K9rVLtT540EPJwmEjsQ2NpWwEYRGnEdOZsKcWSc6zMCrFsT9EVBjmMz0vymgwBek09U/TSO7
BXqZsVgggy7kUJbbpctjzYqWpnbmsx/ZnvRmjwqKTHbcxEj1RmoBAi2wVvpuU1ASXB96PiE6efCR
7sLeGl3DWChPzCEyAZsrLVCOWBF4O8ezzZhfBAMs2H2VkEeBJkFiw0Fm8A5PFq/99SGk4zyT7H6f
yxfobDtyrts6VDC68wfILlcn4ySV+kc6orWdivR5NendTOYlMBNbBlR1eFM8JqmhlIGLovE2oPD1
sLwi5tns5RZ1csG9H4hCVN+1/T/dmHPG6wkIUnD7JocDGsibtSUBdghQE5T8dbwzeNMfhqJeE54M
0rFG3yoE25Pd2QPjF/zosvxnSetakhiWDkif/GL9/aNub+6bIQ9J+KSVMDW3KDafNS9QYQqu/8hW
vR0z6uyfllbLCM0wtmWCZzoiFzq5fZCCxAC66gw9fOSXsJBf7tzhZd7Nj3nkCOrypul1spbaKTtm
KnDUlwK+E6TsOlkBn7SGXN6owMPhfC9rV27MLyHGRrmHO0uxAU9wbnXvKbnd6W07QSacJ5p16q8n
EPj+TlTrPU7YvkTM2wIjq9O4xEuPSBHYSZFLNFPhtOV5wZCWTObmpINli3MxZIt/izZ2YOrampa0
qldE96r4GeRuUj8BapkDO5zM2LgSk5ih0csuYZmSdgacVmOF9wK5DADnhU4Y8eK5WVFw13SWMivI
CloExs2/wvxahcqAOyR1lAn3T9XPvy7QvNrk3vxm/fQVtiCuYG503ejnsVskqGsJA2e8Lq4BOhPO
V/CmJiEaJXjZ2O1ZIB+Mgfog2oUGMV33yrKmaSqfre7VYpOP3IE8ll9C9avE3h5PrJsyh5hUmefN
Ka157YX0WHxNaBLKAJvx7vxHZgYJ0LX1OqOe5JAm0zlv77/spCRpouTBzlecWbKuTZAjAdIrnEQ6
Z1DMEzuSBuLL4GSEDc0UFC9TOI6MFcoRDmXiIKihkv2YruxgUel+EodNZTDQiW/56Wat5zYPMSfw
8YkR+bEaVtWWspAOmB6EJxLgf9fCeliZsibKoBjbA0UXFezP0INNDlsva3U4WHJDpvreaYJaejQc
FS6Hppv5iBzGiXXAmPcTSDVoKZMPrAPqBrcdf08EFuq69TTdZbvY1dyIBxpZYTP0z0ZCXtmhKhyM
Zq+FcFH8aLbljUYRD2fdTeRavyuIUuvAEi2K9GujPjB+zyErO95LdOSxi4ovumH++0j5PS+FAHjQ
Q9GvoViBvT4hG/vaTU2qCYf27OcGd2ozsANanM5GcYdbLMjBWT5Vh+fAVY41Wx2NT8zQZFBQ4JF5
xW+dzYxd3HKci2T0WMxsVvWzdxYtWTC+dw+EIcDF6J88qAA5ZFHOkaXyIzbhHUuuzlrJl4hh5LGR
pXpSGQJOg2xXkyDnFbnUTRSrkNv9SgUhGDvnLzVtz0YmcVa0BrKvEfVo84V8LR+/teyIMqXg+zJz
c31dYIxm0m4A8FYg223b7P69SLFpSmyA38gxqT9DSOGytCim35R4W+Ond1weVjG3dzobaQp2j/LN
RjEXy2x9DSCSEcLWF4lp0XvekOSBWaxcalizTzsI0Gbc0B38dG4QfVlyb9gn9mVFFnL8FTiLhoCF
49EuW2W6aS5bGDjymcPR+eLAf1Rc//d8/ZfOX9LkbwhxZwS0lFC3HvyTti6p7MoX52dUrO8a8GiI
MshM23RY84B38aA+IWCjL9YW7H0/l41szQ//zTL82xCy5KulC89XXGPjLvYB+OMaqsJupNAOZdb0
BkX6A8rGMpni+urOI5Vv5n077jq61+AKXlEZoPEuEt17n0CRT7UzKZLP4zYiG74aLSy5hXPx69Wl
LuXvk2zvXaaVH+9gUI7JB7F1cYrfUWqp0Mzv/zHETpJ0y4ZfV2vrXE7ZRyadbSKehorOjARhhTCT
G3yPtQywI/AJPPFyAi1RHMqUnNOzEnbHBUVd8TQJ6YL0XuHkOI59PF4PSi/2JtLame96Qk5vQjeo
Xv1gcf9NX45bcWt9jB6iX2dWpLI/AtSW6xUg9B4FcHB6b/hqAiiamqT/4hq9Uirn+4aY1qrmGndL
jtce9n2Y6yUQwEaKCckJTnBsJWvaL4VeZ1rM6W+A0dUKsbhLuBM/KiQ6USv2QKThd9eRYh9EP3Pd
ipFE/EkOv2aiG++hiW0YYrPcY789qI+JyejwykgXFsM+Nfhmei0iDZGzoKSDRhRwkHT8J3EwgqEU
piv7EMShdwEYdjMX50+QsU5fQxUluo2OxUmI9g8yr0XrX//ByDAD4B9/WXo1bhOJbgS+R4NLi44X
dSj6qnnwfaJVpE/S18Qtq1RyM7/yMJ2g/hzW1h9PCrno6Hh+W85vl8ScydCb5WjYtkhPeDWQVZOL
DFLnX18XrGcipqhCHlnf5CWUKfYJSv36mLDts1oGHhKZgh+xyxubYbcyM+21HyLOri3TqFtTFSQX
Lo3+XL4vdlLupMOll2GivbLHLQgIxM5z8tO7hmfzJCHmqxDPjRWBkbeWu6AeoXIw0oTaeerLqVdV
qcE/1akT+8WN3paNop/wh6bfz6C2gj3pq7qhBjI4njo7NCJ0MxR/9fW1zO5LjTVORyw9bOR7AoUV
+kz632P9W9apGwTp7S2WgC2HS4qXBfZp6MHscupwZtSSeYM8UBXIk/lWc6SA9cCK0S8bUrUUJUWI
fhn0AX9ZC/OUO8IR2nd1g7XQOZSM4bqapjBqT97ZJPcoAu6KnNQzxlnBRxEgyLo6xAh+tdhA8X6U
HqAZ+d1+y/fedywLaY1XcPHfv5dLVDp67yhDHTopnTXVpvdxHCuo/tfJdhQ/JNY4kq+Ognwb/BK+
OSGAGazC4oEmmc/4D2EQ4tevXJ6AGDW1lczPEhdR7yvwwS4oh0MH7IeujJbLcn/CXVzo1/yRqNqQ
07Fo6Yxn6Qdhzn1DgWq7EOiXcJZALCSEVAOSpAYBqITGuRtjMkMkrohQxL8aH8cyB+TkDf9zKE8n
W34+8U5v+6+EFv/26Lc5JWjio71BZ641ttsh13J0N7jC3Oil2bTu8YJyrSkxT7QEBvLJLEG3Fx2w
XLdFnBfcOeZn2MpGC7wBK/gXTYyvUnm3gU8P1riqPKN3eAVUDBBNrfecuTIY5KEGCkBXSgOMyp74
sRAtbhdCG8PsAvGE76tGBU1JoygKyJHvdf2JEqbIeZTEQsLNCI2wCg3HezU8T6LM4kCF6HX+BTod
iItnM9pdz/sslwl1fOwwl4mCgYPRJ3Gb9kKa/48It5A6hw8eRrn9nPBVHMFN9ZEK84ndOMKX1PzX
LcCGl17R3uEjSAnoxR7Mc9pNnj8vt4vpkuUsq8pTErdFVHbIyNSjOh6s77OPe4viyv8OEmvxM2Vh
L2KAqCcGAuTtBYUjoTo5fHldhZEcESp8ujFpwf60uXD1LlZmzJPW4JKZPZwU07QrTJWVD5WdH0ZI
jI/02ivmJImeSImy9Z6i1Wzww3cCAdT/kic8LKQbdIEbKFxIaTtiJ+PMMCZCyxxE5TiB3G1k5nDg
oNAoqFMNC5/jldy/iKAWJtbwERR3dmRcs2shOY9RsRMkHt76feUEVOZgR8bzOSWPuYwdcYUkuZGY
fgFTjDoRJDX0fyOivXRG1U0hWOHbTxFqFjgK4isJ9/s9dkJVGUDBy138D6TEGBLiCcAKKbHRNa7J
sQEIh2NQoJkeEm49mL2719OrEndQ476sYswyW5OKwKC3CtEG8PvfRYzLHVFR0eo7r/HAfYP4ADmM
ukTmjr1EFS/lOfGBbuUKQrc/VTj3Z47HXzlJ1ocZtgJ4FIzNeQ8CgN2ATQ+9CpFbgkj0X6iVLbMj
uIHnajpPPjI/n/hUvT1Mb0x9QZm9IjgblGac6WY/BMhlHWFWhH1IYS39/Nnoe8mAB/7hVf0H//bV
6JafwWl2yorgo/nJjJkjBrqXREgwA26z+yhPcbrjwBRVZ0gE/RSmDjzOO9r8aDUXCZ7qmHQM2xHM
oAPS9JMOOEmqb+JqohV9BwOn0ZEzgxauYyvGmTXNOkMuqjxp9gpJvoCcBuVIkstMxujXPfOzdnGt
uXhP/tok423bLIxJCCmfQaemklVOEzTHBI1UAjRattkLHkhTpBqNWUqP3h8kwJ7o90vFSIa/oQG+
lFgXIFyFvzevbipUZHf6kMRc3kIP+cMqrL6WNSsKRC5pOv8cMX/aXPBzut4s8snAKDEQNDkaM64X
bXfSC4dYNfiNXO4SgASill/IX2n7OLpXiai0yxPNhhZTgsR/hEqGDhUpfIc8FoDw5jKIpqd5KFyt
Y1glTKYy+UmfNU78YWDzAr5QTr00rUlAvixbissLgwquBgDujfJT1rwlLxpQFfObWvS2YKgYgmg1
YL+yRah1vFsFDUdfzq2rtZCzg71Lwn5o0CxQhe5Edymcvs6zz3YvxLqe/ZO/Vovo1gNMoixWThd4
+fvnrYW3q+RWD5GMLNKcIWat5o9LyHIS9EDbOj1/RcdUDRPGRk5NlDIt+txCI9Oj/YitBTb4zS3H
9/BUCKLgIKNEGaSjOvw4LUg8XwmjIWyn28wpOrYUq4003PAirTr4AJpAgsZANfBzi0UU8TwtEvaS
iyFNUf4F712F8/Z9l+CAj5C8o1slg30agfihxVrA2x2iIiFyIFaRpJpoCiLmrAnTnfzdVumR09iN
+LqFShW/BX3rW+S6VpHnRalmfVdyNwTaWk8lzgPxZno++5cEZArTiBIxi9zoCB3gelCFTU4pHteO
2YcSzQaDYztmJrfcH6muB1wR3fuq1ViW60RZER7Ae7dWUhc7iXk3ogkKdHczcK377MrIV7KoS7s6
MsVBFpFw3rz84VJhaqDMqHpmZyFtLu6Uo/GQckBhxBQd4rcVk1OV7yb1ZDtN44GrKulOolS9xlpx
CB+d5hLYiyxKUWPyfv3Yws5HZ0hCZX0McIrJcMgDQ/fbzWNvD3a/WU7l0304XENtwI7GY+qVCqZT
9j/m1vKp05A0jwQlixAcqVJkCZZSG0YdKRjl+RHZxCJoPKipMgB2jeSG7hUBeSTPH0yigs8Azxo+
nPtnALchMEAe5OlqdRlAdrqapA7+5OfvxOOPtFSLn86iAuRnkriD29aIAEYY1ak932EVnwLtox5m
80PIlkk5Yd0A9DjZs1lxSMJ+sYFKKPclcYFaLSyHkOgL4/ZDbEX+TAso1AbzrTfzI+aE2P4873Dc
pZ+Khi7jDyDlFn3geXmFY/4S9L0qhWarJcGIroPNwbWuk/0agWNOuABc4dCr4FFppw3efDEiZNzV
3jy453L8xd2xwFAQ76lgyYmd3aDFdpKdS9pU3Ha6i/tNaP4I/P7jU4FePDwE3KcpQfpNeGPkEx5W
HKazjTz8K/VVr9l9tWW87sBuDqNmClqLntyF5BazZqzdgTB3dV9Yn9Fgd5vXV41UkDa2w3nQba2P
p501WpPugMQ1Gj/FmS0QgCWwnYPuJ4ce1t0ZxWBEuveSPm8P4xpLUgblENQfslCZNhS+BkteZcUb
Gk43eK7cMgDzVjB4RuI00i3b4FaD5k1ZFS2FwMedD5WcitNDjs7k30YtwyN+NvHy3NHVoTXBDcmi
18WLGqWmpovBhV3UbQOZ8Bu28SW1MZ72le9/Ge5gfvRcFtg/59YDzMQQpJ3dAEh7tSu2p50TrmrZ
n5lg51cSsHP4ehYVq4z0igoOHefhsPlKCkOoCf7Tol4emU13BduFYzYa3XFLl1+w3yIc5NhWeYD2
jpD9zQEt8Vi4w8ZtSFuRgKbggv7dPWZRd9kzuAYUb7NKW0a5GYQYb7PpVV/jEn7Uq40g5AYWCMWG
iHr7mkNwTDZ6axPswUOub9vcgQ8upd61h+YyGKODrEQfsHFE2xcgSDz9OkXg0k530NRiO0QkrmpR
4ccAmATYKP2N1Iu+b8inaspIHMIYamUei+W1ap5nQJMWzJEvUD4SJTppidBSmTMkGDamUjCJ173y
7BQc0yQjEfHsmtRCkMsxj0QWGbRu6kiI9lhlkW1cpBwfMA+n1Zy6QWf7IV3qDWBmjbFVjFmf2xte
BGSc2GwFu4AhRJhh3HdkKTMldcogqkQ7Asj1Q4EQR3N3B1ef4C0fT1r21XvxpxZ/KLhf4UJnaLUx
dp+5Nlsx2HiRlKN9RLQl0qiT3X7tuhDlZnMut/WRWX2MmiqscTAM56652HCFAr82pEviFYNLVpyL
amG2VHfeJvsFPSee8Yyi2sHEegkFrqhGnBEUO2315bXRuDiwQIwXjZsE+YxDAD16cIcASSeuq0vW
TEidr55y+wMimqxh6WnKRbF1gep8RfRzOJHUeaiN0N0He90nqfSwbXPuL+oWyJ0LDtcFK9Enw8wx
5UPuCXonFeohrNTfQN9CZYSdg6J1u9GqwBm5tBrOYFb9q1qLpjSaS/nUCwvmBCRoYcqdFmj0I4mL
iu8D6gl66HlO1aVPvHmGTN4GfpJV/bTwpC4vI+QKtn6G/aozBYi/L9+q+2UfycQRyPvXHs+6Siyx
/GXAUvCvZBit1K7vdNjizqn+7T9R5CV4QgMu0KZi4gH9nGVdW+Ol5+xenlVW7+9TovxkmWBEHOV2
sdr35foph9/xUJmCYXfCZz2a+aBS0rbCz7AmbVQ4Pxr/v8Iub6AwzLwEYfwplASxO5PzDdYKNLpZ
otQ++iAHJ0ITSKeScJppuXDhggDa8BBry19T0z1yB9iL2Zl2z3u0C/zhhtu+UZO6IZGUPg+Plsgn
zla/XK8D2e54D2SSg7f65Q98q7wjiGZOhv+cPNXU7EYS+qcfg/JrhILF1qtWzdL0o0JSCNoeBOq3
RguBmiDLo4bFKypGGNK14MmJOQaJ8uNo3QYzcY4gi6gtECwAHXXKI+WbNAKfnpNQk7TYZf3BQV+C
0nm6j7zzqhe3AKTzgADzdbBcS0lAxEIICYqNGJ8G70GaU/JINhJZdHddkchf1a4rVw3s4MOlq4q0
BUboOEed1Lc1Qn2cytLVXvN7yN5ZBtmHflDipYXm0uhi/quVi61h/BggjKXOeJSFHVt+kq8f13lX
hCeSnFP6H7xgdbvcfjD0oxNKplH38p+TY/oQIHndvLjX0YzjIzl2of89XFGWo4s1abkYzmmFoqO/
zFTrt1GR/Cy4uzN47YPU8xIeUD2aC0DZuCrtR9eyjpcQULpodMyH3/Jm89jl6pxiCogTrs/lKZ+m
lqSNyj7eKSH91paMEc7e2FbGiG09uNmpXlJ3jWShxy+GnGVRLWkqHXltRp8+A85kf076S/knLEQa
m8U/JA1YBZTIXYaVPGj/C4pH7EtJubtVb/cIYjzVyHI9E2hbX2ZcYpQB/j/y+UnxMOpiBasF0SLv
tKM5h+5SCUdnL8/kLsTdNQfnyBAueXGY8PLhPPPiCq7lvrXg9dZcy5AronspixkttKFVWHBjZLqa
njszlcnbPECZdAAW6j50vXP7fgpz1oLXOzyl5h53yP81/0kBMPElXPBbirk50gJ9p+3qN7R0NdKb
63omIwfB0P/5tMKczA5ij3/4dr1eFb+HSAifVl/2tu0ZMdmA4yEc5jPJcMMcI9aPNnbsa5JXFETg
I0uTw64JEMjoB2HGo7Ol8/BTQEXQIBIYlvMngw3Qu8JHq0EdkfA2pp+YLRwyIu7I//rd2Crd6qpF
i+ghcqgwbG+gmNrPo5SBL8oLTIZXEvXN183aI027LSqJVuTcEGbcxOEpFKJl/gpdlux5+UF5EB4/
3un49PZwePwHMJkhYLbg4WzBxfMebtbCrD1S2wQkR4xZfiIYR1hpyoQeGOUPC5D9hMIoLfyrXpsG
qI0quOs0H77GT+kLzGRRnjCUUpI8pHdZfG1h8Gk0wtIrUU9btNhqIjDxpd5wrdTXOi4VVZvUGF2r
zOnQm1m6/HtsBARnEi9hAZUkxkEO30axWmGhiIgUjt65gKdu+eB0K7iPvgzSiycSdLssPkn8gf4E
mcbeOy5g2RHsG9fCO0VsEJMJHcj7/TUNImreLHY5WLuK0+GtN/UuSIG10qpBME+omt6SoqzSo3dN
bZFI0zSvXPL2Vy1sbEqPrFl+5dUz0IN2x1E/b7s/HsQTc4asOg7D5J7uNbg/3Qfl9B5XrIMXT7Za
rl08b7h2uthvmRVR0V7FR06Z8R9mHXo284bYbBdwUMBZ1ltdivGNnOkypssZ69dR8mewvl1vz7Yj
XTm+ZwJ51mrC0Z1P+Ki7bvRQSi+SftuuEWeOhZU+mljUbn+NgxLlStrz3h7YsbgPgbE4WJ3J0uX7
85tZ5kUfMcn3J6YeDWKUi1/uIOcWKYf0xIPjmQjVnedc77nCJjKHujoukB53SmTnYwzlLFXirjE/
vDErNFVQ6/yQAbSaCtQSHFmZkwMXn26CInfyUgQHHtSt7IeU/whmy4eYuBGXagsDSmG3XctgK5IQ
PUSUKFVg/g23YaBpCW8fE4zjJPBHolo7PlspeIGKApPyQmGYLjsXvomYI3lZv1Oi4O7ZP7iOHCn3
+V+fmdCxQEYutt7vQN1dOH3qGLTcE2Uh7BhzTOl1uuj7tXpfqFjTgYOv0x+ZL59Gs5AMLMwMWcK0
caMsVKJ08kPthS6VqgTn0jJuj0hGbCAb9P0fasxfejTP6uaP1PbMV2kRJwQKPDk+b9P5m5IzT8yd
Lwbm9AL6XTmFeBETUnnJeqXJxndm2SISYZjUbaMClUQIfE3c8ydzfeG92DkG3tPWi0RhTYDF94em
nQh8p2563Nq/eoecDCe/mBWBNy2q2nVHXI/p4ZBJ5YR0q+NU4aai05aC+ORnnF8GBxXupkOxl2tl
P+w4+wUSrVDE+fIEE4wVFyK1Fbh5Ito/zte/d2Yv3pFOwEp5stI1m9RGcvQEQX5LEAzeb1IYUQNY
qTlDHLlyW8y6909pxtHB9tDxwPlz29mMDIqsOeVnpYAj4vVwUx3iZC0fAbC+eGH2gORT81E9nz27
IRctl7yQ81w5xBlb8xEAp+cIWy6Gv+84NTAYJkvLtAEqgjFTK+WbULdwzC3oP+M3gzeNzRFAHnM5
2i3+8SWlj8K08UL6Jnr7yuznhmDRISjCHIT716JtOOAkALh+/YOAYCFwR1JZfBGwtoAR0yO6pGEn
lFNNMgHxamjYHIk3PNIWLaWpmeWb60MIRd1QWvFdikAOH09Oq9aD7tbZpZ8HQi4GrGcfQZ6J995Z
k/+qTTxuXj4ww+2hz07Nwuom7bfG8ioNKpmsHlqVvFkzjy9913O66HE3C2m+Rr326hRJAex4Fh6H
mdxUtU8TNOEb5FbffCAEwPIk9iud9TVBJ3wOK9tQdZSV5IBpb1qR9bfYMcX3IGj74bV3KttXDRTU
3Extc9fuMy7/Tq9O8Uxl//ygt56U77MuW4hBr+FfVpt8VQZHNe2jYFyRT3pEFovHONmQF2X3Uix5
AIRpPaiBjLak8I/09Noxn8NVZD9YIGeLWYsEWvac0NaGcMKoxipHq0+isaioP3As0/hS4EuZ+/2B
YGhhrOCw3Lz8j+LaqDPg4FZND9zpamF3mCdOaSGnLOuNI214sEiSBhl25hrGm701K/587BuVFysE
+TYZ4mhrsEfA8HhtqBy0gowfHW8UC+Yua+MTHJHifDD878v/2mekMfqK5dpJvb5B6dbbgIKcgxdW
bqwBWPv/SJV+oqVBOeKBZnNpmQOrJ/2w4Ro+imLQQt1xWADTS9a1x8oHBnCe2vh/S8lzt4zUVR9V
06SlpyM/5oO+RoNT/xe3VAnw+ZudhcCg6dHd7Hdx4QYhwMeEnts03fwBD8J4E7Q8fR103uORadcX
0s77ShFJc9S/Ip+1RxWqSihXrfCHXb7U86nBmr22h6JBNiJCLaLtXYyR0fS667BoQ4nj/6lTe03T
lsGDftj/euafBapjCMuPdfiBrLOA0p9Lqa7rqj8jO4AsPJerL2ypOAeqEm5wn5oY/xaD7dvtfBNs
59/yugjm6Ny90Z6/VsVhpT9d420CgFuCf9H3B1pZ6zayxidQpw84S9bGPTLCOk77gGJxTkROzxSI
e/Z55xm4HRTewrOSB1S2IGXVPMuUcy+AvsW7LBkWbyJXcwWxes3UyfCrksgz9nA+uhXYByiPZ2fm
9WmyoBVUfxxBdW5MJWbL9+jeGfuzKadd9Z4+PT+YakTK0AoTMoXKUw8xJ2h2HyTD6KnqcgL/vhFJ
txr5bkIqAAbUicCNM7e2Tjky9Zu3qEJSAJ59IQ6M2XP1shoYZntnOIACxqZlID1nP/Q12uPuYm+V
1Ccp9cEdY83HiA9CdIHhipiPD0GGCOmXVhOu93cxm3AnFWojbgPyk5MMQFtV0DaxSyBE460j9Hoh
EgfFrsPy2ImjgLl9HpS68shwDH6MlXizUtceXfYzv8AOOGlaUF6w2GBaHMIDxxaBZz8Rf+g1ZtsO
gLfVdsYV+wyRl6PeKnDzZjNpuqDjz3/UE+8nNScsjmtwDixyquFntkthpbqpf0xITaVJiWPLA/WB
OW6fxKgVgJ9ZS8NHYHV71mUm57DMPahw5N7TIB0WCJ7EzvUUj68hK0TVnhNgikQpCbJ10p+KDy1u
NuFs3H6LJ4x0Eg+Vb9HfbpmmWdq7B3OA6ZmoVHFCSV/T1S/fmT7szAldE3B62MUwXC+sgO0qveoY
GQGEdmdaJ5tMekoPw2OO/E4owIY5U0ZMrl3kSgX4lwTcSZ9iSwNFgHwfUfUURKMueuydTW2SQqAT
HrKNrjwicQ4paoeFTb1mGBIdn8Z9g2AeLhP8MR32RswZmeEoAbz8iXzRyzmyiz73YKSc5SRMR0Fu
s5ium5puny/e0gwp8r4cvRUv4+VmpGC72eIU0gF6tE0gjXB2qxjc7Z4yThGR+qI3p7B1RFCZRpSS
mAdowaLOL0evSVEnvDC3TpTz7hov1s2WufKjp0USH31mwh+v+iaUDV2MThO0y/bj+bSP4fdIaxEH
3X4y7GbhbP42FS1ynm1dkeA64Ykmqu0DqcAV9TU9bE6ggwOStj8QU6j+GJ7iSEQ4eto+A11HtIZ5
RkWj7XTNbPUOmdt3aPdwXsQNJCauSPpRvNrILO1uUHLtRnWRnw/Pxgvz9Ag1d3HK9YjgCCWeouwS
uAzQeqQAJR9ID/BAM8PpqjHk3Re7guA39+y9cXqznLnlfuG+BEOd5fpHENuQeF6L/DxUgytqEDAM
usyx+Lv0GjCzpIq0W6g82UuNwa0onLGELG5l17JmNGisgqYi1ZKDYxHMclWHVza+RIxR3K9pYK3l
JiWC45TZxojLDRSUJhupxNmir2O8+PR44IpcItqzDYf3I6jEzRUZoTI+TNzlCCbY6tjwnO+RfidV
r1kEaoaApfEAZkMw9Zdp/18kw8kFBZSGGlGA/go/o0PJEaV23Uj7rBq9jvcGh3JzHJxLOC9Hf3TG
+UbJ0v0U02fm4viJp2M0YzKePLDdWXUmwe4t2CJwzQY6+0+vu2kA8hyJtF04wHQ5gAZVCSX/qUkT
jMb69siygR7QBphuS+umLxI1JBHIE7bSTj6zdRNKv5o7Jo6uCkWt5AYwoXfuUNFlaVA63ggArxUv
in6vGgGGn/mzLAPANonD6FLgYHIfET0mKI5JDYbJybLBWIlChP5D2/5RIY7UM8R02K4ghoYN8Nsw
oRC7BIJsDvrwsy6nm/oQEG6bhtabpQJtRYc62WFdPGQnXUlElbOQ9NF9hJvvoPJHkD8g0zpZxshe
cZkq4KCQ0tKOhINcHjxlMbPCAGvPxTLDBr82w9lYLIUJXOQwV+I2ur8NDfw9Rtw3xwb+ils4T9ec
tWCOdt4L6Pk+f1SxyAIWzhIvuppvesjWCUxRuZNKIJ5AJCqcIgZ0+8Xdid+XHIkZOsYtnKcXk/EK
QLubOuyyv6GebuMOwaRN1vFuBMIGNkYGYk32U+vYB5moiVx7/eW9gNhzhye7KZZfDTE6Y+fQRUzS
I0LykttLnmsDqn2vM1v6VzDuAiKTh5zHfTJ2w9zjQjkxDAEFVh3thMGTp5Kk2SlQrj5PRx/y+WJd
AvIf6Voj7wrKvArQQaSaWW4hdIIXRYU4QjY+sC5+zInojemEP62YNzQ6ftr4wQMAraLYj9sjY/pu
r4x8TGL30xtpdaZqOG5SYm1oeOdQTkc5TPnvV6MElDGX0O/erttEHRIwseCZQdXdtOSQgjQnzGfN
6ZZsbHJQIbcp22baNvfaoHoEVj12gBgdC+pTRAQuO7nvd1oFj5m4MpCzX+BKWkENKsAvva3oYwKF
JbbS2LDkj5iPjOeaCzYCWnyPucYDZjyzSKn1sXSVCtFMi9BRbu8744bHRXjPkir5JgRwGh+Ipf4x
4fQvwPC//XfWXY1uUYrwQIu/r8XwNssWy7vzpJfJdipTprMyqcCdSeEv8v+wuZxM9wH1Z8XQ+Eux
qljlu0FkpFtbSrVPYhhzAdjSgdvyCmiCyS0z33aX1PxM8OKki9D6H38QJtL9DAA7n6B2FdzjnyaK
h1iRUaCLbD/6mAuZX5Y32R9TMrK6ktdTWkGob/xL7TW4E7fgH9JpxKaisYaXVqDQmrXqhm5SGQLI
npAqo+uiLwJ2EAH3W3aZDrX5rSpBhElFywcA1GTiNes3fi/w1+zA4ANmibGWu3EBamtmWRW2KFLj
KI9CTD4gAvwh/xU6xQXgCbh2N8Q4ZP7H1qecOwoc4K1M2SKQnw7H0oBtkkR0wSUfgZ00VX7K8KPG
4/UvbbkQmZaQjPoCZ+UGWrSaBy32GnbzlLHK8WbvzilHwmqvhLipGduhUAgkKQv5d2jzP7Z/8APB
OZZeN9t4b+b9BfeDwBOz+qg+nB/uJgkbApnAKk8mFnyP2xzIX1ELVoCR6CUIXHXu+rh3l2MoOJqo
F1RJtgt9XVQYRCKSNgBeZ/ZizxyQTGnqRtpfC7XiXnPIpE1v5A5Vi0xaUDUqnuEErWhrSZCQTSMU
6MOijSOOzIE8a8wYh6bQZBSRk0uyGWVQPHrxjWFfCrxRavoOHO4876SJJyZsrLJKjss3YQ9pr1LP
Iow0+5DZJkhY5xW63fhI7ea4W/QQWXbjZLkNhsxfYGQG78qePcvfO9qPnAdg6xpH7P7fG0WVCxey
T4iu9O5ZzmlGwv2Ty9SipyRyI2DngdOk7i0kuEmBPsstTCsX4ysiKVAbJkgAG9rlC/nZEVF3supW
UoTKvmDH2OdMTkGcNV+xApsICs+gqgGEcMIoKrPmpdXESVm6RIDKCuSUDh3SvKc/SG0gyhxbMwp1
mQ4CkGRy9HS4PE2jHA5T1az0EEvbXqITgoT/zx+vsXE10Yu84FO6wuzJkzQm2syNG+7XqZs1fcrw
LJP9RXv5lXlua7fxCioxU4rLhiro3NYONL1R4dlXsJZqlCkmsNK7VtSltPaQ+wyCogkkHFrf9uuu
rvKAN/J/rFT9UI/jG8HSyCOth5SqPjilqbBax1Q/LOxzZiNbnZo7WmwExoPAFkwF3safjL3kIWaO
EqDciotW8i6McAir+9dlfC2gdvzkgfReIm5mvfmltR8pynd8jSu+0RLOWBOLa7kJ5HurYk5FRz5N
bxE4n3vuSkUH/GnYSOfEO5nK5HXYI/lh1i/5ZzmLQFawpGmR8sPJZ67qBPdxUY7kx9ZesEqx5vuw
z3VvDH4pDOO/TPi3bNqtffYSfNI1PYDFJUVMG36JTd10mdF3xQbJry7l6yZbytODGfnRSe+Hz1b5
zYkJXicGDZI1etOc4ylDhc84E/brpHeAMUN/wwnAnk6TeRu+LvmMb54AznsUB53BoI1onBpkZBck
qhYqB9GEak3aodQL+jM/fBADsychZZujH+h4Sog5ZKZ/spKkWFyRjNQ+Z/E7sr/U0K0dYvZfqRbN
0kqK8HHm8hJGvS1ewwNlPsJkwRv8y5f/g6r5fvp/+JrROdTibVEOmWpljXbnZrc2Y4BjUA0acrDT
6vx4hSDMQzRJlj7gFIz/TH7pmnS+/UBNzvRu5/CJ8aEUE9IyK/h86lJAMSGBAZ9J3iVlji6K7XfH
g4IpFA7tLvKUAlnZlfm9qaTSx6h2Pl2HLemDwt/OupE2U19LYu0ILUGZrKUGpFUAxfnVtb9JCFeO
69u3lYAXBKRSHg6z4nFuwymu0oA/XqYqxR+kJgeRcVf0JOpwn875aley8PFNr3/cNHjCzDsXtfuw
qIBlY1j7YYxDZWe3swXzeFx+X72JtEO3KgPThGZl/At5U5J1h9PoqBkzdN5QsMtuSCHs+fOppY8j
NdRHMxuvxGxocFRuznacoaMQD5WUu3hvvyEVSFIits9Av64dJ8zam+jXhPt+4Zy3ZFjgYr7u8P7U
gz3IL1S3huDoGRyDAV0iqRK+llUZJhA02bKmQdDLIf5f9oYt+xtG+7Gi592pqJBWjVWMq/QOrf1f
Y34dWDnykEfX+S0HNVkjazzKA4Iz1vDFcpPY4lZ6ERhdwbJrJjmv+W/wXGWIO7uEzHL8mUsOEkye
4qtj89YOal8KzbF6HkrjdZxKyNIL/r5yJQnyou7Yl5QloBQEnFUORFZsJdyKUPgb8oxfHkHqfhWK
vwigCYDKa4xd67JH1/CifvrpPYOwNn3ZJy79rq4CXHX0t0enNUEvkX5r8NEOpg/NehS//P08ZpMv
h3naNLIAmIErsjomx4CN5xkyleHsiM2u+TKNELqVe0dgWsGGR3a62Dvx9l7L6Ejb5ASuFICsdvBu
4docyf6h3Pn85G9qnGz30EArxUUbOmgnkort2c+63eaIN0Doc8v/w41x6U3ojCC3lBW3ZUwWvrph
C99rUQnd2r+eJ696y5/eyhzNNnyXGdNrJo7Dn7APZZLKYY8fEMdvb46h6Z3sGGPT1gfBU+jaqzlJ
+vBMi0YMhGw28CGJLkJTGxnOT9szHbDdSmmw0TuSRmY8Bvy0b0G54EC4l2cnf2rZGgcASjGOUzJq
SPtqjkXiFlt3pnCKnYUpbiQapkMg/2252dUbqfvkKZLrg933Nuh4F7USK3SfE3Sid5rP64hUoXVi
mybcoj7kbL0r8OcRRxI85QtYy9hVAKVmUTMjvIzY38k/33i06IqBd3dXe/XI/aTN46x22/+kJIAO
EJ2HZp1S/eKfiogvOkjw1iCq9kYiiDVPcHYgdNiZtDUUDFMXtCh769zD5esZHpJb2StmCAiEKS65
wi5/RsFoQHXDdfcQLkhXz9JL4nh6UwcX6NErVuYaspuDRHRMlsVXzBRZBnxc2RGFrqsRyNaZfkk7
QI/DPOtyabhTE1ZQIchM/fIoOZ11y4cPW0J/d5LrNYNulbMUEEnhHTaxGjOYIQyrijMemFMHMV02
tSssH2NMnyrbMDwQ/WcVD/84YprrktIJ6ut4B23vjfrJ03kWpk9Kg+IOJFT8oGMEh34UBCo60uwc
AuzDfaqlDna0uGnyp1dz1hOst5LncYNIpo4Vp5p7Ourda+MyiTqW/DRlXxGZ/8kS2v6cX7lxocjc
0M9MfC1IXCwRjPnu/MgLzfWzd8zLVxZ7anD8pK0EmF5ebfTTVrhsn6DWiiW7GV5R4CjJ7khumCqT
CmG/oBUrIB5YT7CxGJWcjbauTR0NltMfwXVHQ9yBrBJTbOgJJq68SXqhsMpOhn4w6QY0+e3XCVp9
1bhwaXTpLGSEYy4rP3in8/KYSyhJIMCYz6bRY4jBRJa05Z1/9QgMJQ52vvIvFA2THXVrqOkQKmpZ
0CboDsANVWLAaRfBFUZEReHX/hPO33zVW5XSR4yOLlneZaV03qJjLB5veDOXgFeOuawUG5uqXJhw
UFNM+WFDAhjAdh3kqbsY8CW+5i+z+9ugSZ7CfqLoVc5RhhG+4R8EaxBvL2A3zOETuqwz76aygiyp
kuSgkNPxZ9gU9nBsesWeyaRyF8KXtySQyTuU6/o/PIDK5WrHJMXmW45JWoYLa3sGU3WtuFVNKDk+
FI+5Pm3ubLHHWvX9e4NbRoBXo4+ntIDBdVl665qb64DJyUWIQOsoXyrUsCb0yR4TIlp70K/pvve/
xpZFopJD+Fzqd3zubYhcolQqlBHgSIZTBfJzVaoo9P01V+V99IdseizxhDOcz4iYmFc5A61jfMmy
QETfL3qtnpy5SGyK6RqNSbgUUsSIuwLwtVeYA1Nd5QwtzDNa98fTMg8svfm8Jz80wAjeghPRiW9R
v8pjMZg2nZMA2qn0xPnOMHgdxzN1eAbwfnImog00kbwS0RmXfDBbuGAi3ILA36tGxkjKKbnaW+ow
NdiWMfSn5sNrhDynZnIbpp8q9qFyvcRzy4WZordW8cGt+pt95vCGmXZ836s5zaQGPPUqwCcHnBuW
2GD3plpCuPG717XhZjPwFTOYAtAsh1RAez/HjliVOQeR2pvNG+WekmnWoosxmSV8v64sCUGPcESj
KXkBKlHtLhA+USlWhyKAc6UPZ3FoaXyJHJj3g83nbT0y2B9vaqUN+knyJbn2hcZncmFrQaPosIQ1
1FrWTknyAL34zSegCj3IfCOj9qaBdUZrLzTGVmTOgkWTC/MBIcjzANg5ZB/XMi0vw6X//QSKOf3L
WsYX4IQViQmdHzcUeYd/cItBL2wEkQhBrnMY3vU7vZWqOTKmsgwbNwAeUL83ie3WNJsX+DMRob2/
fPnohW/b+ggTgzZ4CfSJ6wqVq+WJeJE/NTjM1OgFKxjeOByPvacb81RpYvNyuVwtbRONttCjQnf4
1cVUlz8cjDmp7b47lBR/jTy/pKhvIb6jplU5D3Oj/jFzi+u8qGLkLHo31/rneHnlTWgG+UOFuIcj
pbQLqEuVrhO9gl/PpYaskND6420XV5KFHC0b6Q2alSSxpHVF34NeXTnqyfgfKTFaAiEx7M4+/SHm
AIhm2TKPxk0BlXeKRWK+K+SjTqmUbeXUntxZ4LEw6O2iTS9CPqGfs2Q+OmH1ebmmO1cG9bEa9hTC
nLqJbeoE1rwKO+y8QIcBm9YM8sZzyUH86NaHpamQ5dTQqYafCMmhF+8nGUW9dd2iJyHaVbJXkCfk
zU9khB8X0TbVF2gZKYBqnpOWQPTM7Bt7u/bxsZqr0qS0q8QS2LzLFO1PEgqIHk4pUq49oASnPCDE
Uwtkt4P2H58h/elfpcZFa/oK/bUX8oFJQNQudow4+pGvF2jgmym2gJ33t1CY4PhC+baZX198EZWU
ix3Fz91XrYSsj5RutU7TgRPeNmDt9BCL8By6QhzsClVw2kDg69vDL2AVKXWWUBmRDq95qFMESpON
kTthflV9Qs4Pbe8ZZepXrBnnzv/3FkKH1WFAtXfiR0JIH/V/vmvr2wmOSklD0eHNSLk9xJa/Bg7+
gORQjQi3HV7fLlQv8FMgYylwJCteeml4j/SG/izwPAkAUIIR0vIVRusOc+o88UXDgjmSxKYnFisK
XnLNBx1Us3HkguMPOiDi8Dq0K98hryFTGYzM91vp6HsliV3+Ox9+812ai/FFBhc3C1xz7vFg/ZwB
2F1cKSDYw8Xgw/b/TgLcKL1ofSCyR8fk21DXwTjh6eEkafGq/MKLbF5OGdei271WzReK8ZFDyaiE
J93IdWX26mdFPKJAqTrQivkRE0aoJFMs04UkIHbvIHaZtQSReefl9P5EETwOaUCAfdUr6NhJmQmp
E1EB2TvTST4racfqFeFhu60LzaDEMfusNLe1IBb4sJdG1hPP0n/Aarblodt6zdJxm0rvsmDp9pgC
EbzjQ7jPMEzcNx+J+BzsmOd+9l1eDZhv5ppAd1v8FQVEgOa/xMXM1V6DoHskI7G94u3rjEvh7RGO
+/rvfEywdIoMfmtpDx1loFYyFMYPbWpuVqlSUT76XhqghTYklUe4scMKLgCdNqVGXxTfvu8nkFcK
wWtf8BhBtKBdcQJPYdxlzpmuPRZtq6nQ5USnNq5LaruwxGa4s62RWo/EYXMg0eOsWAuVWDOtaiCF
GlF3RxKsOT2sNFiWY9lLuCU93dmCQKtBnDtxb2c4XZH88tdDR5ka+Dmjbbp+FmqPiqBOGXtnE7u7
/OQpES76bWaa0AgkfneBc56ibQ/kLD4PWIG+m6gJa8lBOIPbPWbWvsyHM0L1kBnGavkljA/1IU+u
HBgSQ6qoHci2TnX9BHq+xXUtFjUzN75l6R5TS5zGOifOUIRHwJjaYEujLorwXoELdMc22hu0k8O/
BbPQwntRUSKzKGXByJFEP5puaifW07E3S45tuVquuC+QC4pPd22n94uvSb2Njkq+xvApvE4C0eJy
2fnZRXx7vyTxxyV/j1rTL11YywpzfYVi5/fzWhYSrXTUglCU5I75mONobBZhGZcS6rqLmd0gJnI3
+DHPUz3HunNfxvxqGJ3Tmy6OQmKTxwAKQ40cZXMgUxqAxU+vR5XSamw/+Ho1m6k8G3pn75dkjWJI
wuRAAORTWj2mqEJ464ADZ9wbsCkdKMvSobb3uHMqsblq21E0Ad1h4Sr/RqrmnTEiccAesLQgEYo0
4YJfEadPr/Xe3gS2rjgVkgpTlT/w40N6POMLTXebCky1MG8tw4NxxF+csyMnw/xXqZdSgyMAthLJ
zar7MtczvGj69tQuwAxYVVpHsfVchoPlu7OocL0n/EdlfOVEmaAq1bARhDUH83mAG6gA1gvo8tjw
d5pcb4z2sKEGESipYSRwLB4QAHmLp5f8hbH0l257qNTVGVK62L74EidHYs8/Mg05mxKwxUBa0f0E
eg0+c+juV1B+JHUfLPdhiFY2sGPfOAKZu+I+Jf5e0yURL4KA2sbzIkjS0ngOgj0orC1seJX/k/+0
gjNijQ+OSTG1+T//llgN/Mah+HSSiHOLIIQS9objnz73fXM/hVcYMj/n8rFOKItYSY6NznghxPfO
hKhfZs3g1fjN/YuYVkEvF4/ei/QMNywRnX9j4oLw+netKXPM/twIGKwtK7g8beFhezGQHnCozLTA
qGnOHZi/2fWDScGeqJuv3ZzgKGbX19/WeLk3q3bOt3+4AOIw8BrdRuY2QutRR1gcqgPY+bzm5f9Y
tA0syVoEONRNqCctm23oR2Pn33dy83bIEiPolAdlpIxdZ16OtpPqQuEuMv8vH+wd9zjg5BQrjmh1
m3NW8T3cFGYrwDHtTS9QT2Pp2QRl84wDPXFz9HdbzncV/KGn3q54zIX9v6TQFxrDkolGG+EK+uIE
V7GKk2oEKzOTTavXZ4Dkw2Eh0o/qe8RiqUYaHIdvOfpHxJFGvWijGVLyZos4dQBrJRwsJqpX60J2
X1D69yV9U35PpGvXkRsjhkJobntLznXCeBfE8Bnt8kZLI/V8ZM5NI1ArSOtDIkNtk/1gqjDDWMzl
++eCoG0xpk7e9nFQ7tBVzVLuqOnZU9Lnd8hGn7kIouvPLL2MNo+moBuIaf25E/QO9SOd3029S+jC
FOxQ+HQJUt3zMmy6brto6vnwEqd/UU7jvKvZD9BxkWKlZDCK0TXQaRCxPkerB6pu36WrEXi5J49Q
KaNycEhgG2m2TG3KLZhQb+irlpL9cHs0beoqGneED0CNU6U/zzJOHN+87h0hiGPN/d61+NsW5fdR
6QNOtBuxEDVp7mdBm0owXSjr6PWlApdXS8bNDYlqT5wS2CTHdxhP13vb61zxTOCsAuuKLvMWtsk1
b0g7fjnXy6GEHewd9nOSjNlFNjfl72vgHz4ZmpwNsdQOyJvJXLSbUB8RS3ql9d8bJYNnoMxXcMZq
zabxLKnWKwLIdE6VjfdbZjUFexMMd77ZESMHOCvXI3dMgNhOPGXFzFYRqWEyERv9p4UlyJ9BS3/H
g/k7uNMBsfLJ2MuF6Dwd2rYIkll4PVBO3d5yIoVlgySdyaZiHWkMxPKWi8ayx3X750mhDGZNop3U
Q3SuIa4DhS6YfEmYtj2ys70LQOTFABPxq8PUv98dEcaaHi8WkI38WPumNjThlGg+IKE8sfzlgEwG
Yj0QepsD8DlGoZM9JjOnfyOZsrRbA4rZPOOvFadvxU5j+9GhnIE9z9IE8rriJCGtjyz5WC2orw4L
aQVi5Njr5NCfbBjbuI6TAL1xIpAaACcJVHPkwb9cpBbrkgLwmmkWQADzJMTXGSA3w130wWhQWKdY
e/M810hUlUFyheEvf9T+MheCAD3WaXNRH6SDoljpL87J9VscC5l4StbSM3iy7yEHQu435+l7ZGH1
xHODuI+5bY0H2jHYAjJxeU6/Z/xoPKqiwR5KGDCjWaQk1N+JzTxLhxgXJCCFZau+wKUuGBNNcHJM
YnKt2yyJqLeAfbLH3LaXeu3VkHcuJTub6hTUNzdIRJqhTnSSrF4tefpm8ncAnr48bkd9o3bTXHhJ
Enxf8kkFgUdUc/vP67AfisTX2MjmCEG2xadzx8GY+cpZ6EmVW3OgLymDvMNqtxlLRDLm6IZCybQH
cCrMCaKs7LkTQEKLf1viiudPQiRlcG6JoFdHaSLq62HlmaDPx6X31LzmwNtnb5MGE89PeK/wWWxB
6+bm+UFotX62+acE8K8JCV2pIEgpsuUSoKy3Qqcs4lDBzMlwp08eQpjaOQBMYRr4xUSwaJVN5r02
odZVVGIgg3Zea0YKhELDhpIAa+Nuf+z3ipNTJgubGf+xHhgCXElVhqkqeu1rrUB3ac4DUJuen+Hq
RXJv7pojebqXzHHrmTfQN0wu6pFiae6nZc/lGdvPsrjLto8Mg4K9VpJGEIeOnA5xbQkUWQAGBFrz
/w4BAb0TncqUaqud5hgXF4qN+z/kcD94UHwy2vYgPz/IqwYy4Vs3gQI+SbrwzsDyJKNxOCGs0Fkt
T9L9fD79iWJz8o3eR82Ms8dBWrCY/WkwyBIQhboJwBt83vcot4+W2YqQnvFD0ZbvwOurHHBfQnV6
cXzLVNyua7C4jhq5dDyapBIHyLhEqEde9oMbZ3fh9gghPaFFn/lL63tuRmhpiuAfV1kZai9++Z9T
Q7g/8pslQDdqlkI8bM0/+zvOoTiMN20A6NMPF/7fMNKe2zS7s9fpPNBAaKdUcVVA+dS3P2Wv9qQp
f4cBX8rA8oehnl15nub9C7RmdQJ+lwwg3C8tpVJoLZFUEfc8gvZOvLEYJvc7SW4wosZtStuCJYhl
ocqeAHnZnDP4tb0SN82sejCgaaqnj2ICeFuW+kNCnfWp66CvmmAqlY3xyutnzV050uMG/W9O9ZnV
JcOXzRUvP167Xou5k922DxBjJIgZQHKoo3pMQNLs7BfTShqoFAjYRHDcXcAUd+JPKj7GZZ75HY+1
IyEvi48PAVzp003BK1grQyiMkzywVPilUMzdNy2fKp2rLGcjRiLwD3uKqNP1B+LTsXyOdE6HkuJW
KBxDok+Ocp+xM9IN7cIAsoZf38i0jsVGfm9qbZ7iBQaHMklYmR3fEWlLtdiXGWXlo1wSI8fNVQu7
7nfKC5ObiUQk9IqBZOC0OwCaFvGpU96SJZFLHr6PFtjy/HxcppZUpcOr/Vm7ambduhwwiZJ462md
6UqQDiMRrbuRpJqCyKt3QZLP9W5exXOh5BV3Baz83KGx8o8U55nwLAKXUKXksPtwbiDvaH1gY+YQ
mAPVzxTdNatN5T4G9LR0c1vuV1FK6jrzTjkD95QVMtjuv89lkdSoxaSaPObFM+LqBISu/3upw1VY
4phMbblrKqxVS+S6mW7o0VSrMMELE7RXkJxdGkvNs7ZAWaujDiflZWab3tpl6NGxZ/VU0KRVBhCt
SMPPcLS1y608MRPBYm2oqHSdzryqVDuleju7qlslfyQoplDBYyF4QvAc3XoKDpVvCMjobrl+M0P4
23P1DWnBTxXJMlIkE72fkwtz1SdczNAmPD4FlxDhap0K+4lVbE7Al80//7oYqaLihbwppdMSLXvK
TOLqwojr5vR8T0KvaRA97GYRYkYb6UNYbJxK6nnCKV0At8aeEptLa2WTXD7JvLRL1k2zGJtvqjVd
ULIkFumKNqhWIZDn6lP3Gt1ABGsMBDAbCUa6DOmz47AbpUtIirvFfYfaS8Jyz09438RFz6NH6v65
PC8f9IRRgMGSeBUF8FnkNV2hi6zMfLy+lHBXNeNyp7b0Fv82mNsA1q/0843y6btIwAGyZLL2N7VM
5FjFqVtEKC4rlZ0q9CQnvP6iIwJnauZXgJwtuKAfLduEIxbZ80/TLeDwK3vx7FpldQitmeZAKZYH
srpzlMrJypwq1/SQB4I7P694Gl65n7LLAPWXv2BHjld2VJ/ntBtBI4kzx3X828b4xbcDyzk+rWyc
/1oBcbry2rEw+TEIaQooiWs1Ay5poE6WVUUGw8IuxL3Zd23toRSJItSqPtXCx+TOck9jAqRs8IyP
9KuGxb62UQzZe2g4BXp+7aK8LySah1/7X21OiyhA6tOVjHDKarkftNNmQpQDxZDShpspQ3TDkyMd
Dql4sXj6eke7wQxLXltYuUHR47v8r9NzTVNclb/dfrYQVoX++NpekD7EnYDnlACOasTNQCohzKQ1
w/CAdjWndkj+axlh2QBXEakataFq74ar4dLaaA0JNWv8bHMSaSuyh1zKSe/Vg4Tg5Fx/VHmyrWjn
NoIER4ySO3xsE6x+Ww3CD0DvUyjf5Nn3Ia1oT4Rhl662qi5+pes2RqGBaMc+ho6/IhsC1WlWo2nj
hq43aJwXh9N/hdwCCR91Ygz++z2jbjHuaMujZQ9n0+fIHbEFsIC9+sQ0t43m6mMq26a94RTxqO9S
7TFBTNRCcJB0x9kypFyi+xlX8dPQBfZwZkGiB4yyG+2CRA2vw6axKCOKJF89mfxx1ZM4sy5qVGdV
mjiJXc/0PnnJZZ1nBALzA2Q4Wihnd0p5+T2fMVkp+9okcqecakQXV9amyb3khD/eQ7cu8GRnZfLE
Z185QcmlPie5zK7L5LnSJxJQGJCf67x1uZcVFVtfdsoMvil81tmwyFk8Zhj1JRYhvcwiQMaN0XNj
s4R1boIp+2e/vpp6qgQzJlFLhz9zHPY6CNG1yLXu6l+WtbK7lKUbzCGRGcMcAa1Jh1QE0ZQO+NO4
QzxhkMY3IIG9JWqFAoMRyIkL2mVAQb4OtIhQ4ZVRdHakyr9sQPExQJqg3nu12c+9lYzgwYuQ5zGt
P8OdsEZT4SWPP+gIAlZunEwJgEoaVxMe/lqVlyh3qHtGlD6DUg32xGBiJODGPeybF+hJfwv4d37J
MzyThniC6FfsrjT4oVAgVfFgNfsNRJOH4P6m8eYVpevJESsDNI0aWIH6x6h7rGau7/rZ2wh4WtkZ
Q8695cC8g2dEGOU+LhkmnbEAXAlYLQ+jViHkPWmWj2ZRYrQhFEI26AsojtkE1XCjlSXdsFaA81nM
lMp9hkeztvgj4E+S2O092D2S/SQpoO7xwOGE9EfHuIfE1rSU9d179QwB9OASbZHSLZQOdn7tQcB/
uyRX8aCWdIe3mJmeQrqHPkXPGShcXb9KwGdoKOfH7NkU13meQqXVT+6NKExAXAcpqHkpsjRhBROd
z95BGLmt6+H+Fh9PUUEDkC90r7EB76SKHqYtmJLeF9K+eKwKnDqYcS5livwvHFOQVAN5/StKT3gS
054d5ALJ6453iyQo54TDQvNhfvS2yvKD7pDibhcp/6gq8mQtzr6l/YddQH1gj3707+TZKx2y/Pg6
sk8zIL9dGH+AT8hExbcSOLu6051Gb42OiADFnMj4ooERvO/s4l4t+ISae1zmMlchCFy8E8BJTuZR
H8RA/EQKJ8p86blAhUTI0NL5uUg/eEKE80oZJzQD2EX31Lo2CnuihgHWNoJ6Uhzj5j7cfxX0v6ae
7MT68Q4oWUDSQBhF33wxbPMwANIYz+SEVmGOFMBdiyw3C0Fk5qb2+kJlGli8mnJ0uP81d6n9oEfD
eAtxw5Eqd+SOJaOe27q2WS39S4KFxZ8orpW+UOJwWh3FeAYWyGS5mBezWTocfWOTv7I91qupum5/
OAfvzZsf5+4Hr4fg2V2Fo18mfg1XV0AQqn+97XAcsxuJwA+hzy7yN8ODJ4iWi2V+9lzRGd+I0pVJ
gPVZ4RdJiNCslLN+0LzyGUYwE6A7NXFHXk5tetAlebMFM5LPVwXkGmYuauUQDm4hTh9Ae4/LOFed
1yEBr/Q5Do6uJLkoYGaoinELrHXghEyl3/gZXctqOF2VLQT28hWYjKZvuVr704yRD+mkJVBL2TVH
OhKjfKURbakk+jh9WTn2FaxpFcBClC710W8ssE9pnZ8jDKFlUvC9yqJ/+6FJUku0tCzHOvBASLdr
AUehAhgzQe1d+EaxZlh327DcxmfKu6GL1A0sFz+MHtZ+M2y2g2KBTglUvKmWwwXy1SeX+1425d3m
BUVD81ICFVZ6FTpAHMZcGfB/AEv1TuNDEXTrzILkoAD5H/yoDpSyBylmb+kpR5AEORbgMF3HRnoU
Wbu8k2gCh3sWcVx8AvUIveI8RH+WpcNJn02YtknhMuhJ0QT1sO8biSJDi226BXoeFNPkO6EcabJP
w53SDMa1cKPpCoJ9OiP8obBUchiM+egcpVvPSaYmdwfrEvj7ynrHX2yLBYTzLtXTNouzqy8+/OZb
tcUrj/RN4aNUQoar0lnvDMnx7Q3POBZuRwp0FxR3c3KfmZF2YhvvgIrSrPYggoPAe1IF63f0osvt
8mcBuHi0tsg72J4N7d15K+lyiexVWvHU00glmn6bmyoLGb66J3C+3/T/JaR+PUXVdlFEkb0Lm7BR
f8opU13+vLq2K/F9WHKnY+QQe2awtEI0iMpNv3kUHtyv3WVl4G7CzipKTe7DxJ1QmUGUtkqT56aL
TUbuzFjrvJEmMA6OQXsT88YvX6mRAna71lVHcIUAJHspF1XGlXI74ERwrAlWhqHeM+D4+amNVMdy
RGltQNgVpHMyGLajDqtWHcewwYIyAx8z9u26ULViPsdw4HeliYx5RdgF1TIFxifRgSb2yr6lp6F+
QdM7PG+q6uSvjxi0I1UXHJo53bvYOtt4a25UcSz+Y5O1Xzp9/E93EvA5TKxZtHFfqaDg7uA9Zq+i
/WXIENrouxeVvGOfLlxoaHHliWkQCdohpptKH2m63FH0tpfwgmE9BEUxwh1+SsDeXx80DlcU/m2p
CrS+u93QXQ4T0Me4Oz60cATAnmJsZS/jXI9ZpO3Ngwzmy2/qE3SepM2YgPYwMMrtiONmzqBBtlJF
lA75/Kpao48dxXEESawfh55UYULEt1i+vvg0dLdAzBG8nPFTLhaQ9Fb3P7LmtofYkUCZrPZGBF0P
39Cmg8jPzTWkSkIW03N+o37mC5Dy5XL2nj0jQNR9hOzSPSguR9gfcXr8SGmR2i2FSCy+jSLXj0DP
pGL8/rN54qye9tII4no3oBSHTLj3yzBcKpbzQoJxpVeUFxgspgSBFnIrqADfOwdObjpkK5Smi7o4
A+oJBf81z2IDWJH7F6ki9MK2Z93bBLaWfZey7jMCw34hbTAFsUR3rxp+yFDY4g4kCwKuZoJ9z6/k
dzYmkYYe4N7fVSeKsHwO5ypjzAhZ/PqK2vfoOVX+lm7h8u/96/rxnQJM5zhzExquhk4UQ5niG0Dg
OX4NBATcDaB57jJYe0vvTd4IY3aj8oWA9N8PdoZsAAJflXM/FQJPI9BqU2GfPlerZNiRQlIdFEf+
ZGjoicaOAYSTmoaJ2bpa45u+iwqQ7z7l27RIjUzj60pQhQNj0lDT96m82KFb+KLvRj2vbLoqil/S
Njnzo/ULuoSSO7j6ESW3pV293g3NDkjc8Y4eyWJi0a7vJjNXMHRO8GsdOPKtVfR88LgMR4sKDE1X
fC3FRNnnOOETAxaNLyU3hBd8Vu0IGjuFXphHQO29846/N8WCb8aG37C0ITYHBUq0OW+d+Ptc5D/Z
Jb3TsyfZBLmjmMpoHQJDhCpxEuZSBGlekKsCzPsbtEYiwRL2uvnJo0Y2LVRskn2gzG8GCDhdIFXF
3A7PUfku157p76ooyFAK2FRYwuNLBt6pNgHOa7O63anHabdq0E+feYAjtTApTbUXeAICNzX3Mw84
W6b9oPHvgH0w/7jyZNoViKVOO6CBBQM51LnypkPWARjsqGar1WxbYWVHC/FYcO+P8WgJxRzAQrir
jc7I9J01C0KaftoejUKAPWOSNEYVffNHdeRLmldAcEm29M4672zpCrjSCCY2VX6qFyBK0ujmmc7v
Iu1DQQrsG+CxAFPErYZZUG0agmTTJthxTsIN4duIB4J76yn1pNX4bAF9ZU/EQIGau3aUdcAhtbqm
/s/8EWuAfheJSzQigxJoTn6hg2HjqbHW7Jrv4g71s2nqL7GfHi9vjTzPZcsBjUAixyo/WaLntXYh
eED/TWi8kLv29Yx6OYsloh2LR7wOTpqhCwTdHe+hVVxna2GibwTPa3B8WOjQKsAi4Rt9Z3Hb+ebc
GrGE/ajzq7Ga+IBju10X1KuihxgCWgzO/wssDAt/KovYklLghEX9cUdlmCCLvV/iFOWVm0fNHIpO
BknslFOkq7X40/OSfyDZr/YiA0VaMj1dxVABoPB6XnhS4t0gsb08ziJ+BumjiOADPm8gLe1dLyiN
u+kLOOXZ7/dF5QWzFE2QLoH/zevafSOUpNT3Q4esOEZlXz0bu76nezioljP5TaeOvKlq5hzIMMl+
5ZMn+Mf30gUW/cnsRyJGn/n779n/2wrjL6DzOzqncwu/DegfZxCwZao/nlFbehlXVWbD3Yyitf9X
zuninIIuvET3OIeDfQb4PeGHCh5BFYmdqPXkI3/Ba96BZVy8mnGz0eYdDA05koQEp0mP6gdHxUMD
RtU8NkcCDIZfGH6erttfpQ4TxumP7IYffYMV/ROPghAveTqweVzwwXTG7o9e0eg31gMPLw2sFbJ/
6UFcC3wwRqE+lVnLx138cJThGw1NdDwrp4+lERJENt1lsFi5swJff1O/MNOG7D+9eIi8oh3zKWc8
uleFjs6e+Jv4e/aMOSGWU/g/hqFdcqGVGC98Sgw71iZv+rbjaBJWciSn6Wmxr3pTYuSMlhx1JnrN
kAa2Ihru9JTOLAHWDE/A3/SwJ4CIrmZDTdeWEszHOz9axya9bhsnRsBkc8xQv1MOlIKG06CwcxyZ
YAqTnRKJ3c3WwtaV0Zh5H2d2bu8WM2jITMrdrW+bA5nIMf/scudtGe458F3mC+u9Sp91YHvjg3CB
IwZENuwukxXjl+s8A5YaXs4KGLK0dPUPBOImyFg8nqKaa+Ty2HwdAnrZIKKybb6tJxxhZpEmFB4V
puh+tAwbm5bHd/ieeKYping85+uHPQHTMWv3n/7eH8uQObLp5zaOLBylQPZy4TEYC9uOIiDfFzkz
4W2WNooM66eZDl0WAu2/gvcCX0ZX8fQz9li+4+YZt06d9bNOivLCAS/ykKtTaSehJzqWWZ8VN4Zc
pDPMIqADqwklohl8xRKZrJ02k9tbgDgBrRsaFlDc/IEZqUHvldcRKAbCGmBQNI86kmocbxmUJrks
b/GpGIKOBDVDiGqmaUJ0pee975SmsDMl24HnZTqkXFg/DQ7Kx69Dh1LMDVkA2aSEcrsREveycQVR
WVOnefQk9l/T0ccE0Ur2dvloAweMm5QVmPiQVHls3XZGmYqHmEdPMwudAKXzrIyKdYVYF3xLA/3X
+WsF/c+HKQZgJiET/FSKzbpB5RHjoN3E8Ro52aiQwrRMOP05TF6evyO79XNBRrtU/OQ/jZY6+G8x
LU1RsDQwPtoooPaesqPwPIeOjU/Sraf1slrr3uy+mvZOxr7+nUfFi/HugleD6jamf39nqUCm92aE
rxSFdfRw22nz/DITSA3XtPepBymcAMwBsir9MbjhHIX727lcnG+oMs/8emAvgDXFkIEwdMVforvv
C/B/H6WAZFpWV+X2pEM6ydqaWjTIjJBPu8lpdYpbJRPXgzlS6GSvxUveYIWdr8iXTDXGdOWKXtm6
F5EyoF53TLW1ZrZaBob210AHaRY7nyKyALW1obFBsv7em4gWKNEmk20Rr4LrHbYctHrbAwsPvDQN
kky7XyuspVX9CBk+Vzy/CoZZwYrnB3twYO4M5b63dEU9re85X6Mt9Euf8OXii3XdPVuSdbOwt1Xn
VkqXGfHCo8pJxAOnUVGoJy125Z6sHQZ0Vi/lFz6w6TSpqGrIDQbxuyKAZ5dDTmwRbu+1OZ4qXEot
absGrVDP7m2iUlvmOIZnvC0AeqFai5RIpS3Fl7kjb6mICtB3cQ/4J7WuUcUqIsJ33JlHRdcpP4N+
5fgQLrEQ3U2QrpZX8YHlSCiSeLTObwoDUU6DYnbP4l7shWPS2mFEVapQM1vr7yoe495UZno3Z+Dy
aV7Pbl6Fg6oZbP1iT1hwC8lJNfxzifF6BlyTpt9ICa47Sd/2spxSjcmm16CdAIxbxBCRzXe6/Dli
NIgZEoLgjyzwka2/JlxGuKxqcjyPXzk/4QtDXGKSlBQ822xDleKNQacwD2Stv3KeQP99a63wcCR1
Z+y5ppWe+x0lL38tak53kwEAz6tg3GabUIn73mpn7N7W8i0ixwb4CQg+IZLf1vznpUEohRPqM7UZ
6NY44gV5IGmeoiTRFoMOnI3wU99g2ZnUGvJiauqy/JdpO2uK6pOHDrEcfZZi8ssP7WjyDYPzghV7
Xg5R9ublx9MVq+lr5KM6gdr04MBwnZTJESEKYVwpjtBWuLn78OxyKkaEOeUV8mA21FSPLLy1ptDt
VHTKI2abACHWST0jXLUIvvNLNzmDhRNEDrYsPiR0A58gBOn3hdwWvaEAncUxVsIk5UqpO8nWus4m
4737l8M0Dmxhk+KR+ERrtL0Lc0ddPFtbzunO7dWzfti3FsoUDqrW2KoAVbwYxnTQgzRNkPDoJccZ
pjsx14cM5sT0NgzXegsuGUJrJzVBCk+vIHPQ3zUQjewAiUs7nrp4w71B4zJKsCQohBZ5m0+oHEnT
m2R2uAbnVgaQ8YYgV9+SHdOfA4ozD/eQR2k4hjcgNXRwZys8TY2vcfn/TxZisX9rUZnkQ1zno96A
fVU7upiRyqtnVECP/hgGP9IjP0qeF09PcICJYTJQjhxHrx2sv+mDJsPCSVAnM66QkOS800jA8a7D
W7Lt/1NBPQY+/F1C7WRzbbmffBQ6Cmc20rm+zAYLelwdQymQdYlvKy6RuGgbYspeSkj8Fd7LGRuR
/8HHn5vPph9oH/M7WK5oQf8UbkmcIrE5EnerATu5qkS/MBOB+Wj/0Q02R5Dl93Ea9inbPJBVM2M2
9BmxbC9ryisVH5F2kMxdAv/j1r00vmEnPO9wlwF2tiaBhJIerykYm74MDEM1BF+9UPamD6gK0Gyb
UXjrTOpdE5J2yJm5yHxyJFJjDUa+7FS9FpFEpd9suN/Y0ymkv+ViHJsk87x9vLEu/t7iPeYq5l13
uRmq26FHoQQuedxbFaB6EHOTSmiAEwZllGR8dfnzhH/3R35YP4jLNXXFkqLGOEVE85d4ebtwI6wk
FZ0X3do3LfNtJegs68pWQve8Tl4GS9KPjrlP6S3+6fz7VHvYa0Qqgp710eehckv/aVavhYpX0SOT
Brcfvav+FkAvO4C7Qw1m4S4faPtaXLyXtuaJnad8a8wIGwVarj8D0vS5p85sEI5aPmtYcWzvcAHx
V/Ivf09OabyKaqVREeH2wRctPBCb2aTRlBa7f+Fpq7MiGxMDEhpfbX/MzZezYMVkP1EGTkm+J1YR
X1xr+u1K18TSR6ZE/qz6W6iw20YOiUxea7W0TLRaNk85iWzSJmxslGut3f83Rw2C4sz8R8uHn6vO
43/yok/caQ/oXsoM+vi2XAyPBAGT4muKj6oRNFk8XykCLa6dybxQXMcw4F1hSTosVURNo3Q7o1oF
iL7NbKARv4xP3ULtFYXheTlcQf+Nvj87ea/npodmudaJ+bFc4Z331xMvx8WuzHJE/a52tY8vTRti
pnndQwgQH47WcC9XkaaS/+/Iwdmrs7uRlTG1VRdRiARz62PrervRa0NjB4XKRKZLoaSRAgheQJyY
TfNxa88ScEGFw9cVzH8WKWIDLW1/aHJ3NLh6nRSIELSPa5QtkfWLgmsoSiVyVrK2wvRU2psSAY5x
NA0mtGlKf9H9qBsvm3VQX1FGXLhLoIIwF6KSv48PRNkoS1QOik+cVvBYavQsojTlFnrGhl4IRSzT
8uPqzC5qGwfdX3x6ZEdWOyj97SLNnKOofChuTjlnaOGcKQ4vI38vf8kPgxoTfGc/6Wx9jkddbiMy
EDq/6lQul6pNEh9YJEjt13JLXlNgAcp9VXlGgqBWhgFiZIEkiaTZbo3wSuqwOt5ZBpYkMXhIFc8w
T4o5AfVL21dI6VraYxJu2lD6Pxi+yAJ6nEV7oXmfPl+2hyan40pYD+KuzmO7WPKloAC8j54BTcq+
NnInyiymdzyJdUcnX985c220KlKuLFmVwWvbUcVNK2wa49KqLoyTYSIk9k7qg4ditdODzgIKYCV5
IUiy913EQoe5cLYBvaHRoHr4fI9pAKR7R4CLQnbwCFFyffqT6CWunkmgHJJ5R3601zltoY8l9FYS
T9N0MjpCVTN/wHJkmYQS6JrNQHezhNfOHMkoWGM6JpPgJinMBXwYQLGNYbOETOUbZ/0jCbh+KDMz
5iE5Vq6NQXcoXgIGy2PwYJeBdGUXsEd2odtpfCV6UGWhsJQgNcO65JGm5Iv0WFgsY3foN5KDZIEW
t2NTtWT/rI5OP7kdjoId2QNxhCgVN0mIpoLe3smcY21dcNj/zADoG7gyuD7CJuUhNiENOxrJIl9D
nMMBWcCKQ5llATgulYhwo5eUTq2NFkVq9lvxmdRgGebOPidOnKEgVUDxltVxsbQB5T9kJvYwTLIa
RDaAchjExgR2WlxXcykTSSnj2phrTw9w3VngLp3fr+v5EQotSTOb+V2qECBIo41lcYW19Z1LanYD
iUe+nTRchQDT5l3lOJ/hDobLDyl4QuY73mG6DwwOPUtnUz4gTdzk9pE96jyHtuW2aeV/DFLVOTVQ
13rvlJ/s41ploWMJdYlkaFFoFA49I6h21WlQ5G6W64HdN3oKywCqrDNjGU3kWeVSJRPV1U4kUD37
ubjTTF446hReu3QyXBun22csR26HWSlHg5M/IPipdEYMMZwiUN2saI/GwnrLuL2czlcPfPzuhEor
h7cRPLsoG62QbGdi2+sk41AokaKMsTQgDchbmQR57f643JxluOeAYyIdWntT3FBF6d0yk54HUChj
NnlaJhZJ/05SEB97OVvVko1SbzV41QYFGCMoEZjfnI9V+KtrRDMfYeqcxDTKSSWKsLuzTWJyMyeR
BSQkCmPzidRoifSuNUrqD+F3JOgc7TCfpYOSRxkw5ju9DWiQH6D7Wx2sYl/VKY/g000VO0a4o0F7
J6avi66SfQtlqOhVTroMfBi6s/P1Zzs3fIc9RMGW7b4ezvF8ywRd2qvssGQPpK5zraLVtWC4tK2w
4vizxFCkJKOuXfrQppjOTNwINpe00ReUIozzARACdjJjeoVsKkupah+NKZEPmrOpk6m4106Vy57m
oOkXjSGa3TDilxn3+WaKtkKSnyQ+VndacEA7wP4sE+u7s3Ud7tiB609rBhGbQPgEX3aVsoAw8kd+
P42apVCFwmFJXRL2hYeX80zkygY9A45xusaQknYKQRCcX/CVoTvfBBncXrBR1YkAxTi1LJzhuKio
8RRrpNCK8ubtXhgqRxdNvJaoXbyXLlvBYTf4YOq6VbtqNo87w+jcUvnfwoAHYhBfr/TXOaATotXt
p9eZ5Xzye7Eq68DYn7pgjxqvxQ5/ts7I7uWaYOk5zLJm0eIKBYXP/9MMrLk9RiJ3CLZIsT70AmDe
H8hukyyCppnc8KR4fRW7naTuNSK9RaNHTQyNX3EQRMxmoQgfvkT3xjkTIiha6rNkQQOuNxWiZXT5
6Fg9BB+iEeCi5QQBn6mdd0tVhR7DUGrHxb4eIFbnReigyZk3mJReYvzWHQWiaUeIHZRQZ0ydPGnG
Al/LWHmpzq5PLRUwPRDConiysYgSAWcLiyLFG7EXmE1vdvhpCSYRvH0qYbLMKUdgCSXhCAoI4MbX
AHBp6sL8ln+T2hoQrIHioDU81nz02ji4OZXF1gvoqjZ5bsg+jqpC0aerogMSgCvlNs94jlfstP4t
wzgChNyVlOBdj9eXdzKIXTQs7HInD1PuUaQoYolBZ+KoRPGrmltxBqQPVJsrzmZkAMentXvWuL+1
Gvoqi2bzyi70OeJ1d3BGCe191rKpPZZuPANSlx8fcMma/1yMzAxEKQoWCIM1Di7QmTp8nEEcSGvh
fj7CYGCk4zsHDiOoH3EuAEABm8WLxBFACMiOk5IhX5dbVdrCBrIeTTgx2qj03KTNBR0PiaaIfq0U
GYwlrHyPHFsXGWN+0JGhCFOEfX9wmlKd+mvtogXmh/2RYBQvHcqCPZuHSh21n2uvPWMwfkVR0ve0
E4joiEH5d2fmW6kzKh16YgHzy0XE+RrGtTIC0s8HvtGuu3x6sDT1expzTbdA6IWehy8GwOX90VDk
NUvzCJaGndbs7R2Eu5ZfPWe8YyYoWpCtTUwU0ubcLqk8NMQy4GKXaFCyMiW/c8ShlJHk6Wj5krHI
zjDLDIV2Fzqq8cBo/fuLAgvaVuL+KQTro5Qj4bFGeDB1HfjcZOmNcG2bZOs7eaSKwdpK+s951GMG
GopFYlPsr9yf1CvSMV/gbNAnVhQ1SYLfaU59vinwc7QayGDo2qI669zNL2pTJ5ttWj0X/7IROMzd
NDeBUoQi/a5l62dx6qRnS/dm7nB7DmWmtupuUb+PQd3cYUevMfhmwD6mXiKaZD+dbi0cg4YhqCE+
fpdreEJnx5VUcQ5IL2OHGOucTSCZbI8XDIV/DOE3RsGOAsfX7+6gII+VqL4JGIsSR3WO5ZizWZsA
4/LQhFoVwIZZELJ6Or1GGvDvw3lQ55bmeze2GfQqpd4zET9haJ+3UsRhI/H9BuL2PAq9OARz6L0H
nIvtlmjaU3n+pg9otoPZd6B/RNFjpYhyip3SBq4fcTKEUuU/pskr6Z4eQO2TEnoXdPXVi9DzZMu8
HYiWbI1//ZUS4ZZhqIubhapjk96+6aDBZaphg5qhTUIIedn7jjvpNzV1tQIuVcA95incHOxxVjPU
0vEIjn/FJRU0xD9KtJVfyECR2JGCtGU16igHCAGz1rljHuMiZYJKhKU8H1YN79sYxtw0J03+3xLx
MlVs5mxyT7lAFu8I6Dx/PHZTSja1b1s5U9M5mENiAt+iTBzO8Ich7LrhZiWRT2KSX011UiZede6G
oQN5wum+vjjMUlXnxxzegEYiiAqkj7kycpkoxSGf2Am1bT9z3DMXprYmT584YaWzoukBFwD32fdG
gDawa6+50ACSBYXdRG/PReJxdeLc4XelrOxk+EVrbyLtRm+kuIdaxHcnDh53Kl0KwBTHJ5Ewg1/E
J8yFgIm9QFhwJHAdfjNHt6hoRiFPIp1VmC2jFojak2af0O3MVzdzkm37lkeUgMy9cVIQYYkNSCg4
5+6J1FMm0zs6x9KlyQx1hgEBCkyDLSyV9A/poY1wfbiRrjhHF0aoTotUP1FYrBz7I86S+PJafcCN
+2NuQPZmHc5hLAZ7fIdpP/7boLWNNil7/aZ06KeZvMClI3nQhkvkux9K+sEr9uYUo5oNix5FkEwh
KfN91Z0u/rayZDutf5hudEMMjWCbWWy0T09WOEygNrDKVZsYGuquGI9t52g2thBGkAfpBb/hK0BL
ynVOU/uqO4cIVjiJWC19Vu1/jWiwGUmJ7RYq+KnjGdJPedN4tMjqZk6zEDZyYrUblOrxxFotK/vC
RHyaPDd1eSMHoklrWd4705T/jDt/m69mfBUJnJ9W2u2jAjY3WqVRrIeiHJQcF1aeNkRHXmHU40ex
ro3NLHYFCVb7Ffm0ZUGKvwG/mdmILiebBI8WA0PyhezzpsBXoZ6j/eUzQGus1ZhVSurblG2DebQf
TRO3fJ0MMYdH+bS1upLex6ynEH+RjvhkdKuRYk3/yA2lbqX0EDymlXJ5J8MBnLKiHaCvk3XlTwGy
Lks4KVuqQV1n+VWkPH6W7mr2qFZFLhJP5mksQl+2LkR3K3gR1BogycKBcLyP2MKlQ7OmiYZyrO2N
GY1bHWtpGDe0+Pe79ryzKj4JBrwTEdHuacofOfBCoBT7B9Q+3r5l1EFQ6iDHnTmgpZPFDGNvcUgu
0QERvwdNaWEPueGWW1XNrmm0/lQVVci+veJPUI56kJpgMYR5PM1R82t6gX88EE6ygodesrnzl8Vb
Jx1lAnFA140t/941gjBQYqqzsLBPVDz82aBZjed+UOGcn2l6/gLIb8VJGyGJl7PHETuhMP4ApAGl
eyIsiZKsLuVfO/5QPxDcSrpG6tsf2q991QOVeVggYsCbg7xmOc5AxR66VFUX2i90anbFrTIHR9rm
lf30I0hPSuYVgpnzKvFzQpRMRBDsXZ5obeLn1dzP8gsEDNJKVA+Dyb35qLUPsrom9pzbjm3K5SAh
IpfIyTpZqFojszM8OG7EBMkCVIfXL4cYE/2vS4ZxkccSe+Jk52MPeY/72lUSPuBdsEPIDLMLG6Wa
VpoOVN+tgFmwfNnAbVRqss5C2Fv2wL9f2ZVXVHcTnISExneZr9vv7ywJ4pm4liH5iQ2W1X9Nv2lX
K+u+FtFxvOkZLSn/1k9V5ISUD4bO+GNIveTxVMf9kbw9CGe70naZ5ZcfuK9uEQQxv42/yzPUO1mm
cYaaHtivOQtrC0UetiV0cNa0YjacPGeHHSWCys4eT7vP3k2GhOSGGM3pJDy/a7AEYuEXAaDciEKy
HcKE10i0ohHEqN3h42910r7NXMa1UY/y+/EU7F7OAWZmA3vQfjQEKqE7jUeZQo8FTYrgh/A26eiq
tnMtM1ykvwMzIH83yASJvSDAqAHF37LOMBXIrT6c/VA5gQcyxpK/1+AzOGAdeV/WQPrd2CszAYZ1
HY6JsojPOzu00z6uyL3X5dqoSfiE4u4qay2vVgx004/43xhA1J83ONXjCU3kAh3ZiJC9C8yxLiWE
zKHumQqjd001SiOnwGU9PJsGP/OnT+amZ1s14iSDcFg9rUDbWymRyCc4Abp5LLb3F+a3whzrBAbH
Clb+qf8dE38KRRW9eqpd4GRqeR/GVdNAq6oD3DUXcfXPX9uYnoY9apqAWa8ikQxyALQxYg+OL597
XpyDqqlRvo/hOrp2T4a0lugHOS91ehYHLq6Opgv3HqyoaNKcc+1Xi3sSBP8tmCN40x6+908uTwIC
Qkglwq+VCBRh+tfQb/FsaEeuhLRlxwaeL+OLjJTCNfwvM4I5CSoqaqoywefI3v6GQHVTYiFWmz80
MWsXevIm8wMLHOUZp5x+xMV9J4EY6PFmySAv85nDgwx1L367WczaXrkRLJxDaGjXykPkuwLqqGCb
NsSDzUKi/VN5f5sf/S8LpVBu+NbDZBTeiUrgpuuu9zzfnXHIG9uU9yUk0pZVWJBvP2JqMRbSyWq1
DzmwEuDWxMf8hhbgjdZnW2rEII8MCDSOtHuHQQZaE9EZsv7oR8EW/+qjkRe8opeE7O/xJHE/wKna
tzDXyRNdHPpdUakxuY6s4EA8RzthVLRv8eM+gvy118r/mpPNb/ma4nNGGcR88yKn2UIuQqLDQMT+
QvX+gYJBMyYnxdUc0jN4LxQSIjRMQ7sAA+KdHzGcN6ay4PuDvQMOR9zuZmuDq/lLpRayAoQ6LM0T
9PTlwdyw5FSR7K8/cc8ExUz9r41QTym5ckqL8rM7tEkYr+C6vNX+Rlaac8/McgE5t/Y6IjX3dyKJ
fmdMVfZtlnXj5RJzVsXwk4Jv4wMY1W/NQmDVV2V/SfcvU7FC6ZPK3KLyrHsXszXgRyvZEqac5V3I
gg+WSREvoDy1+lf/ZE/tnR3H/shwAX1wjMzyJCZKndEEZwSyevnXuNvYAydD56RfT2XCSFHc73UI
fYZjBo+terR99ThVcMJs991ycQibU0ewxqcfWdFuGqafd0wxEKYw49RV7bH+Wkul76DXM94JmKww
VsZc/Y0PfbLpNO+mJ2Ah3YUhx3vLFJwYERgtzhilK6rweXiIG72+zaS2v0mbuzmkmGTDkdbRXRar
Uy8EHASB6RGUgNBgoptPiLjrz9KBuaXUfNL6NH7ltAIL4xGydjixyZFHGy3F1HCcR0YitpSuUfki
KLEM6888aEv3V8Qijv38Zkj1AUArsGex8E0nPRkXQ+z3xAGx9fT7umzx58UTWSGWk/FJKf5RK+wd
1CYAQKjfbX6+q8E0sjzOE0Nu9iBqIy71J7cQ3trwAt6ujTKsnqm9FTyOK/O0Vl8cXvsZ6DHgrVZG
KtJHTcF+eF6yUVrLacFIBETNKwGhdV7CmvLUcKBS5WOv55iT7rn15Gp6ZI36e6wUyrp5UvSEAtW/
6Z2MJIvqgY1a1tfa01hInOtNtBsR04jgJG/im9XnuadtLCwozqJxh79C7vVyU5e2AxervemgwvOr
x4aF0BUdyQMurR3t8fBqaStIBD1g2aw8ITqZqYWzilD3WdhvstykzxSKe+Qf2wJK0KYjrNcThmqH
e0p0C+IOmmE6JsTa4pXZapp2pAvdW3rfI4MLngaHlu85UmwEQ/gbDrSsJu15VC9HiXAeu8UiTJ9h
pwF+BX1sjdkt2/XTTM6MHnktpPkE5gzHEq0uqOPvuzvU6msEmnX6o+tPAieE2YjQtv/95YFXbdki
+9AhoJpamqTSPGWJ4hiStjgmbI4i25IWa3xTOQmGJqQ44vKcTeM10ny1gpeIiyCEvyi9FEGGnNXU
d8HC8+gH7SVmWldsq4iGFFRXWk8dY9GJf+gGhcuO+2zdsJcF8kU0cxhzhZL9rz7MFW1y5tVWnERo
S7j3+EyvAb3MtqnSRuYx/8N2S3V7iMXrw1yvFVaIn7RCK5MHJTKtvnJYKRNc4Q8ZP3qhDR6ZO0K6
YpN/PGY7HFbRj1q27a8rDOXo9KiJJgiVTtgN2XiyKp1/3KFM4UAJBjbB0mb6ZkIxvGXaNNcXYv0N
RXz6uUm+DxgZbL8VjiDle7Fjo0X7r19QIKDXdNFX3oS7WmmYK3l40Qjp7bPpCT/WCZrHHLJqmhCO
PpkFlINhMWm/Z1vDUtUNAP4GtC6mcMsMQILCndVhxiOhbD83gqJf1xWpmQzGWZoLbs0SP5I9qC4G
fwSWT9MPqk4iLC3LdbuW/XBLwGMbSB1iuGgzKFfPQ9gfC82zXlZNvV7FzbqsH+UVBeDyIdaiUlUk
hI5kMbtZfgcazhGr+WI1aMMIsTrR6i/QMn6Y0SjBXLz4FJBIqtZWCrovmqyfKZRHxhONpRMINHC6
+TGJ+tiTUhoYtFag4mfFp5zhfe35D28fWIR4M/s2BS2QN8MJGSohX89HJkHdkicok8djEHdZ+Mj0
UXoXoJhtJFuADbeOON93oi67IfzGOWxxRn8kR5oEbGch1nknvdWR2txLJQnAITi2DbRlVKQgRwaS
HljYjtSo0SBPEpzun728ck0Xw0pRMXC5ogs0rnORcS9OC1fiy6HmfdYBeCntY5nMCzTQ9wLG8QhU
YEeSmWNImCCSJJ/HeM4f8rHd4/brdCVkIn9+REfslPbZHPjL//nW2gFOijyRw3hXMP4uz9GAUcCb
rwoLLlPCcf5QpgiZwypEU4uc2pThL3rG6Wnp2la0zVVs5Z6RB6qtF5ikOLfEmGDJAiMNXwF6+DED
owZ4JdBzbhR8zdSaIvVNaCnVR2mZoZQGywhsbUlHoe1T2ZIvz0eZAb5B0FUfqG0n4yap1v3OpmgI
gVUJZA0wx/wz0NF8PisaSmp6JikCsdib38M7IA8xGvrqrESUtRVe/ns7E+7KOibOYa3U/Yi9cPWi
my1/NmyRI47MIgY4vbAgC0RXGi0xNwbk2xXorDDYrrNKJ7F99IF7gj6Ml3W7bhqNsnseo5ZxI69Z
tsgGp4XPqZDDn7HEluyPmAi+ywn2F0nYNx3w+/K4JsUjNbMXjPoRTERyqHXxymzTmdBJ9PmsY0oA
SCxGrzchhyjLZyTUlryxKclI2nGnPUiIKvinMZttT6AMsyVAyMbBe32Azu5iwCADD3ib7H0isYUD
E4hB9rDfv3JWdCyW/ZR1VJXwmNQRbrCndUVZXQ7ohJeVxCCP0U29f32vYI03RvdE/k9/8pcnpEGP
KED08EubvsSdARaEBIZvmWFfVdUUXDdPYjO+FmYp7d8rvkWyWldBNzTJ0R9dpvQfJiClTRKplGg1
JchMkcYYnKCnXNe9pH1j1qFX4xlxXV4ACBoj6dZRGuJSVBFD9JZBfdpAni8+q7rn54BKD9ig4f5z
UTy1+teHyLMrYHzblEbuYSKJKA+9cRkaogsluFq4+Y/806nQa5eO50WYSVxgVHjg7SlFFaX0rRJJ
XHxU4HxdEcs1iJkUAEAFZZIu8FPy2HQ2EaQa/K4rwMFwcIqG8NpYw9NxCfpZBZW7eXqIkDWUDJrD
iGp56S/o//7lw/Ps0ip9NHKzI0gp86m7AmXXv/iGTQizFfb3w1d7aEyYOZjxzD6R3QtBOaupgCzq
C/wy6kvDajdbDUg3lW9Fwl9uSTI2P5N7rKWidFDjGtiDlcvR5FIHQoi52BQE8aQlC8w9gZoUWAyz
fs3mTa1zACMvYfdpcjK/SqoADdoZYP93cu/uVenqW8eZuvdLbhZNQbsqf/gk7Ry3c5Dvn9sidD8R
wRFUtXwSmbBPq5Xy3i4MXacNX6ml7RdCjTcxm+eM6Hh2meXZ1drkdqsKAkf0qbcr3ELPYuEXkHsI
2BAA8WiVHwSOHKnEsWgjVK24CTw76irLPCD+pdIvgfShnOw0QbvKA6Zt7Kz5zJhz7VONbtLQ2f+D
B/Mpmf0WR0ex2B5cnPRAdXarN3mI41MVTkRw3/XHPOwz5i460EMec8gpqYsKLsPwd4cYYce24TsS
gFqmS98TGs0fzcvJZhADwXF3kPZlXqq/yIbcqSyBJWt2V9qn4l38J6ZrcRJIk22mWhJ7kLmHcluv
vkYuQi5CmQU2B5Va35g+ogfmGfCW6S6eDZ2+mAkIMK4hEXPvsbVhlKucGJaAkeqGCXJ++jjCCDsE
+fjmS3lOf0P5hWIgVnu8/F1VZqzhg11IEEYBuPgIdH0ctEDpXikbU9p7ydqxZfzeWRlU+qGHxL3Z
q4yeW+aO05AcoxMW3VeA8CXlo7qziXz6rZlrqJSkBjuynjCRvR/UyvuJr8sICSuK6+79yWo23upg
aGDOVMmRIie5CKUrft45q1m7RpRxiYYHNSes+NtOPiETrrij4k0A+Qvap4WJem0RW6zMbOgAGpgc
RdiqYB1tpy4Lae0EqlmALQCYwc5A6HvPFUUrljOn3pgBldrnzViDgbQdtcUr7rnYE5gKZklIUNMl
H+Ck2Wc8nq1hU6Ix87iRbbxKLJo/UjUBHJaUBSCgQ7MiRvS7r1a5/4X2eKticTuZUiWn5/Dqi69i
Tj32v3HpRKH2LmESPpiTSGghbqUF+AV+KToe2AZ8jmYlVPXnf6iiftKz7LRRFoktJpsN/y0DsvaY
nxsvAH1GrLyfQ/dmbCL6fcf7V6cmxEQXA/WNNZmgisiSrugXUQtQFgUyP6jeW8mtgPwLbgwayN6J
BeYaYOMQk2SKYcK+NNYJZTAjAQg8od1aP+fmIKaK/O7TdPZeNqTbvlPRcGMrqP29rOyCr4jxNYKw
0CoUbHl4nO0qFLJEFjHzAvN2YNOMdKDXP5NP4bA6MhdRUixJ+X+RHlSZPXei5rQBKTGGMtY95weG
jzfbC4ZOcPFT/IAXJ/MZMnMRguVrPy75EzqLGNENPVDGEdgH2T3Al5ylORg7DzsoyKwMaXPZeOXF
y42MJkF0enklKNRDLtB/094pbKF7uUYsOhH3EP+Wi5qEKrlFQlkQ8MXgL5pruJ+wjp/dG9KaTRdt
uPp1FcxNkXSgEEwYeGtkPg4gIoO+nuoXzcFd4IJvgXogauZEOz8kI/XX6Lx8uYuqg+FtMaslv7JS
cTWYnX7TpWc9i8C+rhYCPNVpnSK9yd5s/VjYo7r2dV3VN8U05/Ok/3EtOhFVwSrpn9PrePHPRxDB
eHWfYDzSJlbHIW4h0YXceVBnyxpxqI4BPXV5qe//hXwB1FX1yRgqafkcKAYYKEBDJ78Hy9CJmj1W
4oH9b2Cgv2ahHZiWB7YHZdNraEyBJrGgrBdbaXF8zia+ihBaxV4VkLu7gld6lsoJcP7bGI8VyONX
givMkIgPBqO0XkqPWrTePYuVrUAUp2385/euAqeo0PKeb1VzSl9/7gVsxLKuc0F99vdIx5QZI2tO
JHO4AIEQhD1paTcQCa8o+MtJbYO/HZFRdFsUBJYadse4kS4JbA7EfP6w5DQ/LODd3+llyAWZcG/H
JKq5+fA6VoBjoxKeseh0eT8e9F6j1feqfal+ZCtbb9PpAfBuRR030gH9901AGg967B57YdX8aU6O
oAg0aK8jCvMKLcRVRzQjh/CEGEh550KhsYVu1IB627zuF54A4dY0B7c1Km1MUr3EA5igRBTDgy7T
OsLTUtMjnA95Lmlt96ed6COYFGdadn0ODW6g4JDrDVz+LX0+nh0gHuxtnHYniXtZaWyvuu4axvzp
Sb3cbpKfn2OH0O3ZSjR6mBT7+i3uSsRyzhtdgIXa6UsxFYLqeMAj5qAVtpl0WXoaXlMjNpWibRLZ
CHKJIfBCj6P0Z2XVxnPfuK2wY1RkCHltjLr+JYksvz/5XzS6fGcgeRshW9TzRD5mpS8pCfZJucNN
kRKgTKgabpQYN/rMHmm8rhoXhbuIyReCWSMl9Rp9xZFTUTFw08gh/NM619lWv4zNLg+2mnnHX07B
p7uJQsdyTVL8uNNszYJs7+FHsdIUTf78PlEbYi9apn0oiZD/W6dK7QHJ3zGjiyn+bh1BNmkBEIGo
LLhLx/cCx3eNoWZ2TzZx+MLL1nmxGZk8vFKav+TgMt25WvOaNpJ4B0NClalVuQQmjj9aFNpUM8Xg
0hcEbNAAb306lHD3jOK6cxeMyyDtWnUc+d2S/7OdTCFwiGEnqowH9fEtb2nCd9n4bRIyb1X+ZEod
DZOS4vs8z7NrjQ0nFP0fxT3O0U5oMfUkg/6vc9f7ggFQIfQGTtIvJypROTcRB55MHFMko9ZxnisC
xe80bYpzlVG+Sph+Bm6WcDgg19GVis4aFTT5veroQDx7QNdXvEk9WfInpe/h1x5Os4FD+2Vs3wsp
ahruzIu0+aWkI3WbQ/w+Pu9SFVjk23GZCqvIuomJ9+Fqc4GI6/oee0xxamdP8UeZVKfdHCOEf2ov
c2CULhvUzuv3FWDm98Myqh9GXcmWL2RVm606mFGO67903CaXqp+y23owLgvb9E8pvmKZw/a88Kwm
9kMH424ABNyDNqmGeX5MfZOJM6wDFuwFb4H53BpCem5vFpOKJqEJ5BM4sNFKUA/O3naM6wIs4sd7
Bllnl7AynRKxp2RecddxeQHKvnaOyjFDHEOmEQ0SHgOfptRLrpt7huMfWNk4GIDXLwhfi5OYAa0d
VFnRdaPiJ6hb1c1XO87PiSI6FVf3Obk+nalDb5Q/PAAt6LD7JTJzwTppQ3ArlTyowM4eRo0prJWE
41fu2Itybu81oKQpNJmmVf33M15pWzBxJ4HjVIPs0hnMdmjqnwIV7RHuHibTXL0bkf/Cnhjy7qyH
RzLxeTmQYr4MfMPAYcG7EPAyKRvmISaqk2eqtH5Ei+coB3CIAz7tymDqzLDnHBt8WYZuNdiwQ7OE
JetVqoqvQONPU5gAPEa0Twti0L+VNC03N1pdzme38m1yhe3HA1f6cmBq0vuQqzWHLYnPyhKiOogl
ocfJoZrKTuOBs4G+0Oj8O2M93xG6mxV7Q5pB5Wr7ft2y1RDCDMCskPmq8/5vbrZjhQX+/UPtr7jP
ucZ7qvWPMVJZY/MY+SaJyaKIj3bfunJYyxxxU8ipu5NMd4caBKl8piXKoy8z5mE90jG0p6vKw/d1
Boz8GYyi96pcuJygLoeBiWy7NTaMlFVKzagY0OTeBVipcQukT39W7rxrt4vIUF5W9HuOFl14IS8y
DEZ3+QcgM5grnFv9MhpkG8fevIS4SDJt5P/tgK3orv6JJnS4xunJ7z8a0uXvwBxalwf5+6TAqLrZ
y/y5hZ+mot0WRwExzXSPJjEt0838LsVsk4SJzteEJkeSxrpayP6K1znD/gIGHN4nsiGAAiOXRmUb
HGxS4V2Y4TdQJwCEkiHntoFztf/ibBfAUvjUI8KY1CLs4AOuFk+s3dyGpKYa0xikazL+QRZFCrr0
6c4RDYb3h+FkcQNrb0iMqgu+NFr8iKpBYtFuijGhT38sRg4ijUt3Wawyo/skJHUBMgDyjR76C8hi
tVlsIoOzVLcDPThJhpbJ8QzoaKywkl1McTh0iYr9MoDSBxXH2ly0v5Gox5xkN9fKs/xCYvRDOwdn
h3uIyJOBPj8wezwYmKifmPMhygCWlWR30yYRGcVlhYW66Zyco7iY2kM2tV1FflvREmRBRfTFa8Nv
jLShrktUpY25SVG0yN+fRrZmYhVHwVEX1atdAWzgoh+52uGpB5iiiintQwZrdupJCXNGGFm2FqcK
lyLWnjzZZt7LnKm/6ggbMjEFHJ66FnxNm9hd7rNUfOVDjpUStqP3zFLdSpukxG8egYJ0e6XpqMEH
DTJstIvDLdqucy2vq66DiGDSF49zQC2/gGPt9NECVoLCsC2RERBL5M2YfVdboWNm1bwwcZBjqpZi
ja3qkxogv+OzzwFY983e1J3j0Ye99CX6RtJGAORCsoYUyxkLyQ/vbFH45BCBqSICcJdZTDI2Vf5S
w479MgMMpvjNKhasf/5IOqMuyKh6jF9EOyl8uRAUogFsI7CT4czzi1oDvXZ2ZyUwzMNHDSLNdqgh
j1YLruoI43qq0U1hJJKLcHkK4VGFljwSMxe5tlwle3ET0ETRHFWe45M7qv4Tx/Cv63X/SLXGlcZO
yHBehZWzleJcanGbRV34OMr7Pl/HG+Bb4U/xx17p64/Woy6mXKi4aO+sEHHrx71SO3p+iHcUob8n
ME+D/WePSfbxXNi3O3WMM4L4cA1gWGuQ/Da6paek3nmmnN61pSUo8+BtiTRFftPbvzZhA8ZP4Ki6
zchsYBFAxy20nnebWpmDWvifJ9X7FoST1xXLXcFYHFqYAfukwhu1MU1Jvax0SXfGRWV+1yqEZJry
dhojFT5sGOyxF4fK+d//jeoMgL5gF/T5sRzbw4xsgTlez6q6anzSeccst0HvGWCLFGhgwhGqBsBx
2zg8UGkXBBCoJxYb7qtnYOizRd1FG4x20sfXjusrQgwb7JGTj3j+5g+PYor3m2jFUE0+L0bt2zdc
6OVCNN26Oc0GPD9G8M3uaKV2hYqLfhdHSNtimTjbMiPHOy7ygFjRnUUFivTkUuUT0gOJOeIMyid9
WK+am/leBCgWU8z2wK4/7cdhs9BXv/dgXfhoF93Lu1WSztI9iUdB5laYEjt+vnWqH8jOywO2QZvd
DcKQ5M+E6Prw7dn9UbWQP76YH74s+DusiPlcTeVYnRIP1brg7eu5j+URc5VMsOiXwujONYP7vBCB
W66p3gR8J67LHxsDszh8UfaHnvcpctAodrTOlupWHLjRPSkBWkMRFzcp1O8E6FPWXBnfEPg58Dh+
Hzw3cFd1sdkBjdRDat5avjrrLuVVBgx63rEMRYY2n6mADbwzbPtpQ+UKWGEm5ximlbatnbExnmQ+
7FzzyqFKIOw4GYYHk/LdWPUYAMcI3P4TGQH1/NAsrDnzYLa+nFmaKHLzwKXZdMWodCJLtaex8TUX
Odm2RacbfAhZLXewq7+F2Hqb42yT8c34SpT5F1cRF7XfgGNW4OjkdaXZjAlpBwRVW3AlIAgHTr8u
TPeEXIf9BvTJZyAe1PC3NnXXm1l5mW/8fV5vtKO65q6uCL2W5hzGA1wAe7SeRg/y+CAO9pQMAINR
axHYTHYx2FKBC7fUC1RwZSwRobCEV3VCpkGV5Acoq4FklqinRyq1RievwUS9YYkOx05DdrWlkwhP
NjTg5mNurSUQnXTynQSo5jfCKj1GQAiXHvyVspD5g/kw5dsGCwH5oLMJ6+LbIjq2iBWUagWQCJb2
+GkgJGuwKnJjoj/crwfOKuc4pu8mXnb9mpaRgqRQov0Zzw6bx+yQ7cmPW3xmmJJz0Dwb1+rwQavl
ml65+JCZ+9s8FF5rmzO6ofC+pxGk3wF/SJYPH7ryjlgmXfz4BNZCPOeobAJ5hp+aqkDJ4B2tERb/
7HRIEx6OrNWftParGdDs37/nxbJW/mIy4dui370oUWSdPpzQBR4QmXE3pBhQoqJOh23pxM0Pfhbj
PjDPawL/bv0YdBpubJ/5Iox5HscvYKnq/Ofbmih0zUtg2ui2or7Pslehl+jvPH8/oWqB675XH+fC
MmUerndg4zh/sDJdCzrCC9IX42lEp/rYsw7s43kySwGGNB7yeRTvwBAtWDmrODW7MwoG4Hmze70m
azQP5y/cjYIJbkj6pzr84HWMl6gjpKJbvgSew59ibbeRsCLyCUwSNCUqwR6tsBoWJgofbIW7shWm
RKNJ4jCp8lhE1ws0kwSlBEohH53EEkAdcFdLCFHY2e9VzUVC+neTui3IHyYNLQ+sjb67QYPJeMnd
zky4aQ21wfjjUC0YUKZlbzwj1kiHstXN4WHV7loNy6QTL1NrMnIM+2tadn/m9xCaHrx4IFb4bQUI
C3rFHXQDsmZe8xd5Lx/BPB/YdTIX2st9WTQCajJq70+sH7QiIZ6f7J5Z195ERkXnvBETdJMAPew5
hq6xFO7tqFmP9U3uVIfpWx9FNMaJrYHcmqp1k6kUY7Qs4B+8ds3RU2onJE/p8aO/MzecxNXBolGr
HAjxub49pPPsfompTq0NNCvJXvcBdD2vG5WsOHL/YN9F9MpUthlBQLSYTZvbo09V8fYb644qrBK4
Qa1PnAFt0NLudPmlAK48E9S0npxjheEJABPO8X+pI9kdsL1/VVbnIz5XQRQkLjmorTBgc/RjpJVa
X/dqFrwj1OCSqilMzM6OnE2juOc4mMAENeS+5Eci0v2dv2WUJZVXzN+ZM1cMuFygD+e4s1Z91cWs
yPX/NRpo/pN71E0BQre5ztNswj4KrdyUJbyxTLFV+9r2hsesCWgGe5vSxT+JyKg03xMEyk97irSy
J5qeB1du+rlPNwEsjTCzZz0bI9ZNOGYljxCms/uYkh7JsxmICsx9C4TfBtvuN/GTCNW5RjmdGO3A
1hqeaK4paWt3U3ILL/6hyMibOPqfs445AHaThM6hR//7v8EpZG61v9mK5UkUxSI5agjhSbYUjf5C
3gjzSkPAsp89UtBrvoSPqZC5vP5I5DAkBz+OR3J1BCaVjLTA0qrQaYWJtP4+kDTd+CSS5T8/7a6g
yafiX+EUkGoOx3ZT6e1ok6A/8wOHFK5kw8JMoCO+8FZJ/Xuewp/hrwIddmvoPnIvVVYBGMnZikyW
FtciRq9ruplzCSaJS/3uHGxUliAZh84WMu+mYKjr6uhVv4gAZ+mzGCidULR2BxovybPC6RwefLLl
cgJmVtzICzkt26mEXgd9dMjKtTUNf4j0II8KaBSKEdJqZbBnsvJrG86bo0a63/AZO44+7DPlecxE
+PT47PLkAjQNoQ0tVriWqNAlp9ufvjjrdIprKhN7GHc7UeqSlBNGswXVszKSIJp/FAyotgmBPFEm
hIi0wY1sOi5mYOiIUB+SpPycmCR+3fvpVIoSq36vLhgdEa5FzESk4bCeAe99zuaw5UviJHHdk6Fs
Ka8f90fl/SaB+RNfAhyRlTi+Y9BoMjvcgveel9VAeQtvGpztaT0dZPH9z7zY0Hc7VaJ0LsEi6Al9
zCFpWCG3tC89rDDzKnzmp+EE6S3bmsfAybT0a02nwLNufNlzQFRZgt/YcYGzKY5hwjgUftCQb50a
K3c6x7OxpEYbukbY7NSxPgFLMs5smY8J72BmQmV7ztS2/GyizWyE4izLlPgdrvOC3//haRddGIFE
a6UD55d5Ipni9WU32U3Wttl6fN0EcxVoVq+WnPfFB2HESLQSdgHBV2b3/Mby9xz+pIVFoXabwMET
dG9VAITmtajYyXdyh6C970Ba6JB5J7NwgGcmRoHA7tPLPdjE3bkWqT0o5tRU8v4NSLX1HJugX3qs
mZBzIOqgXqSUr7XFN0nh6Kwa85IXlv/AZxU4I1KnPPHvGcD2iW9ziTxUEpv5DZv9zDWJBC4i7zkV
SXeixXU3w3OESfL2GmwoYvApXr+KLwm+3vbw8xBJv7PqPrnDOIqQt2P673+lbWvT4hHlkrsfAXIG
mXscS71xiajHWdkg1afCqiWRMc7jaWoRmLpgp8B83bXJmOYIby+aggyGeGUqHzD/dkn990ubKn9N
gRQkH4QswC94jZRmSKmRnG5P7S4t4STtLmwYjBm7jcNkwPibrNCYaazICkOUiAZ+5jfzVcG0VxEv
YnMTRall0WK3YHBxNzw2LtSKZ0LQxb4TOJJYN1nNkM+x8fxhlfF5LqUFBdu6OljU68bqXFtltXU6
RKWlWICnskrdr5bhpCxF0ueml+rJfOsQaiYCptSNiIsvXBF45n1+GgE+eeenkOb6COU6AKaTtQZv
ZVq+91pblCBqpV3Bi9zdbLI+k3crgAw2H3nhCcvecSLebeQgEhPgmekoxkKBDMma45zOP+wLp89u
j9bsmA8teCxpjHLPRUCwMQNh4ehf/uEDgMKgS+W1Vc/ZyPy/DwmdSZfT4PUiEodQfp92AYr08oUv
ZMVmuoTi5z3tgitCNQDPFp2+4tCNygq39xFWOmIwiw/JFCdLeL8XknGMQS8RNgCOiYM0nWUPokwW
gFk0rYeJ8EjKhFsmlxZNskZiw5ZLTf+WZb/lZTAntrTXdECvZaSnkhTbguGsvQZf5VbXKBgcsDw0
lGkEyRsMd47J8QB8uhKhfjlEvtSIIS7Ak1u1F2gImAF4X22EkNXLE/Xeodq7FcNCT7mxGoKzUh6B
qukPwFW3hra8U/WfLLrZSm37ZU/MKHfKFF3Co22FDqJklNUgXKr0Qn0wV/oCTTVRI2cjIp1Tx4yv
kHpiiq5XD5qDLCYovnnkbZSMnKisfO9WbiMokxpaTs7WwtGHU0G3q7b0DJbTd9UoglDgp2SSRvy+
xAldM84k+2nEPLMAlPyTBSNqNDvwD3joZlPKgjMjK9jZQcjuHcIRCMeYkcnOFt/nBesETf1jwHC/
jXd4kFikitiWwXqg2trJcQ+BbQc5/ILyXjMf6Tu50ah96LiFsgulxwVv8gIcV5knTz003Lw6pCfF
KXrJAbcCTCrQNTAnPfVBzOjbkqmlwgtIRiH1R2iuQ4Q5gtv9bTfvDizbWOF8yHZb1Zq6yEhybuMQ
Aw0ZO7b4vfsqRJ7mJ5MAgpunAymxPljF4C4gwPzDpq5y2o9nOUAB7L7f5jTWDLaN+lLCpEofHSu6
KE+39p/OEvugaoslLtao33+OyLqSuqQ7iJ7ShmsGGRW38QGagwNdexjA5zleLNs4se5jaeSL5K97
aHz7FCs/D88xy9SePTa5rNPniioQ2FeVnUdntOxMiBhLqCLK6qCEvosqc8CMjOr4Ee3Or7kJTMga
1w3QnLT3JZCp1fyEvyU/8rswfYmwncCnoqpw6rtZF2EaRhMFeD0qlXAR24bH/1+ElQtB20Trdzy4
Qh0UBt28HAy6rE3RJVAD0k2OBocek8w5MJ1quJ4XdF43r/aSLNAykLXWSm1SMInGBmFA5vvsCw6H
b1Y7gdv5sWXHOYLdIyFK+pYwellBnkiq1oBLFpLeTv27BnTqQClPYE6f1JioKZj2IxDEn8VcqgQn
SDzlJjOnU45I2LuOZFR3QxuWOc53yjMhpq6JwUx18jl86mC0r8l9uaqwtOJ6QJUK4TW19vGsL39K
aC6VaYOSKOc9HEmOJUVbJ8aQiPmb70iAfe258kf95DlaxX3AumKi0YWLo4VkXHsjfoSppupWkbVe
8iwYZV/XiyfW2IxkJjQi8/3cxen5AY7c3yS2S91NnrkruumuVmV8lW8iE1JQdEiMvZCdmJjEbBu1
x6gwC9wFkCoQ1raYwJZtl0l8y0HjBbwtO4B+3OrGE9SzGYihckJBAPwqbPBnMcpitntS2xXO5rIo
DGL3YnDpyJc1VLyv+r0CPZhpxstOlbyQuNcqX+LiNXVl7tdTjbKCRu9gYL3tTbuSm4oGWaJwUItw
qnVH1xf7eZq9qi/QGQ245nh5ofW8QURu0H8CcCzaXhjiwHaEMUjSJcc0r3dNlLTGM/1yShek9Z3U
ZZcOFs1yDTnUe/zjyAvZCYfZ+p0IqPtqL14dvYxho5qqyHGK+/Ib8L6rvHA1IoBTLhHPPPJfR5F3
sep5DMcUR+x51GsiRiM3kkoPQAf/WTdC6i4TeuUqcfsYFff0IieOPbEm0VFB/3RoL0yb9aSdbIMT
RnPkjDNGBRT5bi/6sZS9q3CjizWOXjrlSqdRxZDaLCptpP7ZdckiYo+pJvMUxozfItlJ6hXrwtsr
jXLc9Wp3AvgEKmILsqHCUFxCkAIexp/NBLvG6dRVxeq9vLb+Ec15shlPSR+Lp3fqMCFbKlHyzXBy
D6zUqB7V/x6Tp320UYXxQYuy6Tix5x3vHpGBSjYEfDtNkSGigI/D08eAIVCysUCGM9oVZTD0sF5z
Jn0uqktmhZicqntTby+VOFrDmFLTG3eD2VUADiGk/+6EIl5Om9fSjUcZ9QkxQ/e4+lk0+0Cvsb+E
D9xcFO8qSbVeVNyOMEI3ow0kb0s35W0w+o2poVu7nrIs+Ic+a+T+/GgPIH8rXDPj6g6CSvqZ7qNE
ZhViCpzoPRSSJyoUO+LMhIgntEUnsrVRDvc0giCFn6npfq47L8VK2oex1MA0qEyU3EDKE5WEBJcm
vYWRgugC/RAy1YBKEa2HjJyQYLZD1rLXPrRsUSpxbRHju4Hty4ZPxM0teQvOE4IC6a7ViVRxI8Hx
2bber+kK7UrPuFEHQfB4zaiGuqVZtPty2CyUzYR+uLpSp319N7HtGmoj5NnKeLgYiL9gbcf1VB52
iWaO7uzZf+xLa5rVjklub3ZYkTd00jrViULlbhzLlffTuBbGRgEl0h+Z3Frra3ff8TgO30Mzfw2X
c0GR+///mG3Gqr6WmykXklUamAC4rkEszd/321YPN+9lN2ewhBqnsk7EOGe5B3FgFwhhwRAc6Cul
tAlq1FfCNh2gGv/3FfPyqKDaWdrrM2QSq6IcJhfO7jK1lLfQios70lKyeLOospQpIWDZPR8dEtk4
ESzN4boaCY6yiinEExs6yreOLbwpv8ytspznZNoLG5iWsQYq2MAI3g3dISRwUaf9+Wejuqc3KD2R
7wEW1s3Uswt/3xe0ouFANpPyH05xZ4CbsIBfkfDA29hqYvqTEmCOeE+0218eQEt47EeL+HF2PDxr
itjBYpsf6a7L0v9D7S06egZZwY20EjP3s/zpTDyOPNxsEbyoXVkBpbW329pAB096JPnjJ0lLFkrG
lyVtMU0Pd9xnnhdwQKezHiG8HZOAKy7UKDr5fntD/8mzH0NfTpXDmFVdYFFf7OclwYtaViDbwjq/
Hp3ZEK2i/jPCMGCB8ZfzVVFHzve4z2kV4LA9lLIAIZRVknhi3i8ID++en8zYma9LEfy9YMIRyoTB
kTiG/5cRfwl5M/sXa7V/j9D2iiuzSDqbE6rVQ5pFkrtDPKIuUU99VyQIW61PNRO9u3ou/wLIl+bx
O0s1HEwTNJaSKL5wHFK/ThN7BFA4ueKad6JEih9RX1Fjb5cp5Tnj2VatJ0Jqo5JTSufpvOyGuO7g
NhOQP9JBYOmCkKd8QGz8Gr54R+MgSz61YUsMOhwntdhBxEfmpK70SoWV/N5VmXxw/GLt2m2cSg7S
1627b5/XvBiVgalTSrV5ra/WVGkJaI+YSVZIMOJjuZyisn5d7IkCrpu1vJKHbyHPBbRVYD5gA5jE
ETqG6tvbMqotCMoV0nek10PHnuIyJCo578md+kLSzVAHhsOQHNUJYzCUegqXwyer0wqVWbq4ln+I
xTAxAts81hF1nFRPqcpLxwcE1CvpPXjUrB0R6uLIGLE3Ml1N/5Bow8sZEDQMrtGJXJDDU6Ctt66A
dittXMWf08yNRhFDRlYfIX2nYGbXA7R6kUZtKmuje1ZDFCKoS5GZr6dTRxSqDD2fXjoJfg7hugRx
j1xJoNpHymnBye+MNCKc0kZUPZNf9e+PDlWI+5JqidSqz6xFDX2RFS8XPZB0Wk731Oi+I2Rg77I9
8wKAZ2amNoulskuaijvJ2nyo4fJJpD0z8qpxZgsPCH0Xbg9LLLQXl/AytjQJfX6iu6x/k8qC9hjP
3AXQgGaJHGi6F1C53r/FyedK05Or42o+u8BX+FlX/VV2UdCMJskAHG6EOY596M+dEk6qHEZSgRbW
QS61hGVvC9wOh3YLPBVdpqsMiG/Wg8UmprP09+8r8mJBoO22OkS9WFrbE1QDzY5vXCxCDNRY4U82
6J7S+7SFibzdTTzt0FSorY/Fwmcx7vJsIwa4/6A6yLSz2xwwbb0bVAKL7kKMF2+WuIEWFK9R6Aq/
i8u4vjL4GdJfp0SJiKjE1UWd11sm9blYZc5XVCcrwb638QI90v8mlzsuHlPzaQ+p76ektfQoifaB
sEFxBKlDsAyEuEwvcSfTJ2CtcJnZ2QTuX9BgK56gM2bQOnTz/9/s5TBtItXVq7yYuJ3HNWe9rgC9
eJR9604QIbfM7LPc9VFuOf11m9Kvh2nVPoMdhQUDsZRsuHFqcK1d0TnjEAKI9cSLRDeAE6jw/mVj
luooSSKO4ud9JLOJRF60iycmOId37Wu2Cs+nC0cWzgnHpYAFfC9C2GlTLlH2oW27DLXaMqHUHA+a
E8UqZ1BuUzS5/zaCitcVHkefIERneyxSIs3gXSsr6fiUEfJL4v4EOShFsaoe1VzRzNcEig5xUhiS
bAYqaxbGWnzLePEDF4WTcsyZY6KrVL86n0Xjebsy40ash13ZqHsewBDg61BqlZZQaKPxIYJT5dh0
TuIF4e68WlYY/lSKJeaGAz0+4z2sJl04fxT5UGxkxlr8E1PwojIqEC9yDQ6+paWI9H2fMitdcDG7
7Mlqmq3HOTNjUt2A8u6DyaKKdmGlPiSv1cT2cetY8Ae5RyiCpYddQ48S5/uax+sCPIqZ8bMYHvb4
0+aSSiyjwQ6qb1Yi4G9W9hIx3h6vxfz2iA0H5PW4tvJLJk5z8Fd1LIL2E0hv9z2xU61nvEM5Qsct
mJZMuUbl5RUCverqOfSB6Q4Crj2b1+8L73ePgZJgsS7I59T+2wjsdQ7XB5cTbblTwFW/2w0rEluI
fEGryhjqfRBpChWpD1bq2eR+Bxb5/lwELijTxSNC3DMYp+Qdc6tIInRtr4oBOJhhHVM8r6q10UQD
2iaGSdCu+gFm2REQcGqH2v9wHJ/3yrTjs3FFA7+Oz3vkfkQ+bzZqclBr8ux5a3kdytzw/Jzty2Nl
S12Fi+YCOmwIPc5l7TPwvoDWsvy8xcRX8GB49WBkcUEAFlSf0pi8Rnf+AAvACpB7zwSg3L6VG9HK
CBevIfy2osmiQ+54bFYigsprdIW61j9Q1keF4UetLQaMSXGpsE8FydBRvDGa/T/25m6KnVfTBJ9Z
QxZdlH4SrcDa7wr/NivOK2gmhXZRd8mMAAqozZIz3iLdmeEvpiUQdB8zXfFocIkEVc2xSAlYZ/Nq
w9+XRkELFf4yWOvfBfo7g41CaIVK/1h3WV/lUl32y2xsajJ10YlQWUKeX8jVxl6Qkv4kKVVw8XPX
2tuBOSX+OtwTlwPPsJOZ+chw34YTld6DFuQKVxSvgfZcwDuUpQjb92avZm26Dzi9Fvpvg50UBoGF
IopottX8cttTlTqnWeQ3ypd5sX7brQ0lL5aPjHtUZQ79Vqhfpjfndo7ULtNpd4FohtYbzvbE7wLW
qRGLS9cALA5S2q3NVp53fTqW7bjoDh1nE3aFVH1ISOCLEhhYQVUP9JKhblhoObfBiKWgAWNZf3U6
RVLZXJhWDbPmjNQKuRLNn6IdIwrtML3dUn9PW4i52ImctNcY+y9kQGkk7MFvBANorz3jMraqkUTR
CknKtk2y9HtXSV+szGhr3KPX+fA6miYcLyMqrjpa6RIAktr0FTYcOBXq/OowQrkDzdkpIU8blmtN
gnKRKdkIyfefifLao0/JzZx62ZQa3/jDMl/FrN2Se0OQ89QtKMDCjYqPgoyfH/+e9uxU4Cumg9DF
ku0sFYRe4su38V9nVdmXAt5/VLctbKrDOv/9qQLURK0YatAzfjy9Lojq6dkjRrCyFh6oXrtXhZTV
o5MLaoafl9BuryxD/5kgX10OVv7F8nJwV+AbOf8Jfwmbpx+XdPgupcyPlv3bodJZm6CgW9l5u1ju
fH3x9QJ+n9yrObvN4iPZK7G0CppY3h/5IbD47hHAUgZ8qUMHu76YzUKoWdGUH0CBDUmF4/k8QF5+
aJE0I/gGOrwuLEDl15GZ7obBOBCZtN4QRF6ZyGJzB++vWS0Wz0zu7UZyXTPLLcM7BU6cUIp3NLL9
Nw0XfGsfIUXnhDeJw7nnVt1jJ3koCgYvRozx4hpx+Cgq1dQbWmEEsE4onAJ4/XBYxyHh/1pq1RCx
LRGmw8/a3rdlXLXqu4tJhGkbDQNbzDNfJe6z4E5I0fvarjnlvHeNuoCinrchH9libMU8pxJ/YkrM
xdyJmlMqGJy4sl2FKcdWckZXicS7GNrEXIWmoJVL0ZZDYFOtIsbf99kBPNFWR2xz5wOWjeIf76HU
fk1VJm5k7sFRkzY1Vq7RsYOFHkfaJztoRLQMuRVz6ODcnVIe9uQAE3Esv3IhPJJg1ZryqXbpIDWr
dAsprpql25+HsNyKe0EyC37D2785aUNDUJ+UWJeWMCwJf3OsuOUKdVRGMfUMMSoHyCNCKtzEQDCR
jE6LlsOqpefBTTppIrpOrse+YNCPdG1KkQ2Ye1frRWoEIhTW9s7UbuzC6zMzJvYGBy/QJLuYNrBI
8L39MbYFw5cVkQxOVAWatfZAl22/oGLgdc7+gVg+1Jv0FZ3IKoqEycCFWdFk1WxGfvNW0dQk3G3Q
/NmfOhXJIvGsuKIRM61hsM2CrSTTLzoUBptLFGph45APByf9LDThKbUOwV2ulMnxqKiv8c3Wh6tV
iN7zPxc68jKnszW9QpfvAYMNZRPpR5R+7kLiYJoMo0l9ImSwVXp3YDPQ1D2z6RIqlaquRFMOyn9y
qqd44MyO1oQL7Dz/7U8Lj8Nqhmnp5AWmPsUwIOVwo3beV6WjAq/6nl6gvH5vuxdgi9/LhYWOj31L
OH72EHFsFrksqJAi14IKbOdKrKyCwqU3WN240BL8+Da2UgYo9ZKRwyEhJ66/prwY3p2hHg5Aw6Z2
Ogf0X8TfWDUyc8XLzuFqxTK7bFgI3vcuqKjxz9WjLLwwKIZo0Dw/blgeG+g4laB8wolu7A5LgbyY
vbjs6TRoJcZ1T3h2RUdYoflSn9ghr2QI2r7WdnqluKghqIykrCWUKlvYN9QNUmOUF9+mINl4m/XR
ysv5hvHTUftuFgkdwVREpD4LxSRreHuIgyoi1L5oqtWPR8uBU9ow5Kb+eSGuW4t043T8fJf4Vcpm
qBInA5Qa2t29Snkk9dBku5SFRprcKJo2vnOyoLGP9Op1L5ABBBb06ntRb36QK9ByMZcMuEVJgn24
XvNpzBoCD0uuVOXVP4n2Qu/OpExxBBOXzPnpyaViSNcxSYAetvOUZriskMJX2vzGlTUz5DR02uPF
yTtzxcdt3AXEqG7S2Ao99JbkTspuyCSv0LxNh3rrI1nBEqUtCcyTjGCX70dQeA4wFA2BS3wpnjI7
SOSs+4zMBqPsIo6BSpVBzNbKJQjkvfzrYoJ3hZYHAUt9n9JEk9TBFXFYM3F1ZG7V5hgIWROVBJG5
VfD+1IieTaA84nXdra30GNuLN8xw7fTdayxDberhedyOyCIi1ER+CyZQ44dP7m8bQu94tRTIyXJK
EX4ZND8qSYgjtXonrDaI6ffvQsQ+nytuTyn2PxX74zLmqYkwgaZkxt3Hv+cUu5aWz8ulPTHpE447
AVt+m++1VU44Oz4CsZexD0shqlosFm2+GA3J7QIFpwV6poU8zj/2clhXN4INt9i05J61w6DJd8GT
wcFkKeRexAnmF/iVIlSR9A7g/5xSvG03RFaxbZmvspit9ClwgptMRYiR/RAY6eCyFfTjErpYzlnh
Tcu3po0X7PXMx0rb0B9iZxFOo5nPmr9ELlFT1JxpmxtIrunbSiMPSd9Lqs2pHXjizczpYIW2Oja4
zyowb52vO0nG+OIQ0O6xdPMdiLdH1mdyjlMHbx4eh+4PPIvWD3KqKRfbRtO8LA+t76eCsoE8sGOZ
XuRC7Tc6R9b0gNTz9VKipet8OfX9Xdn5sMBObkT5hB6e5+ttWd7mKeHZAR35+dayoh79tepjUB2v
4Xi1dhraIN9rhiNFFaAAV/yafKrRQmN4mjZ02bMUoPMOV3EWDwsQ8bP++78BmebLwLI/RyFs83fu
OgURIbB1BP2MN4fytkK57yZZOxHYR3WuVYf96FeeaOED83qAfMZIoj0j2H8ZOSP/23SvC8bxg7bW
GzPxlZkH6kB5ZdLYXZgEBNbPhoz/jTHO1RlmvfUQznUsy2yXUIwr5S3ZwizTTvFFf3LF8rlWpL17
nac+jcwGzP1gBw3YPUtTXgpQdmNTGnI3SQA9mpxRRRIgnCaXmSb/dpFBa6ZZZ/rQfVotpn2Vdveq
8125kqVq7WhXMzgT93ITavQwFLmbYCFj7bh+YzKmKLE0XkZ6iwj1Qa2U6Ce6gabXn3AocXwN5WF0
/Ze9ZHEgKFfkMmCX9pYdkVE2N3FYDBS19b/bnaSnsL/cvuVikLriW0VarUAJ57hFWtAF/UnAlMli
PlvtBfQsC1HyTMuemzxGmfUS3u5a6dOSCjpdySj2w5LT7WDO1kVbdbPuxx0ubPjaPY5zw54b/iZh
9eg2mUa5aJgkuLieqZ46NrLKwLKuJkDRFUC4rk5LxT8+s8vo+ndZmFyV7aEmQ6FColOYIjl7bHcn
snSJUuef1L17MjW9NKddHHeJyqkYOhqIREgWvrnprhV9LHpJmJEKeyqD3/C1blbLXQ4gMr7dYgX2
sAZhm05Fw7ksJfXn5UwYA1reIsajNv9E3yGoYnRExtnw+rpRa3vsJ5r/yrYVimtmdY3MiGpuNqo6
tf4DcKIxPCfwdCTYu7t7/WE7FRBVteZbvN9hpuzuPsILTP1m139gCCZzBwBF4cYmmXV2KOjlHOiZ
y7fVvnUw/DSpyPqPnr2svxAisYsHCDD/lSE4dbc28wtbwlhndmasU8KJ0U1CTkJfaVln1QHwDzQa
qQSUFjcenribmo28ePmnwq4heZkBWTqd/Lkap/XGsQV5rVBayKj+WBxpL/UUdVUi4neS24ihs0OX
pfq6SOBwcOcjUuBlkbyn6d3LpUz98s3TEQ04vbCreeqU1H5xxaL808iLtswz21w30fMNN9qCrwPm
6vi387tt6AccOVs19IYeF9vBioFcNAGeQhWZRx47CvkR8g6mQrSQJc+6kw6X8pR5n4XrJH2VyX0Z
tox6NG5gsqYaXtSkNroT1G2BtItkoMhdFfUziWEtz2273qx6yB7kDbyYKAcKPPONaRxUj7JweF0P
A5ZMKMyQxQnFOnxGx92aE4A2DJ8mdpF5IA1u8CzrbxUPTqIcy+ZZDpEB2ouwrDVHfTW7nShUbgv6
cnDAY3ITxFef7mZLwuh66b242N80qcNo0O52BNOwQ7FVzuwQUfcZXPgXKdRVoOkAa6GE0prBQApN
QaYs+zW4HjjmdB510t31uosw3GBX5/EmC3xHQO1gJmvuBkyVWdfPS4o861c1F8ILJZhIV8PgIZyC
jY4b4R/1cm2uVrQWUcTbMCvFSfnNwRJAPXaa1pfFz+qnVVr3AjaAHqPoWtJo6dpbQvXxJTdZs11U
pRdkFUOMubGUiUFeH7cL7IO85GYbyVmoEZ5P/h/79rMwkf+t5+NXishF8i7rXvyMvzbtSIJHPjuQ
PGcmHToPlo2hfARNBMCD9D/G605MTnNQja2JlfyZjmNUQuOBbBRMxWY5X/OuluyRlETfVQLe2Ovx
EJf4YyPwJ2WX7t/GpP38QmPzAO0EgSgJNgqRzHIb6Ndbnm7R5FfHDCJlp5RgL0koL0ExHR5edqTq
MjKAZ9FEyy7rRS4ucKH5UGA4C5O3ljz9KCiyFbLpszqe3HEYBCl3HqB/qtL6ZSu72pG7dsfJK63G
L4lobqjFSFsGxku6fIEyT1GJjfPd7oG2VCb5tOqSJFD5uSV3C9DCqinigqscIJxfFJgocR8nKfnJ
ydRVWVJ++NrsSJ835uDNV1EoyIJUAFrEWixMKbdVYEh3h1+2FyNLHBUu7koQPQmdf/Jcy372DSMI
uBeAvD1YB28mZizJwZRzpB0glnMHlp7o0IyjRn2tC21NQzdxcRrRLlSQZhG49eRjWAUz9U0YLkh1
aulxykinkjPVV+2xXUnLZDk6FRDAodGyrE7RpMWUqg7QR2x0/LH+ikXEOLMO+7H+6UmZV9zQFHDC
accB2BI/KkjUxTzjnQeH72nRkGiWES8psUgMCylkyKBvLQrTVzCuv9ZkstGx/4SmlCGNgrljUP+l
QtYN2MQc1MEBx/X3FTZme26apfrpoK18WFcYqmmnuZFRRh1OfBa73QlYh8BAzgBnJkNzxgvUWdL/
tywsKhsapEqI0ue9ULxY3ykbyKPKGIT8gBweD+zYyTID4N1trTUOvBLirn0T6MIpPwDyIbjraxdT
4McNVefSpVqW2W8ZwEVCgz2I3kKnUKwWqWgmmRch9GK7LDCKJbUDtO2HZKh/SyqKdULQeReB+bor
tLNFwRs86akZ3ETbAsiAg3ST88pipqFpUjTmB5p2OXB41LHyP0Hfj2LEl5BtQn8BIOdNGnl9vB3y
5wYN8Q6R+h2q9bwpj1a8k0G04Eq56ag1iV01ocl3s3fwdjazUyQAV53FRFxonZG2vn+ZzVyMsv/g
i7SjodHt5abplrPe4ftRgq0+UM8CuYP9lvIhxrHLIc4Z1oxgMU4xXexQn3WIE6MmOQ9g/af4PXOu
0G3+9BUGoyN69anftNY7Z++h54qG9tC+MJdVpk0VLhDqx41YPNT0Ckqaato5qzIiI6GI/Zu3gSut
9tu6TJVITyaVJMm0bRe9jD0IOi6oUzU3h30jQ6tSidXxo14LrjyQclP5fm4Epflbg2/BkTVP/ZN+
zM/AUaBaGiXz6wcstAo1a6nxFFF4jEBdgOn4vMhd9QADFuymYutSB9PE5SVOlih+P86Rh61KFR5h
wWPV1ETgBaGjCUht7jTXt6IoiLdV3t7nrVWOgHkSemqdkaFJL5jKutl2vMcdzTQasnbVXcXWlk6n
geQ5IBV8/7JGKViswJnM7v7rL3QW1uv6qNS6OiWLm32x1/sG6PHTcUnRPDgBHH3nJThaU96RNA/e
+hMVLPtbYD1oGYnFW9PiBjkB+/j0UKuFTKiTV2zYLlKkzqCC7NxnRTSbUItAu/f8QKDeLZIMNRzA
EImvINTA+J45vxzQSIo4RICIdk9SKCl14S5CcdATkotaIIHbxdommLJ4feLkRJofux1aSt9ImWLW
+4DHO1Zy8xzFIBYt7++ubB89L9DX9jei0WmfkT/rbxXvfbWSpnroDDxJ0MEpWR2uoHA5yXWmYEtL
ujC+xYxDLxFgUyyoiLJ97aVK1PiUiwzY2mFpNuU7H6jXUkY5uRo5JXgrX45HrWP7P1XgrxvyIFaq
wk9ProQyBoQV5/itq8vGlBfljqDYI/Z+rvS4XbAHj0MztrqvqhVEHJB6oXIr78CrJpMfLwNKFfgp
Vsh00a1NaKhiBl2NptqlBh4YrnhYB2/r14lHJM+KQhfYzSP9RkPEsnfM3Xa9LXACj8vP59CyCVOy
+jKnt1N1d3RwAmonuCpDKisvVsRSQzW9d+rT0ojpTfrZB0I/FrysmGRV7m81tzieH+Dq/RlvlW/S
a9pH91rQ+gUI8TbXHWirVxVmR18y9avZLbGpiZwqHaBwn1fCDePcG0apzrZgiXuXKiGbeCSSuIC9
qUlao8iUT+5tEbA1EeNwzNA/VkWshZv8CJ0AmHqwsmCiNznUNvBK88IZoXQBCW/QVti4q/ODRYNu
fBlovlwjvi20EHO5YphJY4V3Bo9TC7v5uEtu9YyRfZNxxtQ8RukbUBX4XqW2RsLOjWlu97XtiE2w
bSf0OJ/lvs8x1wicpuk3M0XtATqB9FtTXmYImuVDypIIFiQ0A0H7DvtL+3TbJ3qBqx8UwD0PjW64
WYw5mjE961u52bMNU8EZ7YvUezRzu3EcV1JhsenwfPmrWkC0V0VNRmF39XXT7mSM4C4OmjCrVobQ
JuVnXv5mMJrAnoVgueNy20oD/y15d/1/mmoo8PJEyIBpntz+qrZAuL9fksuNnDKyo20dTW8wiOpC
bhx4AiwW7t46+HY5WqyIQDFjpwl0pUGLf2NpXai3L1yBjYwEeFbfHqVKftu4G+FAY3cI6GIXRDK2
Lp7VFxLLLVdlEJ0ntJzxFXQN/UOkIlZG6c2Q26rY4bd4j+OcmWIBbpGmr6IuhKHHn+ATaSF+/vnh
5XsvwYVbAm6o/3LxsoxakzaNJ7NHrk9++4AYFbnH3DNlWJd/woFCHxh5coD8JPsHLNjM1oPMXb9P
dCtGOPwwoDDAspSSjInAiUrpQ/9DbhY4OGDPz/Md6CN7KhTZ41Zs5K0iDDotTRZs0GxoGPZDFrhc
M5vWb/a6KwEMjiCK9Q+YYcw9oIePtqCqBF/Hem+UxtQ71jAVw82t8UzBWSYodps98btG4OLsp7Lr
VYUPQv/010Zkkata9OfLZdbAoRGsLa+L336wuXxcpJyWEY3EfpU+IzBcbAsjuRuWE0yKBBlY5jxJ
v+Cz2c3DAzcuO1q6w+1YVG4MNXuweESXFJ/f14uvdMGzkUqRQc1MFKclsPS7HIV+gqlaDglPOaS/
DTi5OmPhfY+dAJvqG7Hyvrh3z4rshR3/zobJTU6KtQVP91TapyF9MmCY1kGSu+UBL0Yt4k5OXljX
t1nKSo8xMvyA/6WFjJlzYuMpFbghg2nADmHEC/l+lMj3mlYvLCCGJb8PjEzpGtRNyMV8jbVUDs8T
mtp4PRxpK7HLkgD1vnFbvuXB/mahRwsKqfUcg7dvu+MgSaVsWiqLBsr4ApBBpdLuyxvBxAiuVV9m
yRyJ2vKO1Hlkvi9LyTE/xrTZuURQNEv83yTmdLsj5tFsw1eBgcYIbUDzt8s2egFmKXIlSWFa1CGB
NXFSmikpzSBkbnzzH1zAZvPQ7x4lhWw85G3I/G22hrOxijxKgILQfjBGGBlHdUsernkvI1Y20Idg
mCKThcxUX4C73zVvNABvz4uLrgNfrfgk9G+AZucgV+hAFmCq8ASSazu4ERFULqI+SFru8b0DwltM
YE1xbGOJOgc7q8z5mtLSk/0ZFi/EDuB3tdWO19+bWdGNYRtgcHOVz0RBQfduJyQV7rXbPh1pocZF
CUQ5wS0G/uL9qS0mCX9BCXybFCGW7siveNjZecz5kQmj8TLvTCdIJAwDrY0rlzyPnDYgYxng3cBw
Zo2pQML6lNJcvT7CaMtUw1qSO7S4fHgypQeSMzfbH+cHFQnogSO445hQ8TcJ7QjL9fNI3VDvsJ74
OSyVZCFqzOTV7quXQj1MeIfA2Tpbc2neqfWPbRu2dGfQPI5vV8Om2ql74j6nsApWEuaPDs3nHAuj
pZt2Mh5Nfds+ufhgF/c2jUJg6QH1YfWDFbcT08zWv5NnZwd7ug+4Bc27tvXyqVjucaFLObGP7Og7
coOSdbvaU4TvDtvjVMj1KCr5dZu3YEsv054bF14G3JVOPnKU5tur5b/pPYKmYBM1DgTp5bfxqcPh
MPF3bwXxk6sethfKUT/QgpqejFS0ux43pIV1193ZCV80GqaHMC8BA9kJYQAZK+4L580wG36Akjgs
STeWyT6lGKM3AYC333Ct9TbX7v8khmmcUDWc7n/NyaMvzGw9aXo0K0Dj3Ge814zmTWY97Wx+dLAX
dgs9ZCju4jCpMSnpO1R3K/K0dLtzCJ1IKwbNHN1lnJ+Jm7vAOOY5bNotZjalfrAbY0ApkHDCfouk
fcKcP0hSMQCXAJCYfTx9bB3j8c8hz7xNzc2j2nR+sO1HbZC3q1dFCZKE7mL2BAbWG+dkBp/OrLoH
N/zefbMs4sKtb6raGfT7qqH/3/7IDaepmbUSPcgv0wVKZoNuXzgMYlots2n9AwobLBARgxBZOPrr
Vl21a8mINNOfyYeyWf1XaoNIIEwFniz+6DKNdwwj3/eLiReClupvLgITJEA+QG4HYRPdiam74ppN
JGRpJIkAEP6MKzDJj74kVIX0VchLEvlIVT5N+96m4NyvhB03HtLIwtSyySN5mRPaCbR3sj6TeD5m
7bvOnCMv0yMAE0othMHjxyVnW2MtgsvWNbzkCBzf00aErb2Fx7BN5t2HVm5TsAvNH1bQ5/OvOghs
XIPfZcvJpXHVy2qPiKCU7PiHzRWKOTGYJI9Ytd9X4uuHICbi5o5bVOAS+nF/gzxiR1g6VQIaA5bh
MmZJX6dpY23gsX4DkU/wRR4cz5b1eVboN0JXTAgqxfH4ZvC5BVT7raNfcwlP585j4UDvyia+Vt2r
B3rHF04ucqfCHZnbAoB1zjwhqCbFvKlMFPfL+p+YskSgIp7+mKv/35bhu9M9k2SbdqpNQXezInah
1PNms/A2JZ0YtXAUcBFxhPqtdFxFkG9P/+dqESfAY+pWLiFPmzDnU+Q4AhbozqKcNYhTh7ZGr7pY
aMxjwV+GFT5FgUayLSUJOCQou2eNvZqNi69NNA6cnIhcMv/3F2UnywGQOTTiMDanVBj7zq70fweB
u3VeI7r6QxYSmwNYqQNcDEvQpN8YkG5bD+WbLfTmDnq5Z09/qqXWTvz4qMS+ovX8zYSjZMvK7pkZ
f0ecGE1OZEKit22roPAJP8MZrVZFRwljBXk3PkrRwR1JN+6r24V0JmKwvvd+XtxipqjKsDYFNR4h
ouZ3IMncD6J0NmIggW117SuUqoKUIEsPSfpkRsBtW6l4epe6aei73lhfRbgIL4IuMIbeQ4jJLc6a
ViAtCsfao2etTbf2Lm0XQtJQPQlYkQiueI6ghwPyJLmKbBmX8OY1c7MgyvwvefY9ris0bOtx+/Zb
YSDMdo1z+CJo5Jc1tecRpciWcaTOnzUfD9KLasqlNQZuuThykPuThXBLypByB+AN7p6DLBIxkQVE
oBMuZF2FOJIHJJpM4KfqcpqLjv/AXjmXc03zs86k+rwrtLjw0rLrHigyPxujFZOZ1HfR7N8TtbyX
6hOzSyDAHwruu7EUOmoRwD6tJlB4icSgKm9eGsPiN6qb2HZkRLqc1jcOvw05pTv7qZN22P4yCMIJ
hN8RDqaVhofXMMybG0SyIuZNv7YearUtbu2lq2eI1yBlXU+ROe8wr0OVEhFnfJNDyJeNgBhGd0fQ
FdbVt9SNdjWc4Vr96/PNZC1VdoYZiA+Gt6VYSvRDhVldtlFuzOgProMk1mFzL9vhajlgTYiEog2O
miZ0Opg6U+5dj4gmqkWSftFb2eVzCGdYBdSAGSNIRCqDVTgYEMhzxio/2r/XMXmhbhi4b2M24o/U
V0+curPk5K8ou8QBni69qumikkk1X/f8gSRZBQoO+XEetsf3Ce3j3k9AV+gCE6/6Ieo5PmgSNMO7
38SOIcjF2zxT6ON+5gAVL6fKQ+0egJnSNAjVLeMIQ2mMXZG/vwlTtPjPpCteDM5aKM2bjSTrKiOb
ny6J0+FwazrGtwh7QH4wP0t/4e2/q5s7Riz+9iRoeuC606VaLQSaBfBAGDQ5BB6amQRyuWD7x+W4
7nFEAuazTaRtp0n0hSe7lF0o6+SNvGd8dQsMy5ssbGFmNVLqoqPfTdSPCfMIUxsmXtsojACDTqca
kkB/KRin+iMjf3zA5ZMAmp6vFXlhgZJzOGv0Tktyyc5DijJH8EXI/e8A2RU0xG4mbIOXFd3dbcvX
KM2bBMz1lImn0dt6gxX09JuCcOTZOuizZuKL3Mlx2WoDJ6S3KDbVmFaFFE3iiwRR59KAuS5HX+CH
t5Zmp5Z0/B8WB45Enp74cW/Fp84FyiTPcNvY6VaCbIfLlB7F4p/tIXbPkqP0ddiI2hjQBJZiJdj3
RGY4LNHJpmp8/iTf7YaOb3WpN9FjmLur2OeVP4sCtiH/sCVa0DoJ5gWnB+k+gJRTt/dZNwGDxdcr
JTiojgI8ZXuBMczs2NVlHxKN/RCqqMFDEEx/29LfYTqDyEe+D4eyUE6QxDFBKc8hslCA5Z8aQ6cI
UkxUj4ofSWVUt+vyVwE4huCdPrzNyUb8VmnwMOJjdyQMghb4y6vhR2oyTekEppEED0dBx98Cfm5K
gDtTn/fsfqLqVzc9+Kh/kWpHe9PSx2IqkhFRO4svxfyG3DAeQ4Ej//pgYSBYu3mX8B/MFlM8nXcM
TGwXcpCVvsrOB+r5iCkK0WUq5vQ/EdzWPIpzIikKMInfDgRBwb1Ss/r27PeWC9Ijegiq/D1Sirc1
HsoSmGF72xouoNsQURMv9bumbynMGWJBcJbroaAKmSDchUA9kJLXUL8qh79m9sm4xLWM4P9/f+DC
GadNNRwrpN6ntSzbf/o3dyiRrTw7J3javhX10bOSvGPno375F++n3idXQAeYQik2J74ogGtH32DO
Hpsoki32C5T+o8ZlchSXYvdYCI55UPka7ZaL7mhlONZ17ooybVzA4p1XScruOxx8lwmF8rTaFljw
lebpEB64Uim3TLV6WdEJrYQbFxQXptcn0wncqShpmTLfepfNKwkDcafYqZ8et9wIibZjdjXVgiM9
uhaAfJBUq5+i60W8eYW1rLe8OMFmKLYlN06SBj1ZS020DsdO7H+kMx88kCGmmTYIVApkEOATR1Mb
z+IDljlynBo2i6OwYu1OFpcXYjFnwIpfOAmcdDl51ciV+Fcx0NBQLGEGe13eYfErL8X0B4DeUcCr
dIsTXo+iq+7wX4jZdNSTfuoF1MrEECXlLzCQvyGjz6agGh/2f25gYcX1art+65Zhw5BxJmqkuK8c
RtywKe7rxfbYhJVKm9GlB8lB9V4DKbp4XNO6FViYier81uvhqHmleTh8uBFoDCewqPktbMyAcnGq
0ocUIJppjENX71wsewIfYvehBSJpv7XD+5WNosejU61nynXSKyMwxp8YcO+ja7V2qBKVD/iLcCCK
1qm/jsOtiov0dEg/+bG9UzeL6u7a1ESMB9SNSOkZ9Z98mhRw2rNVz2h/LPb0ZosOkVvXOKEH0TGg
zQs0wS9yZm2n793+spuPC5lzQ+MjbaNCzpNN/R2MOl/yYYPrg2HwvfZIcwR4ShxaZSpdabDlTita
wynaPZXzhoI97ZxhC5xDl/jLiS2DnY6gjjC3DQbgnI+r9Y77OSIFk1swVcuGMYZfQGz+f0eUFhCv
+2y28Rp6fv6WmZf/quqoS5Ml4ttIX7dnHHynfOxb+tqAmtBZiTm2CiACc/6XRYdj9nQy5+y1Z/Nj
io0ur4XzVPvWSI4mEYYnTupS4GK6c1B9G846hGs6euE+L8Wux9DXLkkwsEkIayRzI76cXXk/61e9
/0o3tAhat6GK0H9Dok3dwGrgtGzEpIxlO7QH8hUtKvtwFJzXbjwU1nAdOMTKTE0vTy3aPTDfWyc3
m0+TVZEbMfLjgaZS7ZZnhG+LxyNDZ5kVAhM3Hj5OhzpT2GIcjOttz05ukv7df2CxMe4+GjS6m+ke
2ax9yauSTInnA9G0GuCXfSB2yxqHdQZOzgKfOB22FBtgEYW2t968YZo4vB7BX3WjNO1GfnTdTRHo
P30KEJfpqcMxRVRDO+KsrpOSDpP7CW3v0w7ng1yLbR6EKb3rR0q5Ws0g7KU4gSXPIZz/kP4Oi5bw
oXUFjild5MxAVOfcdlUQtZhxTbgTQDl05vR3koP9Nt84SOU0lV63BWRMXc2j//5ZSrC73mjmpkyj
6sHMe/wAQCSBjmhJTR7434H/RmZ/5zMRjw9YN7B1HDnnDk1nJuZ2GhXbYohWXhHCZmGpGraoPTAM
Qi/7vLyZw6Vtp79vmk/CP7AXm1Id0c7mYxdkPvnvWCWd+KjzCoiU0wZA3js52aG6XBRSSXVFQta2
5G4TRDTwZkpdV4iqoHR+ByCiWSqggz4/6Uoe3DZSOr5VoX6OG9YeT+p7cygd3BTJyVKB2E4iYpsb
g+Qx7PU9721AEEfuaETVLRYfxOfZe6JcMyjHvM44h3iFuoCMNXiZgNDMbAeJrZqUnSq6VYPtoI6r
6zUQ56/foXssAJ+DILYLWfMLqzAGHKrk4mA5ctX9Hy9JySPHddWWqt0yeVvlRZRdeEvzGT+sirYK
hN6J81ixTrR12RzPJoKVG1T8VivSU0npHsm1Zz7Lo5530imWxYoQqYvOtnzLh29gzcDjvqkZQIe8
9jI1noN9brSfAHVNLLKEirUHTaUMwkSjgpTR17AjAnxyZYCzGkEsaAEL0FoJESM9eenpku/ntwmx
ZvJ2jyDkrsTxH750YIRuiqZJwl5wNqqCSw5E0X9Iq6o7vMGyPfHPLL19BHlaTL+fCwwsO0OclnEj
2n/BsDmCTuwv1o3QhLq68YVGyccBZHWlQH6+I52kZpH65Hgj9NAsKbOLxHDOH8QwJvxuGcPdkwX6
lbe0sCG0Ckr//NNKwtW1OPhidMM7hCyv1rlXDg6t4MFR7GJ8pdc+P5WXH9nja7bfhODdCuj2st93
tmJyNgjFoiQL6VipPEh1NKKy09yzZ+4T3wv2kOBGNYZButkdPtD+XNCGrYCz02WHs7GL3ocH9lzX
6L7J6yIyCsicMFnTJDgzLnX+0zEtW4r+wK4VKvWtvFPSQgibEPwfYA82Y8E9rO2PLumoYDjPuIpm
utFY+fCYn5o9EP/S2HBJccuOOyeQKAq2NOjaVU78F3kgj78iooRZNUjHBkZNHal7cjK5V4czQKgX
pqKDMVHv1zpPBS+p69FLU3vSqGAon1MVhT9L7drMlum2smem36l+3jExv1mgevJjrQX+xCM9imf4
EHx6dq0eEyIsOat7gG3n4CgWUL5ck54avNxOHl62nFamFFmD0ezrgjq/5vaOnIzWGgCowpQ/T+5V
yTt22piJfWbklAd1YFvtWXFz91PSs4H/QltINqFHI6Af/JOPDvRc0sygeSjnkn9i4DHEGPMZzCbz
2wOQQU1FXnQHGmo/OFXK7hTfex+TN1OGTw24UhVFw4o/sdQMfCoQyQZC7o+Um9fD2t7z8XwUp/7k
AmJeSHdTqyTdu/085WXKhw1u/AUSQbRgayjDy/0SH9Hedl4AQnyIZ/dHpcYoc57/FRkRpeMsasUV
whXwWQDjHqsZRps/mwDynAqhnZpYPHKCruxd+DYd/vRVN9Bio21SmOx3D80SvIfRpGrTZtu6BtMZ
SZG/cvnFiQpQEAUrjGQLF6LeXWEoNvlVyG0/otR0OdinrOAX0F6lhtaLCCJIJrXI4ZOLK42OVIDK
GaSMxSuzXv9xK847sTaodMgmHbUNMryjA38mghuO89Jy0cmCNviDMdIJHIS+eR5d7+Ws4v4jMs4p
FHu9Vemu/4ZJiw3D8P60hW4tXgMPaXvHbzOjvbPpgavPi41RB45lFMMtrIf+JP9ZZtNycO9sg5tW
TrNY5yvr66qk7c7hqW3lhykKMJpaC77NS9hs+UNZKA2UcpC9lY3n36LeGwwcQPhcfEAckHxVZ8EC
mB05t6bF0UTI2yYLGRCh8TpCV7Cb+OEzEMopJBULKlRkShu9LECQRT2J0KhUT1Ui9TITpmur+ukQ
bfOL3FDguA0X7VBmyI/OxU+/w1XgoivJQwz9awf8oot4HBgtYCollqTX07Kjtfm+GatJCERIE0Zv
lInUhhXZ4emehQi2K2iu6Utq4+CGSfRKZepYtb5G7imonuvXrRHlxwjStndtzBWjOUQUUvXrjIGy
3NCi2vpBGU9jopIHjt8R/BVI6zUU8EYdJ4kI+W3wbTthOz+q8zNvfcfZtCiLrO0tO+cxhLV7bjhL
ifNA+oZWWj+DC7/wNOPvcvlpzpLyHXAYC7hPi+j1cPIBfs3uK5ivsNDJ8kDaf7Jqvpj8ahvwHC1u
+nK8Vw/UnpQeRQkUZdCd5QTU087Z6mMmVNUtFvQpiUVP0YGQNeuun79SBYmZTOJdPmpjkYPk4lai
CVZFzl9x6/B+qVtZV7xbb8dpB9JmLw99UgyhGTeEy34zhOdCTKqGtQUo6RhkU69M0tGrL5Wfg5RO
jHCTTvIJLd4ap8PHXQntweT6oWxybNzD9A51NgNNhpk7PTldvB3C8UYLP65uvZiyXEkqKvJpGD4N
Ui0sYCxNqOJYCrOgekYC4Yf/QnO9gTYV4P1h6QHZsFIbhmr1+uNrwsbllqW55IMHnHJ/YYcfVoCJ
e89VVwDtU6rBVksStTU1iS6zxLYtK7pMFeORDrirphAhZlr0+VQkNej0uYLTdpTRJjbM4nBd0n2U
8o0fz0P5ICqzlBc0HJCdS14UelG0OiKRo00Icb4SdX04ww+BqwsaOxtUcygO96Jt5Z7/klLYEu1n
lI15ZvhW+DWG4DpQFulyNX4SSg6QPFD0CAv/TKLbONgfWfOmvEYM4nIIP8SZbnTiYJ2W3QhBK6OS
QVKlD8brq33KOoblIM9V+e9W3GMadd01TxWN6biav10Bu5GY4yl/9RjR3RBDPJaHyftBfTnpKdJE
+tq8ACw/YVB3da0Je6SGyhDZZQ79R/dNzGs16Q/RrXqxR8tgkUVHRCXee83eeVJK0zhyekxe9U1N
y1Tc4r70NH99Mpo1xbjcWcOKpc81dFodZPfDQPsA+gGftwjnr9wQ68opt98GeoBiUKJ6HeBDAR4o
8f2IMzmY2m8H41hWrvPaqzHyLG3nAz4csa1po0nPqYwqLIP1kU45Nei82QExBfYmoxXYZ+X6d3kx
ItysJ5LPPa22atQlmR8BeKesfJBRIqETMxyFMnDZsvGOqJrzNgWTRVG/ESbc1mqQHKN5IdrjEivp
b6lQ2fl1vwh9c9UCQQu97EBXylhdeuyLajCRse0+ZYsoMYvyjgEAP5zkihZcHPM5U8iI6veDcLhu
zbBzi+QIVS7NM2D9FT8u2If3IfRy19LJsjp6ml81FfJAzoEi1+PKbo9ZcmAz9L2ZWNls9en5D+A2
e7VSczTB4yJNpLygbbN0GasfGsaqmf3r670xrndxLaTW6Q6hhIJGOCgIgEiX7A55hiIIF/kRXhdM
+2anglxeYCLyIaqa4G3Nipbm6Mdyh5yf07/QIxfkb24iUfbKooR7VVUCdUwvmLc19xqx/+UmkNK5
jQltMMhvi2mHUJYd8UdIKDn/SLPaFqdZ7/vXK+8AVNYK+6zrFjKML7YrmekPOs4E1tpR4dZY+N4g
DOQWOlNy13FTk3GuxjGebRRixqtCOElgKi3N5z3oD5bxvcnPI4oyCI6osIcUyE3wFs6mwSeT0Gmv
/KXDRlLk68s4fcA2MnXuucI8QAXtvCEw35NvKnbKp0K7FjimBOt5jG0uLBkaaNJw+EB9dOSMjLCy
7Nm5Yzv6bKPb1MvA1t329/9BTAw/nypLMLhz/GdQ4b/ixdE+UswHMAS2mS4b4UzA1o76QSOHyeNd
UaCT0QUBcRdoQhaUNXCQhv7aai8vRk1uNqJxfojvMWR0M1/3GNJd9kOEmoIQOV/EbBJ9EIV1T51x
c8jaYSe6uG2oEHFsM5urKddnZVYF2e+uynU2sc1kBJjMk6dqB3eOmrX6g3gAJnn59LoLAk4JZMvs
Q9i7LVR5rVc3ueQxQXQjbMvKuHsOQ3YuzyhLecPW3P5WKHwluQglFB5AUwzKECmMsKxGqBtVeM1B
RWb/sSHtceoahy/kpL1yaU/OxtEac8pAQWEDkGr5tHRsR24wj/oetDSqcVf18aId2wGJ4qSpbsul
qZ9zwrJd6C0BNNXwj7+Z/xjcdD/NFypA/x2Lc/3IwlicG4l6WhB2dQjIJHMdT1tuHjsH40RuwTXz
lb0iaKfzL4cql1QHOAMiZbDZHUojrwc6npZ0yHsIKhsrdmmCTQ+BOo1dqyFtLFLStDmMohPXOuSC
w4KIyzE4lM9tjCVjdBdfP8ey6YtF05i5XqRnMstP1PrdoEizXNe236y0KAsRg+8YTWGO5EoUqOzs
IXd/XjHFnzFeALkLpsLgitoZuHv4Wti6NYz/mPZ67itoPACrJpCVH1WTBJMFVJiJRjscyQlVLYk6
2C/Fm5th92/npYC6NwC7Hd+TDC1R0B+R1jAhcGJTkvPtLxJSop8RcBvGhZJwGO2o0Wsk14kx3Clz
uK/WtXV7Y7RNT1V/fInCbzVzhYpvp9tphL/rIvFulL51CPAVtIgWB6SEKsxKob8DcSj1GHTYMwKU
AG7J6F3SihCXm5M5WEh80fYKVACVo6TgrzoTdZfYrDJGcFIceMqC8rPYFvMlujH3hf2dNfcW4lp0
IxLg4tCBP/ejwtWtDtXkox9fboTFLC3u0XKgBR9Pk7C+IGFbIo6FvxrWBwTLS7zZWJy9wiXNHzYg
QHGNrOTNv3Irr1BWbKodZEsws5E/4K9LsdPE9IC811b5MOlwLSPHyWvRywr05UTgy1iAfMzIeNLQ
FPZ4Zs8v1XLURMrw5guqb/+d2aWXEA+QZ1Hg9eKVhctI4bGsw8DC5h5EVdfJeKQnmbz9ZR4Qqmtx
Zum12r8JpTumukXA1AMP8Y0eqY0XAfbGPO4/OikNrd7hthk58Uzz3JYoorcl61q5oP6oLX4WgQgX
UzjlV/umCv1rT0FySh0LsnJ7aarajFeCtDBMGJFMeSsLFyWrYMclKAJ642VgXNWHNwj+NuG54l6U
hVBgPEdriQ5xlFVDk/FKRiNSykBL7Ifb30qcWPfUGDYDenaGpslJMqHlrVxxGOEkdMkl1fu9NiJR
xZHp5/jwmr2FQ8Q5xbb9qRXiEgr3nMuJaYgKjW2McTu2f+g62mUahTgaQRq0JvZ0u0t1InbQa5tH
FEnfL/mGSaYCuLkvp58bSZQDoG5+XOpBCF27z7dCFfq/LcI2X6UFqwnhPwgo9iwd/BRyvu7Ml+s3
LPhcEA0ABeopKRmuYcksiN9veUKvlrqcwKu9yOb7b/imPCWVSOj67xC9EUR1HRzvofAg9zCX4RXE
mOU26B3eLXzV7Dr6KGkB/eIJ2fAAdpeKiV1h+zsjUUBC/6shxhG0tP6Wvf28ilWKofXGPxmluzyq
UBekcY9hEc6SFCg1X9EINu0uoqoTvaCb5a+Gdqj16SkB55NavUty04HpeIyBMi2fTjnLrREqAdXw
MdE2l7hWJViqsUNxMZgW6eZB048W/76+f57eDvDUYf/Dw1fh6LJhIFpsvCD6RTeUD3WHaiEfN4s0
wLkXU80PfqBrz5FoQJRidQQmoY3ftR/yHgQeMCujc68bS+fGiIhO9Kh4UiwuCMqUYiKbzJCf8Ag+
Vk6sphI4rDWWWd5rMoD4tDEsXl3fnh5YtGe7fbJs7I/mwIyr4rD9gvRn5INN4e1tGbUbsm+Xf5UB
dHvEkj++OVy7NA7UO8/z2sJsuKfrYuUEJBWDldlv7XPuknwiI03fmx+wbMwFdErr2/iTLBz73wz0
1BhC3U6l9U2E0bCHxUbP/Mi1NFe4wpxzNxTXKaFQmioAdoR5/L5sJul/rNuH24DWYEflxXRXDDyH
ZasE0Q/CtyfLenRNtwezJMKiKLmRF0mVjdTGkSOwDIzmMfQ1hrc/viI6bscvqyuUg98N0ffT48UA
5uodAC/sbzZn0CxM8eC2cMPsOgVYMsNbrRFVnWNTPbjzFX2x7tjSzvRQyqTELQHnEQCk7lBkoRaq
0QzX0U4bJIFdxbeKDVx028rXKI8USdM6FWMholzWwOFnxZXeOf7Faea6grHd6JnZFxEGdZhW2Juz
Tiai8aiN+FIxJ/oJH5J1WyZy7kSw79zPrGVJF5XV5iA0WctN8J8/X0g8mIoKAqv4WTO8nxBSn3S9
/xBKpBbeBSvawuwnFa23mt0PwswyR/zmUlLVL8nW15269Q+kiNQRQBoxXNUVUBBnnVfQzCBGjN17
Vg+0yYwRpurSZ3lyfB58G5m+Tx45CKT5AUoaJ/LwP9THqQrSyAFnqFbWUIit7v/yjvbVk72iuVd5
59xriFvz+A8pAMi3g5SWHipvzqDKMv7qLA3vDwFMiSwTYEJtxhFm8csCsaG1izaIkwflXlwJDxNv
gh9uDn7eNtLY4iwB8HVKIIxS4Q9kdJHnvlpsUHtw8Z1/CW8Ea4F+bAkeB5Mnz3SOcIO7KYaqUsxk
L1B71RidaTq4vVlcyRx1uwYfAxcDkkRGb0UfJyKb8ZFUHVgpgTO68CTPde1TvdY2mi5BgSyq796k
Few4mYRCpS9MLYtL03vjRLbeOeE+PVaJNLDTFZksAoqlNH6pnCmXuxJDDhvLrc+mkz4iHqvKZ1fw
Ezydcxki51IKNYU9wBBfuITchBQAJHmtqPqbKX/pO8wwrhSCA7houc41qRd1gnNRbNY1+PFO5eYb
K+7JrMl2/dqoxsHko++I1Ci5ksZA3TTlVjYDUH2FhXVpymZJfcVmWdVqKIJIJMth2oTAYLAzjh8S
xRgStDreWDZoyiRtSlCKpM9207fV4q+nlrOaih0U5cHfC9xKL+wEHLlM5PA4YsazG5zJqcGmM2PO
tWc/g37TUeaLoljHPfGi+LHhJnhDPLE1wEfVSFLcwmJOTvGYWSJbnMeryN1sg03ci+keZZpRlq6w
lKoIOihyNydQfWxscZYAjlfhvFVSUCgtSWrCyoLdnOR/7LqrUerPvlkkFduYzoWWEmC0PcSyxydR
AhTnW0Pbjlnjp5F2pMeceQ7fT4auGtGgpxIfXGDZVozvADh7Tz8wRJ8Epk6cB2LfVayRfNN19cxA
CdCFYcG6klxMHy4YpogsnOTPQbNkdQWdrfzBisOMpC1GRhuu5boR3WwuhkOS3rQKIv9AtGs6PmoS
jDYvsUD10Z2wZ5af5Gy/fuKrzqm/ywKKvorW42Iw2Uo84QbWbZ2y4pMtMVwYFC36JPiaTHysgvJf
LMcwPtmtVYfNgefz7795NSYf5sSSHrcpHfJ0d0T7Xk682L++0CoRvWUYWDdCS6hngIJCUVCvNAdQ
Xx/lGw6qBVcnbUhyTZL7MWakNupCikdqU9miQ4DKfr8/HFGrApcE2oVRDPi3IdNpZwVkHtxgOaKh
kJGR61ovMtQ9erGqW58Pzlx40qgARluVo8OEXsrQBt8i1Z2EAST3cEcPlLSY6fYrQ6MQWAfbofPG
tnVgy7bJKk5LlKLIiFGPLU/Kdht8PfcAYxc0+LzIsXv9ln11m9aRq5CWxeD2jmlAlubI+GM4kAu7
h0hjwbfgfA7Tg8Lq8Mz4C0WHvUXwfYXfRO/7vZleNW+qdovJ9iIoQoiJdqO84ZJ2TmAan2GIwXit
IjddTt41F8xPVu2SpFf+VFm05m5C/rZG08a5jfBf+U3pUvN0vo+H2de6VWwUcaogUAenn14QDdDl
convnHghqlVO8J2ibwQeERqOVWDf/Dnko8dJ5a1c8pDZs+CQQYLLOEiOJ2gq0xCxhRuv3g5U2JVD
fVjoxOyA8JAiNgT/kD4G88v1pHfHPxm6lANC2Cz93xDrBl6A/JNdSzqHhSJnhngA8xtdLuoFKX7g
IatEHO5i411Qhci4PRjbb2mRvqJRHLSJsE0hvtvB2xMKkPYMgrQyLLzxR43YjqWA6ri7dwd95/fD
ZV9WPf/V1azn44K1P6XSEQJ7Nj9Kn+N8SfozC6zPT+lCVHrHFmCPtYVSXxFfMgnkB2X84IbBw5bn
4562ht4GfRKiu6y6s0d2Gbc/uINr8HI0vPg5qmBwNysDMjmMWNeiG3UBzM+9g9NT6TjH2Zi9E78g
VWiIDmeic20OaUHuas2KFL/IAfay+8yu3axDaguK+O2RL1UQfpCGaxkxCIlrW81Q3tisD4F+/Qon
0zthPkpNu3cFjq+HMocInKzxoiTztgfc2rz672ngqMoDIaBVYlCmql9q6GolmeJ/K7+90fTQmV1H
QIeJI5j5eHm0tU02GNz5jPVzRihftuUPr4sWSnyhhTFC+NVMFHxCn3ibS79mTEIf81jx0Z1YkBc+
SrXhx5KqdyDKAQh/Ap4vd5neDywi5e+in9Ll9YHmrEbtayeQfjRvg/UEuusd1AwIPbcxiWfhqEPI
IYYuMZEwXBEVKGfZEaR1PhgcuQL7KCe0YufdtnTjfVT2CCbVD8DM8vKlMGUbbDU4Sk4lMik3rWyg
1OhHLSp+0J9DvYliqSa93eQ1KMIe2silcMkoOthdhM5rDPeAFxpxX+DYTVv8DoAXLnfIu55sSxKY
OXAlbacgDyt2FG251qqLZbl5es6j1tyFwFHx3l6xway7z+EnPptYw5b9rxzALIygnyTHfmNlsNei
pQUJdLUWHyQU3VqH01/h1tDrtE4A+ZMlwQSyxRciXLD1piQp5T3KjuQWxBfN7gDAsJmiY4JThktb
uAoitxkwAUNQhyimNWMbFtKTngm9PCd5yMaAZaWAa7Qle1JgX4tiyBQMq7mFt7ahzmUlnGq20wuT
YnL2NscWXQL9vbgMWDthPLsKImmPJYlvgZhvC8t3v03KwXdsjrCUyNNLR70tYYBHQgmDYKRKZnns
PnneD3Iwt0jMxSrHYeg2ZLHGamc8g2jp8bKaut1XMxBk2UZDjvvEr2OXvtp7+1h8gAsTOsg/qqDC
otXrKuadddmcZlt09XJ++FpoJyuxnOtjCZCnnYGHYKzh4OChbCraU55E1ToJKOTpHoQG6k0BeWDo
Lu6IM0RdXFgCe4Vqf/iy8oJjtwGSM0ERs1fMYjlt2mkIyAOUYFMMaU/a86i885eM/xUGVE1pBVFm
46PFsaE/1zK/ARRvbdL2Ar4MtEu5RjdfmJ0yIJgUyREUTKmjxW93IoYWdaTP8a+EBmOgEV1VVaJL
8fE/vUy1/+WdHJGsDuXp5WGNW+NA10mAfyF9FDbFyLMvErtho+uo0huybbtdEPiZ1hHSVYJgqsr3
Gffctcd4DEz69Ut6HzJdKuKjVluaW7IgYnpATH22RDhTUkRQPaOGhIVfOD8G6m31PWy36F+/QwLD
13oiu43ydJxG7p6AEUGv4y9EccXFa89DSzcl2AoEBm0p73ZtLD5fbUFlXy2X7t/BE5W+HDwuWh5E
akfCte+UrRBntm0A5ya/w+dQU+pG3D9YS8l7fOEy0nmLug7C3JkmaXxSioTKF3H3BaZDu9UMQFGw
HTzRASqdx9L81uMzEBHc60shbD87XzfUJuhtUKU9nSkPl9TJXqP2gB2twZlsk3vRvoa4HkcJR9fL
dq+ezuy0rmYiwNYkBnEGfaZlQNQxYidLv5zAYQAUuiT8lugU0lmZ7PW2vas798hLQ0ZNbV832DzO
XvfYZRyjpAgzhPCuookv6YTX3gUxVnmMm8SHBnMUb3L3ZqxRKNCgNEC9lHneu+CIzPYEaPnutyK7
jyRUyY4JIGFkkq7w/525OusKy2NAPuR0Bwqvdt6gfFXbSg7hwYQg5JAqj/+wCUBeT0Z4tAgi/0ff
wVtB6uqqZ5iCjXSzEtmX28t/Fn920Co6SY65MK8kagDS1OHhI2e9bt2ccwkvYRZXjljTkQ0/3ESp
6JmBWesaoLIDCRS09exGlYDR4QDaDnKMAWJKvk0DgDusCzygvbJssD4FpIaOWQ+T0LqCVYhEl8pz
hoW1UMlJmkRF/d6gYYBRcAh4xWGrqi5W0j+1JvxPufrT8esNTSrsDm/2+fpoILHaQfJo3NendODA
dA9P6hghQYzmqCnZTAKfITbUMbmbibo6gONKMZUnJZv2ECJMz6o01TB/UWDReCZw2yWfz2shElKG
hgoKjPItvywVaNnGWkk4rsxqyWzyM8GS/GjWPT4A2fgDyzLoelOzSq1cpHjoPNUEb9FKMFZvYtBj
rBoYZIYYafuDPqRZ+JSAT4GXA7MP9JAjOIIDMmD99OFiEULOM/1oOU99gwBVHR83sNEvkqiZZxK5
GJXwti5Ckwy+G84yvlCdIoY7tpVoIEGHc8LNqdoBxuW19+i5vgs2eOAcGr+uxb95L8zNgZGfr0DU
Lz8m79BH3ZWgiU8xMvtpQLeQy4NVQjY40rk9EBa3HNzxv2QIbDBuC7ZpDfzz60sDB3WJgiusCbLQ
trTiaKP8gruZb/yiCaY1ZZzjgLTOSpZ/s0ydoDBd7d1bnjzLHFeAzQq8N9XaUZXHqfEbodJ9fZ8n
2hYhwjPDm2+/TpOJ6uSHXdz08ecRsSrPsNv6JhiGCajjdQKLLX6rt0WwuZHhMTl/vGmBm8vtOqJQ
e6AS7bUIAx12AFuZKfZBNfVP1K30KoKH+YFw8e5SXkY4XTlfwXK5SIG/2JD8jUtPE7H/vyiVqbji
rYTsuR/5dbB5b+QKYaV/YYUTx5ndbHEgxOMK+lZMEuZrC4jOTSxOLm4lvO3eLa1Y5a5eSxbmmEzb
LyTimytJ+Df8PaKktXGd9t2eHpziiE4mKKwbNEyrK3+eis8jO+OHO0MWqPYEr/uTnBfg56YlJWy4
huFWxhuiaH6QP4ESaB7nQLB8KUYW2oBGGQ53d2HftdjWeOJjr48WpQ+isYh3mpkxrbhTIZ/GWcQn
0j+syQFNG7nF3Ay3mud+KjDJnwlFKMlZy1uf8AUPfDSuJnHNXfDqYbpoDnqkLbRpvlqMyzcvH6ke
ZDEsalxloxc2q3nDwbSuoT9KmIFpLou2cAr+qIGZ9UkqXgxnMFHqM+uhAwX1X5s9hfMLtlE2Y+UD
QDIFiIll9yjFKwPYL9TvPvajkCytaTfE9rss8JSyaZuIK8JpXQDPfjvNFdwNtzgnPFydu4ROJBJO
t4WcDkcI0i418RmksXtttZSB/bt+OMVhTnagLdDS6g29yJcqR1siwuzNBnROCWFYjEk3hNnImma0
y1mynffqJGzWAuiaBAHbxZ3TowX1F401Env+Qt2FIxq2DkA1RV5dxD/GDw0Vbi9KNxWxdz9pDBZG
XGvF8qj0kyh4ztoshTdgGsKeaCLrEjYLRynKfgHWmzP4YSPgS337zssEHR6DdYQYwcgLyVu/RLQ2
9dJ7BfntIJlxaVL/ghUL+oAgzcZ7wIqodTawBkEzfYcrtWG2H56mx4w0M+YiUm249FN/EXPsiIby
4MKM06+fzNhIqvwGqUR7MQg9QOIXcASPoVjTSCEKXST5JT31YoAOUHdtHezw8uMwhSdKD+zxkn3L
m5k9LF2F4XBkb88y2r3ifiayhZx7lcpn88eReDfLfNZQFQYKGAn/pWosZRYytagGLtKJnkojnuV9
LkPc4n7bYjj9UwcaeVQi4dDm2mx9uD+N1RwbBOfhIm/DvQvFs8hYaCJUtmRLu9ya/pyw0njMYK8s
88ELmnJWUXFUs4ZU01TtaJu4UQ6eqXNAs5LaH+MCdVCVMkbXVefnsnr8YXaWtoaYQdqdOJo/Cdyw
7M1dAY40YuxirFgU92uL6oG8M3+0gAcYvLkFTtM5SJ04AByaWTIWKuKYDQXtkmn4s1v5tj1zzkF7
pIGJ4DUR7CLPM/55gd0HSBvt9YkNKZ9/uDBwr5ctND+eG/JGDqtmcm/gIMrOz1nzJqA/zjEqbAWG
1LDhU8+ubNoB31Melf95rKLlAOLLR9VCARqDke/X3TYIHlQdDETQWF/XjAfZ0R5zhGEcYokgrxwt
v1gEZ2npuxnZpsZ3wuNTbp0/eZtYSsNS9jOHNLiiUtGK7kSnZSWJ42MjipTyt5ojvXSptFFinY4R
1Gl8EupBswoyUcDEMyPVjYCnd7vo9xXOmNsnIuaxWV1TjU/uoub+mO4Znx0dgyc3sNoS1REkcb/f
rzG+r1fJ6vHVocI+9a3HXWEdPAewf4Q/6D3dyl5opDCr4aTUE/9Zt0zjmMXXxXeNM+wA0cfyT4XW
vUwNqsTPAETEsq5w5WnL20UNc0q5dKskxCA5Q4sDe6+3K2k2XJLs5eteZLoqfp+4CtTmyj8SOpTr
eiLOnXtr4vU9Z/sdAL38EEtxUV5QxwOpd3ykFTT1EK/YsHZXSAn4hvWpu+bwubUvrtJJuoQurLAk
mtpt4evO5tzQqra4uLCM326Plv7AVLVsEwRiXBx0jYkE3E+NXgzhjQ10YpHBPRVZ439RC5xLx+l4
T2qkVt3yeNNE9GRYal4TsiwGq285ofBcV0py0Gm5qQdaujqtAPmARmVD3VeOFWX1rP4qUJskPaUj
MkqKMyNDjXdYpq95od0uQC8O+zWRvme+4kBbErDegcVBbN2j9486WvvsbkS+3SyQ7mld6llADVYk
Rx92+hRORWn89tlkxNwlRnqtHbsfOvoWckxZ2OD6rrsDZvPG/B0USuF7bh4OG4w0/9rL/vkFMr13
nyIUiV2GIcZ7t+G1fC+5YABNmzx9uSeLJhy6rsuOZVAO4nRu9ic0RB+Dj8/L2clVh3aTT9ZlMqQk
B55BryXF1PVRxlVyafiAPV8Uj1JQMDsXR0ciUS2+GGh4aUG1YisFORdKNt+SXZ4IkmDa0mP3zK4A
Xf3CCJxMmCEHqC2PXdSNoenqAEwe9GeR9oqQxaJfaHdyAC/oYNgRR2DF93JizoaGfZrDLDhjcXs2
qImvU22b949v3TPVdwWhGjJrdwhOPWE2mjB+aeXC2WqkjL2/sjGDp8WCjX9md7zTXyO2+znx7rPM
JzlTKsjLHSSrXo/n4dUwWxK01h/kZQ/G6ihoT9hAFrl6JQnsoud2/zx311ma5kDMWW3IjWB7SSp9
ZRQnlZ/aW52h5VI0hqIjmoQSPbnl4WNuLykc5YidyUUu4q/1tDTTefT+WKLvCbajIZG5FB0aSPde
NCt4wTEZ3ON3ciLT8mT7rqpOFxxkK9U4I8u7filfVx0MD/SkCXpoTKgziRT8kL9J+o2Aquj2HtC/
sFUh8eUNM+16eHgc0DNwndR/3bL9PqLiIWClSMjU6Dw83ADQtmHxS6kp7FnMQbrR+5nLHTIilVvQ
NX+63SF9y3naTncyPSok1NskllaPAXN/J76H2bJxe6klxLQ4z8E6ppOESYLxW9dgclJwjPFhaIrD
ixrAGrxrCivz8fOHNnicOKJEhomVtCWZPG8Q47Pw6N3nHIdfoH3x4lH8z1hiSp2+Cw9zxv1NOI6Q
DEdJwzEnITI338rDoq4kc14YHT0aMvhnbGfvylA/1y/zteJaXPNEWiAlH1PbVOHxpPUtCoDDey9M
WZS/+Yz9K/P/kRZ7NZZOy14st+e3TqU5R5HOqx2AknSnPDjWoPL47BuRJ6GiOjRK6jQCbVMkBGAc
qdgzqiN317KgJJ7JLEtN3U/OpKjLz5/ODoBsvOo1HvDgrA7eu8i7QCDYxqHWqbbKTsBr4xikK/7n
w0kCEaZBrZJQHq0eWFimNEQqgXDJxS0HlUYysoMeNJeYUbL8xGznT5nv5gsh2h6RmgAsPxvNk/+V
ZI8aS38jM5nQ1mucjGG6aBT6TP+c0Io/s9Xz+pjsNY/OfrP5vGN5Z0vERa4jldzXRTAWwruyCXxI
/j2vQ7N8PnoPWCfscEZfp5cBTn1sp8GsZrX9HKQJzGc+cOhQp5SDVl3MKgXIHaQb4/1KoJkg3prU
uQ7/hDNUHc9FwTJdfc9OUdFbTpRvj3VarmK5iEo3DE/I5oY4ol3fVMRq7yMe1J9jYXbbHGTbzdOH
XV7tq1tVKeUubrttJya4vym+S/vkGuBZkPi9nwU0oqQgTMCfCBB1Y5oBGd77Wt1CXARAikCVIK6f
zN0iEGT8KVClEIuDCeScoA0DbhSTYseAWS8XVoEYWQ3VO4N92GYiiBv7Hgrn26wE6I3qVn+YJa6+
iihVyOH8peiP80yD3VztwroknuhaVO9XDjG3G9OVuoMOZ+IcJ9ORTUYhiNFqcifktloU+0nK4/Mr
YQ/QKFG5SDPACmywByKnXRrffQ0RXfmFWthqv77MUdmUbxt+gRvqkmd/S2H8nAJ3lNxsqOfYqqTz
QiDIaIst6CP/bUTeZIUQ6dNU1kaf1CHsXKJWP23NX4HTomdlPhRDxFB+hHOda+zLi8mitqjI82Cz
sJkN+yOUYAOyn0JWpcP2LMt1tR9wzOn/YQRn0LKMtJ0w4xYFkOpmp27ZeTyq71ao9lBOddyOgPvh
NLDNHMdTqdRd1PKHsmSh7IlCKmRgjbf1QlVwP5xnbL0meyIPeCMHP3MZWvjwqfWs6i4wrBzooLYR
NKANi26M5SEYkIBXe8Ujf8c8QrQIzDa/YewFKRGvhGEPnrlVZ7R0wbmV6zihlhtLO+QBhfEA7kFP
w/1eOEtHxEwm/o6iLadxebOUvTIa1hX7zrBzqoqKgetAgI8ej1T58DsC7/YQLyiGzz5DPADgELXO
1QNp7EhG/2FN/ywIPz57oG2s2MEcdmohQnR9DUoSO4o2dUpv/IeBRcbVC1naFx36mZej84T7cwDY
MFG6HVG6OHeP4PDvvdybURPJ0eduinmjbLG+zRj7RcKRI1+INTATeBPGjXVXLmTujELLnUaUArkc
SFnzgMOGnvD/sMrCT62GxFXy6sBOCE+4wdvhSEJGF0Bi3LQqsgVM1jWuzf0/BT8CA6l2seiuNDcG
OPw4Y361n1KzYKsZ8R9c67RFPNRlLkIaforLq7x9mqEDDXFc5CYYvX+ZNnkun5TtI3dulYl9IaCM
P+1ubUCeM7j/1rhVskXelEreZjMiGS+p3LICZeurHnvCUTr5fQojf0s0HM1OuZ04Njdavh9WWNr+
5Ep8DpoyX0+zsdLNxZL2Xz+dISvZSZ8+NmnIUfZpvydauWZsscML1nWt/Ent9B1WUp8oi6r6MMVg
1vwJh0bdtTwjLaxbF/sQUs0lNYv5Bg+hyD6Npy8GByntQbl7/bvex/va5MfM8d93hIajf+5VGDbN
CsV8aQs5sPg3ZS6wwvjAHTFwxqzJ0EXrZo85PhdLq7tc7aje3PoW45KY1mD68+DcHgUQ565APCfF
+b9e5gg3mPP83V+UIJMIfTXxpAJFIXyCU+lMxaW7HKPFi+L79loylDmItDivxuePWGvAPeoiPzyT
8PS6ZKZavhpjkhrSQ8bqniv6abmM4rRn/FtnEde+lUsooxDCKxQxUujGQimvQr8/ofB+HZoXXfA6
maBDtVKgSehIbr+ctSfTNcVTORCbkMbzybFsvPmfTR8dhN+uTFHKbz5cbbb1e+SLxsAyYIm40mWJ
qEpH5w7Tx3qMkovBLnlFRoKxJ0qX5hEajC7ExWvP5GttMxY6HVkeiyV8M4tS5RK6WjBMnfEG2yBg
H5TPOs7uDdqPgEd2YTVaFndiOHUM5ouiG3W1IcmzPlnT7I4wBjpX69q3Uumbj6gXJK+u9yLR4D8q
ZVsi5b/F7NMAaPIDzWj8XO7zq6otxkHF4oPbhcPi4/mjz9rVCLbUj20zLjTs61/FBOsQH8fQImzr
J2m4GfVtqJAEQY0dUC4yVsKnXJxNeplGcTSKLmytzfAOYP9g8qIebGOSqA/J1l6mYylp85+Vwph0
8TOdbpdleKAMxzs1m7S7jgqFr+g7olIACn3TXJzw1gGHyPb1b2FQiaXo7KphqCruK0IcpahYUp/Q
d/vMlbxNbzFB74JEJhov9llWKPQS899oBqrDW/v5f3GsS0PoXLvmF8XxLOgMN08YQpwAL5T5h4jc
zjyiZmD9GmUfr8GpJsNRqQE0STN0SJrXu+vjCbiSBP2NTQFXQw+PWZg52lUwksrRW0zq8DBxTIIA
JOmMLKq1QRJq75MuRzqSzS5+B1dwNOeU0i1xQQS4m9ItBq9n5OkunlWHWYN/S97vMzNtix5ZS2gM
wuD38WtWiC8xt9NKUQZgsIlbBWKwSZKgxwYYR4vEL5q4IaZH66v0wTFHPlUgeE7n419tXojSFmGW
QXEydib9zfk9aBz4qyd2w1IIwaMHx/qmXBFQOn7Zp9uE7lIqZUesnnzpeeZXjrx/LIwNv8PlYQH7
vfjca+evDcJXamaNiwK88cmNTwUHu1xjYg7mWs52Ht6ewMQIsCWOoC8HBTVraYOjxmH7+zfC27rn
LvSKl5yca/BMKv78ynclMR97e2+7qhICbOEGHQNljUgdEKrqXuu+DkrQAnRXOCbfvdX3Izs5CYd8
TFZTXRDYmeN/Oh5Qn+tbqFySij2eKJPVmZy366Ap4rb71N6xJ6mBNjmacgTkNQkOurduquusfQ8c
t83BwYrwDCzIiKzAmHqlYTHNTN4pdQ0hVg/YHtGl3CVGrM4tQvJldXpH5gLS+7zKWDzjmC/tTvf6
YFE/aXSDKXnwp2T/YGS/masK/yskaSYc+0Bt+FNGXnYj8yWpOeMGIJJ/Z4XMQHZ4sVJBMqIikS3W
K1rf+uJN3/ZXp+kX+rxBQzMPQwsvnieb9YJyTeCh8hkwgswYsVCT/6Cv7SEkzsc86oaEfjJjKzhR
nmFL0/gT0nffarV+vYj0ZUU0Pkynz4ye3qQpsn90CUZgecqJVKk0Sb3WJQiQjVw6ErboYVg44eMg
xS80wKePz0NUKgoPgkkaY89UzYUH9/D5UdsMTDfRf2RevnoEGNhjbd4X2wvyCqyWwju8VQ6eMFkx
o2YajFCD0sLVkCshmRKjKx6HRPKTF7voo+2MJVyk6/YQHJQ0kLNGyosNr6TMwxXdGmDaSPYG9NcK
zsJ5GsaRvPD5dJ3HlSWwnRxacx2eRIWHFR5Lc5OJ2DbvoXP5VH2WpEArDofw6y7WF/A4bFA/RZFb
/CUwSiCza3RLhmK2bTU1VulNbLfc9SoEtNOcuzlLJc0b2Ux06dPKWhzB3Y9Y6zODTAl3Pc3QK1FR
KE1Z9PV7o3acaaWNUURBe4CqT8GB2TB5fgqF4toQTv4esjRDBQD8Py/uBOusn4tV/xYQ5d04kaEh
DfY/GmqmJG4ZhVVbOTBl/D93Cnu/d1VAJSpjcJaQddYAqq1ILCw46yCsvfE85fkEU/QeCA7fEtkB
Ep7Av/7XrvThoWI2TAbVMXp54x2GioiJ+GQqtjsR35k8SStMXqjYECMvO8GIKnSx9QINvrAlo0vG
70CSDNiMp7nDLyd5Tcow0uOUW++KQnd8SCQrztzDxktj50Ymb06BEcuKThTSs/PweviTOXZjSDS/
QgnQMHFGFAwfNJjSueAtFEAIhKGaomajcwmzRy66T/1qzOiihrJSgx/i/sjQM+s357GpX7ga2c/y
pRf/HxBfa4EYPegHNWy1+OPBUz9p/Q8ilpDmhNi04sKHOSrWhyBgm6WkgZOJVBdZNVjFD5rhqx/M
NgwlAmGStEV6RLMIC1dQxNOd+9KwkaEXdDLhQGMUxUdj8Sn/146GSRLy9VZTpWS7VxmL4IgDdCkH
PimIdflAAqhT8RZLmSeOFKgBojgZjqdiE/TiSGuYZDFVwBq6I70YQLxYa56aV+EZvgiv6RhHnuPH
Nlf3lGoAYHoZkET1T/naewULutCNcIhX5oNM6f2OwvqCSbsboQkdKYKxdR1CooFzs13l7aO8wzG8
sVkf0jvTOmjdND3G0AXeVqDSKyIbNfo4dU1Q9UKvseLM/UlBX3hmhjpSYeQZosNjY+cAHlShJE2D
ThVn1F8TnKQTSXNlCpvMpSIpaVsvW0pi5ThlIaSERgiuktMt+iuIxdUxi/t82N2ERwFCYV5TTaxJ
aqN0HgDmQyZNHLVnFGLx0fc5UpL9YIB22LR1OCWZbv8EiPxgbbgnE81k2P47gO+S9Nf9OLlDoPiM
+0QuXwv09owjhM84sLwgVg1alSCHIQDatuNUA/FacZoh85P7BJIjV6iILWO+vLdwUer0pzH9BwsN
TYYBnrcLTTR9oc9DSMvMlDO2vs5NzmpAbyLkBjP5/v/QeNz6YCo3Y8W8nhD8yVkI7ZNQOdJhjEJF
Vw41z2mqx7TF376OZbVEKNidC0iXKBRh+QD6KXm74WAlYe0fptuUcil29hcQb+8EzOs69tx+5D0R
DMipeAydPpghDdZh1Z+qDomWB5WPXO3rXjrKWhUIBu0VfBvWm31rdJBkNOzUOtdEELsWrGuEWIib
/9LJB5BvVpynld7vwl9FZwZx/COvO4fatq8i9Sbd8JPavM0LRo+msyiKyu6mL4zvjNLhXCS8POrV
2tAEON97IJPIsh6RM6rhACp4EVBctaoHBi7psrK2G8YLMNtSKqmBkcF2h70vSod9Eoyue/z7KEjp
lauS16ZDJaSEPJSYvqQl3RkozrajjbjbcMZLuDBvtUpe4gHF9z3faY9aFA3z6YFflRZeO6Wv/564
9bihJ0D561bVcDJlrysEfDMCtyusM4+5kFCVT/SiaNFGJ03hQ3BUvKW3s8aove8McbX/OQi6dKg3
IrvO9d/I1gcPuJdvDHTvdwZC8Psi75kfen5Qr/WMGlpBz6mHbyTwum6yqUhwY0hwspe6iIUIxn4J
gbiCpSD6DFET5PUl266v+3wR92NBFsJuf0jY1qaDYf/K3JUQwFOIq3Z+fD1mLlcZoBppKChvOLVb
zSyszLBDysG1f9OaFIhekyBtPMUllnGpkpaAffUwFe0urx8C2M8Rpgxp0s0x78huoGlr0uWIfDTJ
h3GsaTQl1Lb4pbM8cVazaghXX24XJwvLanvR2oY4islcwZYlZep98omM48AqqLxB62w1KF+yKRoT
Nj3XR3l5RJwhc9J4IsAXEshU573MtxqRMw4M7brJLrgI377XZoy6cJM50LswTpb6QlS8/HR+z6eO
yCinuef1daP2Hd5HTQKs1aZd6eN3IXOJgK/CkdiY8hoyB1cWIKvlEVyz6W8Gh/YGaxTKxxHWIYRl
KAxglPECePsHy2/5SQRt+s8J8RI0k1oQ8mZ1jNmf7dT1azSXVuNQ+s2lAdr7QZibTJVECZU9br78
GdBEhQFXQ8af/Ki0d70NGw1Kx3GbUmQiGs5Zj4k3rFWkF9wzb3RVIpXiGwxGNGCtAsuw0AfjlJvK
vnN82sk8KLGumajyoDm+JQfy/QZ+PnH0VDxDWdjK8/X2jWGAgA/t9npvx5m2tN419IHbfDnFcQhy
+54+fGolNwz66j8x8UVYGl8y5p4sat8MbzDAopBvGg8dwcWytsihXNPyHXCKobj4HJRwWJroUnXf
9JA0VctDmDTk8Ib1eT93l5LV3fZol/2TjgPIS9T9n/V4vpA5SiSYokO36VWgUT/uDaN/ux5530Zh
1ivKa/FeXG0LlAR9iKt8/oriPhjM0BU8zPYwPLAcYS5aFSyOGl9Wg70kBDPqdYA2iBAAsjec+fw9
NxqcBWGS4nDQswiQ8dD5R4eqKVGeur7sJRo10kArNoo9fGdzaJvoxIFJx37fQ4HtaQ4IxW1zYmOn
zwGIShyYVxVZA4Mo5knKXjvFeYtAnYqsn8CU0JZZV+OLxstmTu5wVAxA28iFhWJWFadtwky+x5Z6
xYg6ZDkfO5afPSbJ0ovG4Ruj0abjj9Edt9+yGpqYcuiHHlvDaZ+qhtAMd1sZaeymlu46bqM8e+bX
byvR6atcXnAYEtDU9pA88Sq2mV4mw15Wi1uuGXteAlY0NZVtVwdsk+Sp9B2+54xbVL3B9ndDqNtl
BVuLW50UlM5XJ0xdhJ3l4HUXD6Wgfw3chepGWWk5etiQ/aLMq8f520dgE1Oiotbyq5SfLqiQtIc8
vEUhsuK3Kidzis6ILHjKPjES30Kz4ISAlq/zWq+VHJh8zKemC55FHcC2TbI9mrL0CF31A1m2ZT9p
ur/rcINaOQceuwnxjkrfRkIVe38JlS+djgmJyOJODOEkn2nIGsUAAl3+udzTpgTALBeg93gFdbDJ
FSOGkS7jnfX/ruH4WQKNoj+Fw4dyFhJCXL05cwtMU0U71J5j4i9ROUiqAsG/KFg2UYSyb8uvO4D4
AU+hrUQUhaQWqyH2FRi8/AZ7t8GekP3E+6CK/pyk4mlQI42gPL3pFYcWymS+QGsIG+oIGWBva+a0
8E3o5Ya3YULTzZsC1CobgMG9YqWsm+N02kW+TDVZ9FhqF1/kB+BMtbST2CPN94qDm8WTH4lP8I/Y
l3xYFm1da7SVE/c6dJY8GZZOovaTP6RhYdyRnL3OxTduexFbVnzkxEEAlEWcjHtzzlHFe7+sjFnw
/gcKrfI2oieA0caa1C7QZBvdbhJUp4nuFywb6HU1Z1HAYsNsuwIG7aVYawf6tEdX/59SRBGoLeS/
y+5cdCDwfDeee7qpqgOjkSOwLqgcuo0mPBIEO2rp3qcAgUEWnCM+XrlA+AddqUjuYw7i1HWJWMT2
Yh4NfgOyAaUFkYE+9u0zEoC94zfRHJ3K8Ghp5pCGXdGMEtCz6cW+mZjkXoazdXAsQ+BN1l99TTAs
oivKSenx0+wbF8dijs3arK8ZLnEfSEoFje/JhT2LOFklwcFaO61Ba7Z1vwdtOPYBO7bASiWEc6FU
/Vbs8cn4wwiLBtspdEcTTNz+KHj7dlFB9snC4xsQOxxpSyXOMbKGfOUDAk4FYRnXmmzbnhJIIE+n
B5hVX/0yIjkelMb/2XPcqz1+FESn6RcdCUpQ2RxJ+YJ9GoLsSvq+ndWVszG888LYKrJu6zkRHTk1
8dJSdhUlSfQ7vc/vHHHs+WzCTtsGAAs5+8glwJ3H5zSGiPGadsngJvnR6uN4UhVg2J/LpdMHja8T
MuIQeHQE25EqRK5afOCHEqQRrHhaPyxBhSxZXnvOkF/O4NvkTkf4+iQ9jEkBkipqs+6lGEJanxYj
jgsBRd3Dbr7V7LEWgKmSmVpRK2T042vF6dUEOKGR7FgIUgwn70nmsQdqow6RHB7GbdANNtFi8GWT
nmFZC/pgSYR9rVmRECmqXn8HipbMfmFpfd07PWf4sL+GUMyPvKlTACBAT6Cg8oJYfmS5lgP7lAu9
+AbxEY8lMIgonpkTnWkEHuyGAr2Dk/BM9emcGDD/xQmueivxp5PfqG2SukR06UdSo+mGObzEXmGE
mrXq+Du3ZBVqp6JSyc++4GDP4Uyzel2AlnqLHwxMxn0WXMzxSEVaHKrSmr2q9THn3Hvav4gC8e8T
gZNB81QA3t6LMPuYFXuemQYNOyygTaVtHYZNLfk2LmZ9yMuB9oG2OSVjotna6UFfCjUB0NW7bmML
KVwmKpQcU0xJtti1yVYuxrmeEaPDEfWE3nE53UQx2sF95mCdIVE6F8UMK2MqJ54b9S/cuDdmjBir
lHaLgjSIvL1Fzy5fQDMqcBh0RyNu9LORUBupPdfo9Bk1wbEGolvK+HfCdoa6j2PjkMargDO4rkT+
Z04JYcOyVvXc5Yt/GirxLL+3jN6nCIcGvQFckGapSfUlgjIlDrk2qfyyXsnvGl8imcNNTXlj7Ck8
j7aS52mEwl8aPDyyC/NjC5Zd6cwHbgsgTn2/yNE+4+OUbXKJZx1C0AmedxqyhBM0jleIF+z3aZtn
1GQswax5pgsKAkc2FWQXAfN+mBF6dE/sSs6lyZqq+hQLp6Efhkjj7P3ihlOEB1ksXym/1qoxWw2K
a6jV4vxzg6CG6UF2/v5f44XMsk/OAydrbnr0VqhkOMzqti3ekElabY5m1YJ8e0cHyeSHx8zKmHdi
iSrHFu15Mhcl3X0UUQC/CzLM/FKHnh2hT9MBiS/TaX8qZ97JTrWHl3zaVJ6yG8eBIPxPdltCvFXQ
x46jWa+2l6BJtquwgtOH2DyhMP8BsvzKClB0WYwue84SZ4R8C6YCuZ2zRKzSFtdndpDPUla5fQoB
dNjq7YBMzea34bl5kWJv4TJkvyp9w1RA5kcobSVWz1OMIVzMQ6SoldH47w0VnqRv9cpaRIIVopcG
VTgzihLSUbqyJiE9/rEj7IY7lUuNTrTg5ZCSgoDAa8jWGbXTJoYu9d27y8B79n7BY8Ax2seOi3Ni
VGhWxZepHh60wDTIJnsmJYC8EcFpZ6we6c7xJnmMdMKGakxLiZ6Qnmdzxq/canIhEOSL0aYMZz+M
h3ZyYQGJHTleIejdl1NMXIIJ3fcHJ9DpYeAbE+RYgGX0PUimp2SaqlExcEgrSURjhqoljCWRp2qk
M5gkg5Ww7TGk0z7SdG4RlEKCyxFhQNq0fA4ULXau+Iiae9ZnUlHegiG8xJaIA7m4rInvn/RHZPff
F8dIupD14brKTGPvNgcxWWWbaY6L8G3X3OZtxjbRqBe1ehm0dInbj6WFsVKjpgvvvXpdl8LerFUY
JTvhzNZBA+QEtBuaHqTWhDah55oLRzROv3lUkEbBYJkcgud2PESDOEVSGJxk8DvScaW7D0ok1ERY
Dp16zc5AZ7OpzkxHAb0Fsy/M1tr7amjqPeclp1chV+g19xl01AAk4o/j7b3+HsvD1KtR9p48czDK
cDF30w71H8AaXhpL7qtZwxpARLOurqT5m+KUVT9np2u033neK0JTATPvzU19C/EaDu8Syqjxeytb
vFDpdzCI8OCe3eVzj/Qp7o95ECJWXvlG9YnVlx96ePt1pwKfIS3bAgfjQSZLHEzURiX47XfcTvcL
ozQpqBAj1T4jILqUTx5Qj/T3grPV88TQip3YBBLcw9MijXZOJtLrYLFgByMIwQzY1/ZReanapT+A
YmTKBqS1B/dkDfpolvnl3eJFsdz4dQGOBfq5dt+HAdT2frIDhavz7KscInyghlA1g58W9kYd67TO
PIcMQpaI9PgGSm3m3bx6HBwvOjg1JNddnJPJdAjmBiiIqghgfu2917JdsXyadwVV4fGBJgDRf8T4
xuK4/FSQVZViXVuz+qNIHYlxMTbYEIftqG/8tpUTZ4J4VI538z3IQY4w7S6m6YrOKpAcWzx8tJ6I
0D6eQLC6kKTqhSjGOQVYVEIOMV8c68e1JAroH/p4wtVbW0TLRoqj25BJP2BPYhHrwi9gKYxbQ1e7
58463r0N9mfL0Eyu7jn90ev+5Mz8iMU4gB0nHSGzeQKsIRAcIJBDIRt8QJJuWymGuDG7oA4FTSAA
c7mtbrmFAjZabhd4wFqbdL4LiRNvsxE63D471HQi4DZoBnOFN1KX1BOYjUxBV0J0j+jDmtClFGN/
jBmXizZkxaBdrYdT8ykDV8srdhdILvScs4a7utzTMdfW0SHIrDYEAiOPJuzB2pUrINsdcGKz4Cb6
GFLM3wdfZ8nFtoDMze2/EUxlS6QIjx9Sa4P8Zvm9S+G2GnpWcyfqQQhVZ7+uMfFneFIXFK8ytXmO
lb3sRQTugBCK3w9AtBmCnx7XizVM5t4F01mBKMWMGguP8VsfZl9wrryoePf3qLxUKwWeVE5lxeXq
f/vr64G+jl3eYgIWjPVvQ2yecSorluw3585C2HsOjOXw/v3UFsWBppCMSJ0DKhMIU4jJDuRkE+Fz
JXPGEPuk83pit36UuZtjOIH8G08FquyTeZncbmHUGhqgoDvlEwmDRSxa58b0jTX/KZYlKs0ZNKzy
SD9/XxksvUI7BwLWB6QSlBXNdnknPU5Fr+DvosMqxEVkmdTFCHujOb99/hpIdIyJzxlqWH45iypN
twEzxe7RR2GU4axva4wzLrPxy82BA/7JjteM/dN96/lTNfh3agfP9Pj/J/sJHT1qvJ/vI1UfiQin
rXTUHPIcWKPmfkvJIdAs7ovtsZNw0fitActwSWjxSWnylAPAc7hoeee/6TD+GgWyh8hge8ZbFx3b
KsfTh55sHESkzgMmQxQgdWdR7mQd0wb7ejID6p82GarPotgxGgyO4Fe/oNNYZYf4ZBxGGsTfJNdW
p3qu5RjC7a8sjK4b8ZHdNZGl5v8kS9nLuRW3IW730om47cj0Ch92hwAoQiDLATZO5HBDzJU5zNjD
02GXIICP6dyASdB0eGUHEVdLlN8HmvaUXFyeWhhw4oXd7J3hDa8c4+6VGxXrJ9aMKUYOYoBSZknA
gJkD+8XQVsGVEfkOtTiGyf2aCo6N1aTIwjXdYflqawzXYDpD1b93VjkErtGZBaHf1lMJZq4JBFbc
b9StiLtIshseqQL3i2Px+WH0juobKaWbNuVCSaV+muo9siwvHFTnHxxQ3PFR7F4frVp6LNLd7EsZ
P0uR3tb/ZYohWowj9rCvdTq2GAKTzQ58rHDhOWLcpMzPzQIIm5Ij4D8FMFnQZT8u/LD/qb+FDRBk
Z2U5Jmso3JuNT2h99o6qRrxhXyUSqIykfy7Dn5/LpnfgI9nKljJ2U19I3r6uT0kcjtrabeVhEY+5
o5MfK7iKSL2NRcMIzgX1PRIpIFwbCO+Ht/vCcqXQ7Gp9eKD8QQ4DN6DvyWOXHpSsqkzjnLjNW8SE
tkkGTfAcydBGiPB8Se9m8edCLW28QBAt6HuW/lCCWfE/gI8nqHFLbB7aHkjQQ5+drcwQC6WiJszU
5MVn7gzm5NHwHOLX6Z1rBzdQvffA8/5wOzq68BJatbevYSCigwr4vTAFBREzrFTEust0T+bEwbWz
WIeeZck86SCl7wv6R5eLL7olokpkGWIOGJbO51Uj68zrA/tumcgbI8ZyJGnVSFgXYRaPKSI6lvdX
5FIpjkENKZB0zc1ElDUuj5KSgufSAZ8Xl9p4L+d4rmx/5lYDArBBM9FrO4uD5qCkqiPVb+pgopUQ
Y7vnVy662kQMjA0uGiMKb90P4ACXwiCUZVDkfHxrKVqyn/W/Z5SFOgpFiZh+N5m45ghaTzstMRPk
xb2ukbWn3lgGU7gJXUpQ6MAxGHhhttoSLPEnONwV9GL+mASQzR6iY07UEEVtF85AbflLmGUf5M99
lDMluIsB3SCrA5H0jrNmXF9Jrq76g1CKwPI46z4we66p1eXYPVzOSyX96ULxzHeDhsvqMVusNWR6
Y0yD7t+xF4KrQtDnCMqII873teAaq6OCYOpLbyTI98qe10U8qLcJuGkYhyCLtLk84Ukltr/aM9yk
7tO7geBTW0yFRjj+2Oa0Iu+Ru6Ee8t/KSEoFDFHioWDdoeAk8GZNQ3HKCf2RBTxDviA7IoH2DYS3
KlOtt82kvD9r6XSFdw+VAx/g5HyT8Pdg8mkWL4cBnG8eAmkBD1oaQjebD4+Qh/avKGZMIgj9Vs9j
cnsW5st3keYTJS5UgQ1JAiCVafWIxmfpkt+Ov4jW1bgo6xT9shomiMB0+bmSr8EH8oG4G1qYdNfC
WysJ4upv4kEckA8XpEKM2cSheEOhhOxpFXQ4x3uVr3anpH3fq5J9PGEXUEiGAPRXzfQDJNguNI9B
lEBTazTBwdPKz3EudWL74xdMPi4PBAb1ZZ97uWSAZgrviIysw8sf61dmEeSWnqzidU1oj6sqDBE6
qxV7GkD7OTC5c1+w9dkj07g7OTBCps9x+t4xhkXM0G2im3PpAkHGto5oId+eV9+mcgxvMJSd7ad1
X7Fngc96EMx2Xu/yv4nPIavuaXpCEQrwNwna97xWaaf2Lg80s8ZIa9FPsBLdVrdhzZCcE30eLO4p
GAW5WmAYljaTVc6Or1Fv7893tm3VqJ44epKzPQhiBQ8tbQ2NuuIy6hl0ZcBjhvOaASzq5EZXNLvK
4y9BfI0MmW3WLV6QIn/gcAtaBT4Cd1tsPrGWupdJPTkVRju76kCGDWBd+RdtAcMxf8W17JarE079
WH0MIGY/NsfdY5/7zOsgm+YO7cWWAi3a1asDJHMw0WOqDrsD27JufQJf8iGM9QdZlLR2LT7WcjKz
0AL/+XbRibyVv2IB7DNj0hS8gL9HHpZAL9BI7RfPfZwJH3iwHK4dcA1kd/5Q7UjCNL0h4sWslesb
CcXiP8VzouG+7Pqst4K5Bk/4QaQ9KTrXWmGkyLLyO1CBHQmvo0DV/qgy2wahuxwfrJAAWAS68sCq
QuVfNcVLFmmpMo61AdqzpFOOAqYkoNQXpyfsh0iErBBh0Mw2CmUFF6WrST0hp0jExkC7G4Mh2kXD
G4/p3KBNJVlcgBL9LXly5P/ByYvxU1UGAcldrfDCtyHaTZkcEmUN8q/YID8gh1V2lYada2eS9QJM
j0XVLcb1Jw8Qlye7wDp2AkRQ0zhdYJ5mqeqBmdNl/dt90X/L4CFJSIiYZXnDKHCztl3zO1kTDZXf
A0XLbauQpvFVj+4c6U7Yo+0RW/TybbY1ZEiq4S4RFHoabFIpZhppwqih+/D0FD5EgYB7qhE6pRuO
hQhDDDnP32uUDGZh/SbT1/CbppKQEmVZuOFOnce/OdMiddWvmAmYRMSUduF6fetV7XgzQEjm8soe
Z+Y9RPn56sbfjvBIfByTs6Rg4GgnlAc9poeG61lQA2lJOX6tyIE0FZPAtQK/A5PWwSv0WdP9JZbM
vxbNaJjEm9C+oXwCAD8i8aWY7TVxzoVcY2CdQn5BcIl9KttieabKEQ0qHNalMU3lHJnQZ8UHjD25
3SZbVMbp3u7HIErqgvDDi15s49CXKvnKamwj7YJp6jTKn1ZoSSWfOdlM+PkweAHIS++bxjLOVbC9
12aL/ts/OV3uX5Z3bYK4mjceLfDjZWbVq81CPNYNz0j5t9+9RjbZjtisqJHtvVjaMnUJCYwGXVCM
+WILmHyBbYjh+TRQ/6PIAcb9+H/viBgsyywU8m0reoFqL7DLkXDRk3R/At7P8ZNKLVGQy0DLKGLU
KEmUhvThv2miwOt0okDj74oKIR5KokLfto1cLWRGmZUSJZ7BoPuGFpTPy4Hf7Bpzo5RqzrTlZCSR
HDPWOb670nax5fgSn8q0FQC/eKqgqjpYujnHzytKt9TDkXXTrBf44K5XEZnsrqEr/mG+YArunVe9
LNy3EuCAX32eAp9fUWaHRomvsB56AN15BgGwn1uWmtEDDfHoZOFTpgtVa6wljcwjeiV7YNjuPOEF
i+O9lhuS0F81Z+ck9OgOwsPSu5TWGswjoV+kZauGim76QMaXbGJF39/1GCIkStLtm8go7+GtD3dl
CgztgQ0OPyrGZ1tdqZ18STFaG99b39FDefKtj5PSmK+6Ny85RNw+8Jx/MjcWIdmjsZYrO86m5r+C
u28RfM5BqDquzOQSoPwH//DwOCTvcpwxWNoLSNSctEzGmpwNtnfBG5jgekiGL1I1cyzsRQpUlX88
iaH6aVNeTXiOK4V3CbBF0jz5gxU0nvbx8ySPdt/MAaIb3fD8aGVkBpaNSyQCjzvjoxTby+p9ASh2
ZbCZL9IXdjpcPEAC7cRclH87SnGZ6DH/2yuI4sswJTdoZuuYAu2hDWeV3TcypbzBXxeCmnYFw0Eu
IXvX7/noNcFNCU3Y7CDf0RKAorKbW1SXkpBXMuUhbajeTkPDd0fjyXzCHpj+OJlgDJiVGqWQ91YM
77sdajLoxBXZRflLij/4xau9XmgcewU1rn6YlpPpDltpGdS7R9LrKy+xdI0MB3cHxO7oVaBX6Qu0
VBBkXw+3tXYbr+7U1Nx6C+N3LYFwM60VTQFeIITplzQ4eySLVs6hhGC7xZjsm4Sjqm5H0P1X8lRu
LlaF9+5zkBUp5/tRkp57C+9sJlwVTQ3DiLb5O0ZIXOVx8yovdV4at6/TefoZpZWe51d9HocS+IEF
s+iMp1HIbroP841iBcXREM+hEmAJz6Yi92pEJ341af4r8RhEuc7DFbwwtADvTKjJC8n4bHZKuyqs
Ka7kXrQpupdO7fMvGLED2B/c7Zegw367Kfu8uWjZdugb3M4alAF0I+hRZZeRGASjsKtvFJeu/EFh
7TTbBiYdXK8Cok+2sSyP0PN46M3ubFJQgoHzfAQAhUAEjjq9NeOqo6qXiA9W+KzBCJIqp5drgiXp
vgangO8DlxtaicrY0A8GvpUb0BQ4i8S7js/BG9+Mf+uKrBTEU8kV6TA9MMwXgeRg3aiD+n+sWhgj
TbruCpK9H+8q51kNXbIKVwyNLQ1P7UMkR2avHApHtTGcuNt9R4k1nckI02NYe9wm1Kl9TH41f2nF
qS8qpyuHjWYJfdQvSarXDxUicDGLLl5GqH/bJYJIJrjBA078dJHVtU5wKPKZUMDC2e730j44BI/p
d8Ukn54SqWwb1DuHeMR7JQ2B2NOnx0YLM++qO4h45bMaD6Jh0IZjoPB1VaOkE2SWFo1k6yrqynb2
gto6bS4ffWacKsf1gKDrjSu3JNkrd/EQ36PdROZun2C7oIV3JpwW61SuAQ7abx0EPzJdoE3nBeEn
5VhxM3Oao9kT9ugWOjjKyNwllcJej3AqTvtQ4WzMMtJoR3ePl3a5kgkSc6sdykrydb3qm2fkgS0K
R4Yry1GWpQs6ZONT2ijXHDBi1ppd84TaTGtEjSFDBgWxUIXCiiwmPuxYif0azKVujGYUOz099OR7
kkXOSyU9HbjHDKpkIl9p17iR/nMe6P4QVz6ZotiLcLLJhMrfbXLB9F2hJIUIX7kdIG/5Z+fWTzqD
et4tZ7e2oxaoBfRRp9qGDDGkbMHs60Zeg9ERysgtH+JDA3DPsf1JE2HYLx0kmKfDriIdiJAYY9+v
OTYtUqQjFEd4eNl19CCqjLI4ggIeKcb47bL6EWA9gNKJPyzATCmtuLW7dfBG/wjSny9SYk86u0D+
MvwVCIg+ustI3MzQUxzoAwG+r/XiXYA7IwlA2RldkPO0ucpBlniYvjEd6588sakZaLhU/VGP2DJl
EH/cfE6L5VNswEaTA/0f1JeW4WLgyMYyY6YSl+NUHHf4JV8/ueVMCj7QRxt6GrpCmv48DhH/NKT0
/dvAqraiv+6nOTKEz96WvGSIzbdJ5Xp+3e3xsjj+g5Sz0XmeW3DkLo3zul0j6rf9lJ4wcLIlegfF
fO4hSTVNLUAT4X07+WsTHS6kgDY0OYmcEB/XLmj9D6lWODwUp2PcV6W1Vo5NwvkDQykOYrc1Fm7T
cfU/0ccjwqFhs00xO7vnZnjZ6QP8dynSBJpIbWxIrFFjsf/ckuam3bP4alJXNDMYdEH0MLO4JOlE
txklRUnZz2alIQPt1NXt3pKUzyToeWp9fwijVhp0RVYBCmqsj9tOI/QoSb7Sns8fwrtshRZhmZTd
Jjl9cZudQtMfGI0w1nqlo/Gwm/LZbRZq94uukquKqux2SU4w+CBwOYPhwB1SEJlY3fPP8jGvaK5V
Ivp7tr2Tg3+Wr+sX+JJICKETwuLmE+1fPtcbIlceUP02/iNZbnfyBwDgSmO96DgrFdNRnpJTKAOU
9wMhfhQ/RYK0DHTG6OdCnSBS5bYEs1r6mpbA6Xfs8IYLdEQDY4c76cFTd7ZnZydhArINXZMg8zkk
51Ey2FF4hKfYRf+5B7MnP4kdUopp9KEetowTxxWqeb7GNwMfuw86UXly74gZFDIvfL9UibXxdcVj
lX3vUKzbdeQHGO6Nw0YmQuUXG6rJ9XtUrhBRfkF9RHT2bYTUg/tom6LQtbmN349IqOsaQ2y/8Y5L
6SgWpvzqgs29l1EixpWx8H2bML7vd2CChTtEVxj7+ZsT32DHSsO+CieOr8jkPVvZ6bduAwC5K/Nc
bp1MXI+Ai0W+wg9XMoIEDztc2PHY7fpLD6uulI4RDpW2cu98v+wKKR4VkhmC0pv5d7nS58c/D/aE
KAcnOWNeROGsUxSQg3VhU0cCBZhlDfrc3FHzw6PezyWNPBLLKBwgHC7FJ5LwroU5stS1NnzCo623
WsJCtCbYHKoKdmDiQwUYkC9RvbitX8O2n45BzWGWhf8/9LXjuu6Qcgra/0lYS5intBbGq+AV01fb
NtY/Ghs1rKiPXluyTy31986FoQcD8p9qlQf5F4QBSkRvKl5scoKdWn5TGUIYJaJxUD7LGWoHDLSl
lloWUP6GcxuvwEPLON3EtslvoxCB03hO/XzGSFTbH9hYKcbGbDEfVqdMAn0XWl6mcujs9wIxcoMU
3EIpALoIX9Z0EDPm2qLJjDEhGh4Ec6qOlX6z+qpBoQMZoX5bG6lYY5GWTHCi/NdKstRnwEGBr/W5
LdzDK7WD/sA7IGI+8Vc2IpoDibvLXYAnpHdz3WBmsv2ZS0w0BHE4tB3ruG1EF0XgimlktxXB6kNe
t6CKxgn12XN47M3csUr0LyyYMyrc2ckimd0632WzZ6DR41g8r/4HWmfCdzmddwPMqSgWt7dCjGIJ
ceUsmkCGzZmWKJDMUAuvVLA7ycxLG7pFV3w7WPrYwmWqvex5QUh4QY5AufxMZtmqpB0frUIKKJoz
pe/2cfkpMQth4rl7UI9o9v3gXKDypHRbPz5z7ekqfopgNClzBoKSYgP5eJJRqFSWn4BnMdEyH8pY
RH8fd44EHA84c0syJLbJWIcf0Viuw9wt7Wmd3RtetEQgmAWLI6exyz7EEO8tIsS9qhymbLSYVAXR
iQ+BHB/qUXc5QB0zylNYgRRfukihUsBGAu8bWeVlF6IoESqznZXNGo3c8LIcEmEoWg4YVuiBA6Fi
qjGSqIq8N+0R2ctEvAjOJevOyNsTHUg+RNiG/7sBB5l4eOUShUdeOUV7jFWWwCh+oeIGFGtDotEZ
77FjqUck7l+9oFxCDbx8th/5KxMjWbNR+cKYwf8iFDN9f2WUsQXyzLaaWxo8ZkfTpmunSkZMlcZQ
K43TaOmSiM/TRwl09VlNxX0c0d3FrZBOioEDWYC9Cfaqg4VrreutAkyc2ozibIepWt2a/oXFdGiI
ramUZJBM6OKqi7Plmq3Zk47P720Az7zdvObtuTH0E/CRPFsUcrqnH0O5Swsstnse3OuhqNDfw7Hu
A8rJoawwFxifpuaTQ7DcEPt6A+KfTSzbRlVKarng9iIjhgo8qr0WILm6lsFtGGBzKHZ5ne1Sg8/8
PooBCkQxDNgsw9YvLwG/JVdk/QaD29iIay8pIBfFdGETjo3xu1oK/8pJMxcRzhpzt1rHKnzqWkbe
ZbFbxUaPbX7MN8bdmqz3HSos7oYkgtnOIL6w4BgMBGHkbAERXykPH2/+qhJ2XDV1bJIKU/huxKYt
0Nom10LWROOo7EPwi5cLUoaMN5wzcxIMZT1NwFFUB6EftPM53HK/I8bCSPsRb+up9FMv4FriNe6d
htdUcr/hqPHyTKVdAO2yUrm+tm8xpS/0kyUk3gLX2TCw3Dfui7kmXpu3UIiONuIeo+Pg0pQdBOu/
RSNlYT9FPDGrbj6W2iTNcQNQrUzkCUOdL3ORdGwclBmw43qFpHOi8Vm+ytULA+wViy2dDiot8hLY
3Faxy5lBze455VMrUikfMbnPRy9y+/ykhh5W2i8Pr4iqltF44ao4ZakRyyDEPQ5g5WNvO7ce9KkM
gL/wulvqjakd+gdpIcrA5yL9gQi50Iib0Mx4wGoKQ4J1o2MJjSbRC9ttubqZVw4popQusV0Q4VY5
9QkWXLJOLTqJYE2Xy4ZKuVk1M7g9E8eUd9A6vXg71nDcF1qR0JAlPm3J0hhQHtPI/WHWRKEmS79z
vhYPROvwh5hSBrRXXg77gEdy544X/Cq95fNOgqngrYhHvleJhz1R7Mufekmr2fUzragx4p9q3894
DAU5xjAPZp0/vDNLXI27pt/DPKPgyPgTySpoFHlCBjOUc45cbyxJ0CMu6UFywMp4xXjNW3v1KyGD
g8yOTKxQNxi0RNr6XsEW7vPk8U4vkA+FT39IWshDahOfEXqp2rrk87T8Ifs7FPMT0DMwG85xtlKJ
xMOuV+xuYXKQqQUzfGdrVHcf8XMrXWPHmr69dZzgCA3owX6G+REH7DsBGYeqAA5pAMYqFaQD+lmS
CyRGJLJqn/7NNuoQBiySP1Uwwp/fGj0EpgP2wV3GovGRJaNS+oASEhCJBQYsSdfqyykETCkSYLNA
HJIU/YAtIFc5gTOiI3RPbKP5uzePeQ/XKRhEeX5oDvTE3o7D0kA+DkHQFvH8m0lGJmIoOorFyGB7
XXwheBG9a4F2CLxGx1Ar3jbLrOyaPE2x7eJMYJ7u8hfKYyHzyPswh0kQVoozp0xvN8GaQg2IPOiS
HWHVHNa4RjLxzE0tBsEXrfXNHBZjjJr5kFUZ3SIyH1ogZhc4SDtGo58oXCjzQ0LrHICFF/tEEvWW
kbN5faDINw87IYHEbAbKAcEgrNcaRovVHuoInpq9Iuv4/7vTqZggPHhG+JyFAyzvzFcDA0QOGneS
fTUfN+nB/Vyq+ooYml4M/BhiDn3sTel2TbqhqqTewqR0gfdxlzJaAovQULE1FA/QQZPGy7zHK5YE
9Y0wOzVb0YvjM0kaTP9j8LMbTY0Se74mZ2bzIMYEJjMhouNVGpBMjPOyt3M+LD0Wcvn2G2zqsX70
6IICFbliCbL8Ixev/EPR4cJIqSB8VTeL5j/ftp+tLosHncA2xbLqKsbE+UzwVBLZ8kPUdifUOJ1X
eTG2tJgx+tbVQBDIx9WmyliaKE9xUMwC8DDIiAxjoK20TrHQQqPVZA8/4qLCGwOAmloKtJX1/pgG
9oVJN13quI1BgccgKAkufBcPp4DwU3zqPJGwp58YemPRN5gI7mCwmtjHQHXlDS0MCU3v8vrfshJj
XkYmGnyoqN6wrFUxmxd/0fFXQ8WUHs5JkSUk6CLQ6aa6roV815u6ppXF+i/nd+qqkDddBBVstUCf
R3QM54JlokL9wmApzaYnDkVoCU6LulCFf/nXSmNW07hwlQGxG0YwxE6I/8ykLsJw5N80XWhlPmLW
iebX3SzmmR85t0HN5A/jyL/DmvL3K3ENu0e8BbvzHzZGR+yNDPPELw7s6IzL46y+kNwEfaYB0ke+
h6aJ4wJDirTnTGUF/T8j/wwgGUxsC/aenRw/dI2fLjs6Xqgf5uu8Y/ERDGHE7ulwoQm68AEAk46+
dGhVtt4T0T9wl7mA10VZEvVom2a5XdvU2Jzl+B+f+cB4Smli97W/PEvNkf62DUnM077mSvnCXlK5
wfnCvmkEchVRTUoXUHv4SCKYGRs/qe7tzGUD1EfigyCldg6xGnJz5G4uEFHiNtuc8rUNqb8Ihd4T
bYV2BXnR9Zu5XAMpedeJgTz2apUvVMvkMQ1eshA4tSX9opGA2cFSPRFaQQ46uVm8KL+1KWl/L2+I
X2zZXPvxkd2wfe72rEo8vSRoSahIlvOCvVAGa8SDR9Iejhnw7LR8JBRqLcIRxKa66nxXirtN/xK/
a0gtT3qFPylIDUhJdF31SMf4XFfTrS/wCNEnzK8Tfa26DpPSy1fSo7MFk/D4FqiGRXUm8gdDH8hb
1BDnHiHM3t6fjjjaa+ys626r4rzwJK0qRjQpa7KRLZBCdzEtXy3pHB+LfDyujrChuh9/qHTPm27T
ofMsOAJEup/UdMcdbSasKdxJWmWFR+yAuJwDmxilLRrQdhkRp1iJcw1Khe/eF2nd6mW64Tx1otBr
S0sJx11/IHpDmOCsEXffzcrjxqtNMDY1jbgEJHPFspgkKBCPxnL7ECE020OJqBRVgBNTf6a63u9/
t5x8isyhWAGX6X2gjbb+zyEYQOYBxMlLRFHuqLsbjKNu8ORnhdlzS9pFCW/pVrsbkVzdYnClbBsb
yZzw4z8gvaCzcoArPQlEp0WThHagWtKtIh3rT5e16eDJyw/J8Xs1Xmv++UsDypV6V0HC0rwpUk1Z
aVpRf7sPBRaNM5eG4ofT5yG6RfHGmZ/Q+26sZl3M5vkB3jpW4mstq01K0LMxCtYBN+ADyx5iRqDx
npX9uGlvOrFC+nMdM/c3t5gr/gtbBJd/GN3Jl4tpH4ngBbh1GjMLecT+zxgN0upiD9WasJwAHWw/
1K1d/P//F/kLqhL7CMoLJU8kbnlsQFAaMUjfJ8D5f1nKE5Al/0I6NpcxXXizf23gfAFJqcgaBTK1
/uOJlDDVT31GLrdtdF+BysKHTmq7udqYIShyx5pXpW+OCHXaaHf/4urTLh2T8+reus/wK7JMBEnh
zY26M26clkZR0TQc+Ci2c55B8aj9shrdEfH6gBp6vTPajis2H9SE6XWqm8iBibjAmEfSgKv/WaUV
LY/qgwJ5GsysN16IDpYGTbdDcnqDqlaiBj130BGUnq+zc79ptoW8doGWMwbvL4ordtRCAbAxDVcr
ngAazF2kQBy/XPtiWFaa7BK2AdBqptw/C7gUyELWV6yUDWFdc3xFj9LiubHNrqiyAIo5u1o6VDHB
7umCS9E0JViz07SnT5uYuvMYBrdl/vCnXVuXtHRRP0o0RGpdoVYW5YqsYOTvX1eklEaJVOEl/8QU
QeRviQSjyTgwujKEqKtbirMeJ9UqJxwhzJedHxOReXezbVcuf7RpzAKGbVusOSxIVEzWIEtch6ZQ
biOaug9qaDRGLnOpC5z4j5l7sSufKXQ81gzSpf67XDWdbyfzbGbOtZdEsO12BxdAfzV1prdnjNcr
nxMWw06VTEbIGQlYfdjpM2D+vJklzSJaoVigUsiV7nRl8MRf/PpjRRLlq/n6VbK8y/VEpKW8mtYv
IheJXeg69chCvblT2QnboESZlkMDx4na7KjSR7ZmBDi32ghGIGb2Ku0LlQKFfrkShGJgZVxzSE/B
ZIGgzEL0lyPZp0ys1IxaoRI/ugQ3wEa7m9o9gZMQWrPeAkq9BeeCWV4eqj76Y67P8Npm5Oa9Whcn
W4k4ElX3+r+eBWCC/3JODu8kEOVmvfsPaEWUv20MlTIMMjEaLJKGMQ97ouB/ouPAfW9pJTJiCRTW
mfcAXugV2RYy5iyuhWKpuVeE8WZ30GokJlDxBp/kaZVmkoxc4cvsjMcyNKdejjxxnDdF7X0Sx7d4
ny9I3qIp20BE7agpOVKRUs0Rhp0wHIMXErYkV1IjbvPt4vWnNc4FvU4AreWGWNCSpjrMFwVR1LL1
QTl7Q6QWinc64+0dXxzdqKvX+CWOJUkXJ1riFrwRc8wLMU7U4z+bBEkOhrMG6Lh1bJmyjZoj+F0g
LdhYuxausN/d9KKm9kSlgnwNSwkM9QXqxUy5DikDfX4B9hOt8hN825nXsCUc0I++VeX+rQvJDqzY
iRDxDGvC+nlU05zlNm4s62mIqtalrR5ZJ+rumcRLIr7LqxdeZbR+T5lNSQNNzemccKMH8MAeTVzP
neTNWX/CxUQfrOzYtTpIit4Ik2BEJUW/rmhS8DiRYXW+qj6u85rsOtXp4YTEfgEBf/4K2lXDBS3U
8PBpE58wm5a+otvxDn4pteTRMaRzrgTkGPmlBwNtOG1BzA2/6/0bKjtuJ5Oh+EjMr1eTG7U48rA7
OUqif140Vel4x+FBT2I8mGnnODNCtqMSB+ya7HcIdwFYMk1XvAzyPcblsqiZ69mkh2Sq1gzB0xzm
nj8QSLZ5ILFp4TnEV2R1vmUiTXBteU7419zMVvcgcyU/bpAaByryT63RpW9U1Qzp9hRcPkbMhmIA
gtjGqT+sToc/ul71dfIjbk80qUCXQLKg7BmUdvJpqaR/AzrY+vhZo64cZNWQqVAmchHMooRzTxKx
tmet6Gs+zD8eM2mI51BYl/fbe8hqpLkn0ArxHFs1r/hGFgGxIObrjHNksSYxsLih2FCHn9jTwSsb
BYe/7zdKaVBRJvYYiOMtfyVwhXOlyavSsgrR1HVDYlDrmVPBBDwg02F5NEs5mUm5mKgKBwxRt8JF
nUJveGcZeICgZHm3HpaZrC9m5uRbFh9sNZ1O+tWJ4xIW0/9zTx2rqJ+hZLwxozI/BrhHe8px2KNx
sT/Fb+Im6H+QQ0dmtckPxobBIctp0d4vzj1XzdThF51fD1hweofONLtz/tfBoAHgJsTkZGP5udUk
wk+zOTrIJx/w/MVWS6pejEYXTbLo718JUanfuNfF7Njqyu7atAjbPpQR1WKH67FvyCYOAIYXKylZ
BHRGnTRoX/i1cTHLTUDLNCvIRQBXrNPsmCOgGWoWod2S1ee8usTCYforZej5An+WgzxXSZYi+XiX
WfnpoNYOKtoNxae7UXwdHTqN0JWDcULIml0UrQof8SApNcgIsQjD0DjViUwSKpr0OtA3gioKAro6
9DtKZtCdR0cWVn7PmaKJSY98OxMJYVfrJAFN4n3DttJHzMemD+2odYSxYAdvO7bXGgHPA+XL41lt
tZ9lp0NeJI6uM34Upu4BjkMK9SPvzDEeHaiBIjRBz3E6/lhtMUEBTk+R6xbLnrl2A0dULkguUSa2
z45AsNICtrynEcdZGXWg3G8cDjZhGA04wZDRXL/i9nNtRfPu67AWAnw1Ns3QT74nTlrvb/nI7imX
GAbsoSaADeWbBvguzSk+fEKiAZKpmgZIMlc1vGtqwLpxk8Ys2m27rL+7/p1ihS5TLgzzOX8jsXUM
FREKJTZbZtnvujmj01Xy0u/FmvR5b5UIT1bHu2RKDYvV6I3BG44kjccTX17UL5R7uwEp5mWLg7lQ
ouKxeOs+5SqHbHLEd97pFluzcMZZwjY2pO+Af+C7aQcZs9erNU/VRN/fmAYZ7r73BPjJk3RMKmWn
ToW0tKaKyJ3ml+0zJzd2uPLjB3+PXp/C5BPDcwgCfZdwB8o+KpDLciW1yaHQWgdsVWt2h3na1jea
OCOS3MUUm6h60fGLQbXtJSB/vTY9iu6kuTmYeHrdhdiY7eC6kyvgKFpKNOTlW7Uzs05JUBfsCLaz
d6YmkClDD/zPMVZLzCjLCd4LG/SdHoSkNBrY+CJ993M/K0QMve/3CBqudQc9QuzPfj5myy7sbOgk
q+cH0OX39Au8TPyaJJbUaA3l5yu1qk4Y8K9YiHhqXXoUQRknqRvd3J0KZBVL/yrHT80jCFuV5V58
zHecRZaGLXzjozRy0Bz9De36diEep0pKFW1jMxthL02VggUkZXmHINsRVAG3z6c67hLuovaizERt
LMGSNaMShJsfsjTBuzYUuM0qKnXka7bFlo701HyOtZSLD2G8+vnsrbtJpjg+zDG6l6xfMWIe8tbm
BpS2uLANjehMcizJ1+UzObvEaEQK/EVkg1CC68Pq+Ctj9HvvWOdA30eIUI5ACCuhZ+1LSi7V0eHG
Sa6pk5XL8TY0mB3kvaZ1Hb0SyjfxothAjhh5AUMmelRHQpejKds5dr2csWz065EClVpqGKW68fPG
X5Y/dJV335Y3I+9V5EOxGjAJ1Qo/CsD/CIEfFpOLJtXCCaa8O54KjlGOX+7LAgggQcJPcMmmQ4E7
4TnyM/TwNU/EpfW2G1qYZbetkziZUAmQH2hTfDdEgWMRF3pnHjOnyYzFU9ueVHdYxquTQpfbb/Cg
FZwyyW2G/Cpyy7ApLH7TzWzkMdaT08PQtYQ27EJjpJzzSOAVzj2gRQ5qjZORY4RdjV6lxYgtSqom
UnrjtqC2HE8AO55wkzjXjKAsvhMwbXxa2bmE9V5XoAbC+E2YQaP0D1YKuKagdPC5HD4PJi9YfPH6
BACDcHyzPmfO/k5hpU+VtZiEEu18q/ZI6c/a9E0CEGtHZwU3dkYOthln13KskCFJBP2D+7Q70XHi
gQn1CTedvAg9LLNpP1OL9LIgZKOcqpaLoqGS3un0hPb4BqU799S5myqCt/0JmK3RIgNZfM59P3Gf
ZHOG0wmwvrZN0nnam88v3Jqt5LYHNytxNP1BhkJrOxup2YNEWiUPSbqq84kEVGj/LPGeg5zsfy6c
XT7vsJAc32+w0E55woYBGxXMEHsAh8QUVPtzfmDzh2EVJtBEs1NyENigo4lvCUWfajK0eHbq1XKC
8qZXHLtylE+LPrdJvmj6m4zAQvLw6UvuJ5OpxOw9z7VQAh76xNwu5wOpb6mGcqwZt+5trZXEdGR9
xoxVJut+nQizgdqYIcMxZvqFpSJHV5mdIRLOHypwxvVtIsGP/Ivh3qLQVPxgl8yhNg7eoLfNfxvh
KV7MJ0ej7QkZr0L9FdasE8arqNbwjnBXbR1vQvZZMLUFSp9N7XAgFBymtlUelIPw1qprCTcME2cY
bMqnCBT+mHvv6Za8M9Gk6CGFqLfn5Y4U32FW2ZCWgBis1TV5WDhdM2taMGc2lidS+B9uQH1Iy1Pa
kEKrXt3JW3wdAlfBAwcSR0R4MttnnAHQvAgUqdDWxW49Q0SakLL0GdEgzNB2rWRNd0AujjvoHCJ2
cbOPTGlFbnUTurpvjQJRuS58gkXG0QWghr8IpNPSxLoW4omMo+1/Ik+MH45holtvOS7n5gAjlWnF
afvn4bAvnXUXTCwFMrNhFg1TMeJIPk/TA2vutdBXxukYONmIR5n6ujBIErV8Xo0oImpF4Q71z2uB
+SFxpLnMZS84ncIc6oWt9SP/rUrnf1b7sikYdJBkX3PeI6LMiHndMIhiQgWMRUuUBWKmxftESYK6
p729qCmDeju7dUg31H7dqfAflNSykGWCEFEEwvqjkKzHe3GIkrACM78FkbkcCXRL/0U9iBxPRFIF
XvT6+DVMHjLmF7eizpuPSdG1HYH/PtxXAmLWP/GeIh6OpuoD49AoyxIVkAD34XayYidoafE27XHn
OJrfWIEdpgR0OSL62B6NpInfQJp7dpx+PI5zQ7YQUi8ufjzYGg3EAkrGYNSKqqc0cZFfiV1DFSx6
Dg7i/602bJ2oG9oNLb9eCHZRhXzDkKFJbBgv+PyyAvW78pXryhhdxdLCp8d/kCg4DpQVNtuPTJSz
FZLkYuHOe3tJqfNQgnC+mjyzttC0V7H2zmeNN5gpjFZc1MqicX4tlP9KawMEilJuQHPSiA3NJvgw
8F79DOO96yDZW6YuDfekbiu4m2mkluJ9dq+Bl1GJFR4zoeYpijQu4iuOltHphQAgaB0JcObwlDw5
zSaXLDmvxRKcQbhN5QL1IeKTmFe4ZGKo/mJ4Oh2dsJnv6DVhIgskNqsE+fwutSd0Sq4aD1RhkIg+
+mbznkez9M9rZvtjeYfN9cxAHjX0tCeNyRAU3wzRyaPGyasf3pfZVg1BOuDn1RxT/rv6k9hVkdY0
dtsAxW8AszH0ov6PBLLN+HASovn60qo1cxFW7RPWypIruogTdI/DNVrTg1oFhQeC+CFaMDGrhsPV
+0GwceYvaH1UHX2TJSn9KjVbTTmxFztxy78Wz/WRfVwNIPqT1W+8+7WxJ8a/XQ7hDGwy9vWdxtbY
rwgZigOpXFecnTuRhtJ0rrQ93HmEE3IZJ6G1WW/3n0lpOQru4xXap8AX0GEu2C7mF1ItO5r+d5p0
N2wbcpwVbh4dZlxHafBovpEXEFpLBVXeIeCNH7AL8yNrcCdfDGlNuGapk7557i8rlkG68a/KIKDh
oA356JTAhA0sm9SY4vVMDJ1H/pUqCXl2eTGBb8La41h6S/LQvsGPKvXOKyTIGpApMxb1Ae4aDS4O
gsu8rPZZX9QLLD63gJbyn0j2I7Jo4McCuH13Jj03EUHHuunm+qcptG6VVbWak7QGnbuQXPOfVAB9
T18Dy0N3AtIN2JZ9nuL5s9JGoO11NnLnqrCtzkQAjMqNbuvWLkRSoc638vaFPMR0TeoMRp0s+JnW
LrUs3423dRm/P0OT6hBJIHc7um1yYsptxYrJx3JJKFYPDFrgRxZodvaJZ2ZZb+VUwusi1sKxX9/c
unc96B7t93QFwIjynCjT+BlRTL7lHLyc7vyK/fpvlVxbophQWCUG9xrJqcSSrohuTfsLnNJ2o3cU
A+HNpjSFLOOahjBFd8ghFE9Z4YKDSk1a/jwHwJyXEES7LkHtZ+zcZOU89J7kaKXLNxl2IkMWsTZk
+qMyVLeTtPl8GHdKvKIP4gNOVCGJDSw1zOVOWhkc1Q41EOvBP4AqeUkrMwrHfLQKL8lDn53eqyQP
H60WOL12Xcj0qYOIN2n0oz+0fSzJIGP6AMgOlo9ddue5mTAcKQPFqWnytrFBpLO7SPKO8sPFSDIl
4M8JCRJsJT75yBH9L76EvzOWiITIjKp/tJ1xccw406IhOIZLWHncxbIxR0BLjN5f7re3tHi6g+eU
J4q2qbSWiMWgJZvr+sjEtYCz3JFQX7uHlFBcu5S2mMzjuu5dcLz/PWew4/d7eaZCrxAukPVQQsZC
KHmMkj5fH8lCpz/fE/iA0giwWiIg9MYt1qS/uA4zMraYy/UWYOoSgQnvLK5zueyGEmkCkzWk6ZZo
YVEQuZ+fBI5LOeRYzvVaxrF0HqM40qF5O00UD05bwUzxVhEwz9MtYlT5Aihm1OzGugcfL1ZO/aHT
qzgVnaRrmdmIjJdMnkMPloeVakGChNruel7UBzKuAgvVqTDwpuxlqxQvWdzexsD9ojz1HccRjpVl
+PkvNOspVQYBGnUG2ixFerZPX8Mo5Q+pRZDYntyB0MA3Qx5971Nfze8tetq7ikjgo5mwfu/Z8BgA
Qruv/XSzDwXgtFstM7JEj0Fe0npL9ZHWewxUiVA421VK0wOTXXVWVdpNGtSgpMqze7Iakt57c/1a
TCxzri7WRqrdbbCzqT9qd0ess+4rlYn2Bg87qpV5MchuAKb0HUi3ut6rAHJFdQuxachcJY1CxZBW
qVnJ0Eb6O6ardI7+BGXx+M7DiayLpFeDq/NPnDXFd85Rw4lMoAdEQeX6Y7LLPeYjvtB7UCQ3eDVo
E/opjTOqGqPTJnLrfnqZPgya/AwpoqIP0BlxHjWttvbfY7qIgHXuZYqYUmbAMdwzwJiWib5RMfIU
zjrgt89Mmi+h++S24ihaZbLhv6fFwNrXhfmu3exkquG3Dc9AiX2EcppMK8QZ9bKIBprLWWyotOqK
5OwBtb3njCl/bDv5aNAOOXT/koJTr3uM3598RkIupLGCp5ffbTUgVQg49iKGeDOe5WbLgwv3TQzO
/Y+HDpciBYXu1LtAR/FJ40zXMR/WZi84FJdT4G65s1UPb2+YubyV/OYwLKAbwbiMait/4839DhkZ
9TCDW0ybCkLwJGy3EAOy2lPXId5ms3K2dElthaDX1/qS3Jq30YGyxbodWvuxxu/vxexbZXUpLJGS
K01FpggpgzSxYmCo+VmVj4Rgx5qV9/w3TWEwlPEA4dUTZlIimPIKw6Z2UnDj6OL1qTatlmZ5MU4u
CTXoOBW5plYECXVBtmJl5XZLfyjQadIIIYcqAkhxcZ7ivPYYMBOg432xlVD5rggU23QlR5gqcpYC
4mQZwnROIRyFY/KilmSljKGnxkwYeYJNVv64a9mFjmjfwsKwzabZCivB9w+CVYOceyin4mDW3+yX
hUsEcoj7Fuc/DADotG3dAYvrKxD4dVy5TWHP42lT+x9TNv6vQsLAVnYZevBd76z0P7is3t8bp09j
S02V4sHxAiuOU8c8knmFDi1P6PgIZF8BYTdiqoSwfA14EmgmLkoI5wj6oO8ZKoelQNZAmxC+enqV
ciw5Zxj7AxO9a9Rr+dRT123wpu/C0RM4JGIz3fSJAHMWnjqeYLq/Z4JbmhqMDNv5pqKszNEF405a
fC2uWa7h7Dpy8ATlNb3RB+IWyv/kKmFSs6GqLvEeS2gW8t/IB0pdNtij/OlJ4keT2LkV/+kgraky
B/B43NIH088aU4904oJIO8Fj3GHk151eIWnzq+jNbEkJK+bIFOHCqNSdOmORrp//zNnTHggKSqI8
HUcBXISMQP5BHEKAHNvpqbhOKBpvxkQV0chBwW+IczIXo42fzL+HyGcYGIO/dMLFo+2NKoHYlOIS
WonDmOWfUlIuBkXjW+20b0GEC9nI2ozKkrVppxBoTyMWt6VJj5o12oKfrCeAEvZlkf/RZtVYexqh
UVY/yNCkIoUpsf30z3BrasgAThz5kPpwi0kiF0NKXM4PYSW4W3h5YY0U9SBcZd0xFNuh9x/35tkc
yEbR45IcfS9CvgeQFU2cM3Iu47hJgsk7IgFQWHDBsIS0SJ3t1+tjO5qpYmJc5kAu8SvQ5AJjMchd
KXG3i91CWTfd1v/NVGW2C9lLo3CPyh7dcJfB3ocsVNQ3Io0GJdZ724zVFyM8a0nWuIoz3kftPvvf
S0P2POSeD0zS/z/o2jjD9iyIXTygfbjiQu8v0+uQCyheTm/JGX8YMqOi6HodStGapxl94sb8fFJR
FKud1cCEGOnBgVh7owWVrrUsiT+AjGOfXkNsZ/6+FJEE6TekIqRDzrx2j9uLeEMX6cbbz0ZA4b2z
XZqfbvwdzrwebLHMcP26AgIUOOG/NkYczrtkqN72dvTFnYSOTDRVSYfqDt4eGbo4cp+zTaAM4aZV
88VBaVm1A5RML/cq5AB+0nMkeKieR4StJkgvRzLF8A/h8w5vzBh5OunYXaMbb9BjHnS+ajGh6LwB
IBKQN7HJDAhd3/N6SMN8ycKQdK++mpw1jWFXU0BEo4ovDR2hgYwOaLgkaSnAtxsZlOdXCxOUdXAy
iPt0SXUUrTdu5nU/R3uAeVaUSV08mLI+EqG6Bec2A55FzjcFV4/uBAxjO14XfVaL8MBW0/URGTKu
qLjzZWsAY8WUQ8RFLsN9cc7VcTDY+Ie5ulkKFmEPTBI9M7eOLQeaZhy1nHhkiaOMZ5+IXZxKsNxN
Qdbo/Lb6j12Pcjnj42ZNy35hLdlRw+2q+l0prz8Wzrcj/6CHXexKDN5ynt6Ux5yK3ZcsmwgdIYY7
1NFzJGbP3oOw15msgZg1nir4q77BiCicg6pHW9HmoXd4VsKF8hAlyz/2+uzlazdlWeS6yYjKfDAa
tsxWKq9RK7DUM9TOXWpqUdg1H7gl06UyHD2gZKRebJ1Qvpgw/0LEdr5Q+SUmWzQL5YomAE8eJFZk
u/7dYUExSsNLuiHF7iMY0SLPa68EqcL+/UwqRBn5cNbBlXleq6ZxTHYzhQjHPW50q0bMK1NtTYQO
2qbs6wQfNneufWLS8YWBJqGLS6qKOCmbkbFH9bL4TYt7JF607ngf1l0OuHhtupxnPqs+rOB5FG/D
TrG92oy9LPIOGPRt1QEu62ioajm6sPBMwCV8CiUIuFiJnlgmNH2KvHY63mXBWa76YCw+3BECoj/W
NuoSqdxEo/C2PODODunROgnmz91yO/8OTYFFHQwVwHQKiVYaHMzYsmI5T9cpbsY3Xg8+gRTIg//3
dcW/fx/Fk3Mo9N65v/fOm3v8AGRjWwBYLLJMhvI6vbUQTh17skRtvYix+BgME34smOfriewXdk4m
+6DBGMPJniumir474qKPPbgaFTpCINqY7OAhx/g0m9jJoEsKOqgfZFxWNbE97h7bAYRXgNTrK+9b
+vsecvaz8ZwwbyKW6MSPMaOx9p3UaV3wtKuufyyTQfnfbk9EAbc7j2o3VAug+13DKc9hEdNc7sfm
C5WTdFWbxw/x3GtsAz+cmNbFGy9G2PAed8LMDv6MT21+u//ZyBN73PlQ9VxfZ3I+c0GtHxNqgB5u
Blde/TA2c7itkL/7lISYIGT1URYJ0dVtus0Ka9eXz26EQxYotdWGfvmQWAHO0Nk3f7d5aad1jGfS
7KVZc0GqYv2r656i/oCJIBJ/3XCZkJotxojH/Muoh6AHaaKonM9KTU1vrT96syBBDczbn+lP9vel
sdn9LRAD+Ql8huHfP1gMMmfvc/EXMO5tY6CQQTkYfqnSd5Gky5XLAW1xeAai67fdHZ9sG2fy79vC
ZsbhmqUKHgsoewz52j0xBeX22RZGDIUHgULKeXZdOd/Cda2Z6L7C+4YSCHmshJjGJ+TtXlE8suDg
X0xbnSMB74+1ii8X/pu/NI9A+FKRUStgCD+w7/XRHxvE6HhM7LzMAeDWvzxm2mIMcqfekS6n33Rh
MByrWebILR0PkVU+3RsCMP01ynseMEagSEA2DZoxqTu25M35LIPWJ8J0/SDjLa3Odb4WPv1k3A+A
YB1wEn19g/w+vo50L8No4LmMEZ05xBYGc4+JaPW8R42bigeAwxyKRXgd0K4coCBRUmiemJNHKAPu
OxyM/TIILvhZF92bn4CX5qTQ3Hz72uBEr1IpoCjEnkHlQiwQgMzVHgNj7WDfk5NUYHuH858SldJI
z45V4KY0fYqhyIW0eHXOgUy1cdHnLm8jJ696C98IUAUxSI64PuLfIfksYUHLciu2aLphbh3Cgosi
wpG4nOcpz7pImBW1qdtdxvRID5GMnWuNkBzUmkTC4WY0pPdscFA+rtASHc5lTYPyB7jm3riVxFmL
RHsnt5yIM+lV7xEJj3/8w9MTog+tzL1Cgzt7/GuRgUci/IbDkyD2OPCNc7Ug4NJZtgPktoXt7fnt
l7UvRGG+MpKB3N3m+bsIuKVHbfzSfWiRRqtWs7IyA02BObD/6NjZb2yhCWhWXs06rCuzBYK38vxL
5tkkr8W4S7PY4hXlkQ8tbUyeMRFgVWIbGYNejOflmmwNgATQ52F1NP+I5jUCRjVehr5jwuYH4YZx
27oQbiFaFY24LBeVYuQ5ZJIEeBm/QgaRE2VYP17S1+Ytf9YDNPCL2ZG5/i3QruCWOTUhxKc4Xu//
vs3ZSbF1fp3MYbpl9ZU0arz9yVhL2iXU1dKD8WXxSXZ/AehMWQhI4R33AifGNDzREhcK0TPTXRCo
Ju6Z7ri7ahEf1Nrs00aPQUfXTjblSjvBc5k/EQXTpjaY7EFB47swCnaOEPXVpgRqjJ/Y0AlTE+/M
ree/mYWWdTH5m/uQAv5G2d3qGIULr6HUAaMr4qaOcd2THyowdE0/2TptteSwKYqsWYL4+hYdp3cE
uADN/9vkD6yY04I7/ohQzg9nr8EKp8keAftz3M6Y2hFi9f5xYVYlugNI+2ENGf7ZZrTTPUwo+sJ6
u9dp8e7uClHA/9k+rqKUMdrmVxKP9nok89O1WAX/8HWxOE3xErxg/rrBJy0ApygYIBUH6ewiF0k8
TQmi3v+YNXofzQfbgaiDMAeQC82zFGfLUVWRZG4hWpAd5rZZjoitAZhoNZ/L89N84J4Z7ODM7ipk
EZHcuG2LjeiAJiSljGlJSF4MZKPJ8QUuIKj6ox58h835QcJUhnkiddJHji8xUr0nMWKLvoi6gLJ9
sx+MnDLOvRDxiSG1c3nqgyO7nRSqA1TGO4Wb/7KVI6ldGgFLH00RGtKg2d3d6zdfgstnNKnovFM9
BkIc1byfy4MaWl0A2aDZXfMUMG9npJHuNJEHX2aDX3TICkibNtfEgddRvsHNUUpHH5hNa6sEMeh3
4jMKZofG62xJXh+lsQaBtswVW8UGqaDy37Z61CSznC+hYx/LJTJeQbkrgHeYQ2C0SibjbxqWmPD6
oOhar0bdsm/YKLG7pKHegRZFnte3IdqEvPGKE6DagN5OPAKwQHdfiamdYOLV1sHtafsr81J7NjSA
pQEWkGIZzZ4J1oqbK3Rh1fLhrFT6fZ3CMvEXAqD9l1RVomqXPr7zykq2Li+F+gpVYMS9AXOQBAgy
RdUS+LyDb3F+TD9yKBBb2NGEjbFLSKvtYIirOQZraZvcWp6l2T3k9QNYjdYiuLn+93WCFK0k/5PU
sjejYvG7X+pvIPL5JPAEvL0dHtXT9UYo3e0UOk7lizkqm2nYT9beJW4vRmmO2D1qw9o1knptt52P
SCOe26We7V7yZeXrc64s5ROyJADDVICG8rawLJZI1L5EUS8jGngcm48l5T7SeSHstkU85ssAz+6Y
A2axKl4Xs/kvhxzqDSco7E5WofqplZ1NfU9ADRvctPbNFp96V2nVKKEU6SzH71YNsE5TU57TdAX7
NR5ldd3U+yCx6rcFVuVdlhKhtxETylqs5kiuF7S0Li0uDMrYZ5gzfnOdSqaObiV1Cf/Qd+mFaklX
QKMaNIihfTFNGc/YhQ8JyRnRwW0o5MTGqnkzsQTJIVji7ViAseuUA7T5pcs6SW6Nt5MT4pZEB1IZ
d1CsHhQB9xyIVcSFIgdd5N49lNkjkmiFeOuEWUi4RIVuyzSNKuZpUga8UOnqGwDckfSTPA7vLX0B
51zTBMpQC5ncAMM1/LtIh+nkjGAfZj6spvaCzj/zP/dYxUMw23NDvnyahbZ0pLtMWu04uUeWwD+C
4n8W1TjydFp0hFBl1tT6kuTXnu6ruyKwKOJsuVkbGieTerks6tlSAQTE1iDlBeJdoRsoZuQ7fmSy
BDAoHdrSvdmC4K2fJOKibOaMEtH1dptRaOOZJP67WA5hX/WWr4VdxtMOtknsBhzEXjqZ8U9hHzWH
Y1gymY80al8IvbjsNaXsjUfaOnIzwxHfBCs/biXsy5s0WmEhZ4HsPp6sMUlwqLe4Ed53LdI2/1UH
6IrtS36uoqtuKNCpZ4wEl1gnZFV66xQQJRpyep8IedWw1Vu9xrWxPrxuHQoFotKtPuiRi6C1zlSP
pPQ0Ac9p0FKgRY7/A4gNE8j09I8wbbFqO4DIJSLVzg5ZqHHH5V1VmoA/lQZL0BxK0+OJc/pAXo5W
LLyg2dc4GAMrJU4A1XE4ADM4YYdaY3K62+Bm3r4r3Xz1xwBrdp66tsadvmBLqi0a7HZSTJ+lo3Vl
KATbOGHnkzIqh2In8vXIOZj94MBNdNKGsA6KTrlXo6CGybxv+3Fih+M3Z4xM5bFbW736Uvo3hKHq
7oA0w2Q4SsRyxVSGRJGLxS5coElPNZ/n7rxAhrhtSEVPklFsw3jit55/BTaFHfHyCUGLY5UpObaB
tB2glfjbQ0lElNhaSPhPLzH7qcjggSMqlLEPafalWFLpB/EO2hrs5dsWvj1GrjEd+nF+BH95tMcF
h+h+7sjDudv45ZfVdYm2e/bRYUPXCuNPq2/QILvjDadt9YCmPkjxXtzPICBATJfGbBzG1obe1zVE
V+QgwHM4ZhsoF9K2p3J311Hsynkv4YXfXFgAdSct9+fckrKqt2BQBOyZnPaCAOYoMrdG0/ZzE8HM
KBnGGTl5z2k8g/7gvv2gFT3iLhAx9k5QN4yybnTY034+fdGPYeqwsV8ddCw8pamES2JWio3Gp6tT
tFMPIQLs02YSgBq1om81vMggZLebKWj7KSIyZ2pAI/rJJHbUxSaNcHx8sPIgNPWJQ7ubVjpd5hIo
o0b3swMhIdjSFqobwxai5FqXV7dRu0DWIcXZ52LN/APo/Qx2E0/P+JsFoTLDQr45nAuapCYPawCE
ANjI9G6W3U9w5zrIZNpfi8qmYLXavpDicwnkNnopqSjbt2oOInaUle0dgq36GxCfVhfDUbuUPQDz
FwTXlzMcCNDwV+xQPjreGx5E2kZ9eZoPXo3cD+9oW5S+2h2cu9Ogt8s7LcRsIf40+sCmpVJtFYS8
EQpWPQelMjsyqvxkervH5awiilNSVK7dhkqjXu/4wIq2NewBkuUafJ/NChQH0deTcODmOwYv2LRk
O6xjMlQkrWy++ZcUsli+IXvJhbsTemu1u23K/qI9jYJgacxHE1KAuw7qaba3/AlNmfVla0agjART
Zx9ns1zwqX0iZoRgZ89NyYMcGC4cuJlTLIabm4X2/uHeA2tP3+27bchQafGn+X74GCHhNPSNMtRQ
YYqPMAhTlv6Dn7/3C7UmD9jQCfFjZaj0oMTToIH8uzLqlE7r5ak03zZq0bp4OZ0LKvRCkjmZNn6q
L5r/u30AMbo7+8Uv9H0RTvDBamt4ZOv5OKyf5NhYEN8iZgW8FwnffuyYkxNmeYfjS3vNjJ/B/dgM
SFDiJ0GSZCsV9frq3RDsOuLncWGUbwEQ69526YlahtpLcePoYbN1dSA2tY2c7SAbRSvxv8G4wVDG
EpXNtRZIL6Bh8ZKjqVlDq3+GMhcqz9Bd5mT05Ofpa+FEommoDBtoyp2eSEIB/wW/9F8PO7wT8gLo
FLUd9YlE91moX7v5Z8ex6hKeQh+4Ojo4RIeUSipqDaoqahTMC9DsJG7s0EhHQ0CbdbLooB7xOkw4
+B7y7KnGsHDY05oYy2eSZdIAGgWFfmdSoP0ElNAQcJAq41E9wmjih75BuniEhpIVlKhVkhFBC0qh
e5b6hQl/fXxLMuKeIoFjqw95tt38a7xKzaLBedOoTaPfY/TOVVgxmAsEc2nYjohM6xjZjRhBFtTJ
MFrKWKqSVIHaMqMriXrCSPOQtaHWs2XUOC1UcBc7gftIFmjeQ8poHhl4UhJuKpINV7/5fmyUIebB
ywajdx+VJUF6MvZsCel6gDSBzlLaVVaaCLaNJyRFeeiit5ViqA+Cnu0tQHUV+9sfvKEjEb2o3OOe
zY1hDGjgWpc3QE3+FAagOp5uV/4aW75lQczZnDFoPvS0iUd7lT3n0cYlS21r7OEFFP4/CNCOJ+6S
RSPt/KLFsX68VJzKyKuE6E/iOg2JnqhKb4Iveiu+VmYQUYyu5Vs8RY8/RWlyzKRpMaQrQTEMW1Nd
hhkX0/Vlj30Krz7dP/AwpGWtbLRTkEqaWn2KJaYCGQIn+tRZMiLrmv713NR5rtcZ1irzTfFGy3jO
zHT8PJ28rl6Os6YcVHC6lILZvuwOxbxfyt0TZ+Y7dmPmZgdgaJvlOBfUTBoT0b/8fWbCAP8pbfop
XCxTr2SlBpw0H0WarSc0O2a1F7xqALcfC3NOwnWWAcIugR5/XEeuUK6QNzre8o+dR3lP8uRmlua6
g2c1KVD7DCyDNVEvZqv10LqRtwirS0QlZliCZPjUy07/GVqpYsJcrCWVpsPNVwP5zVH1HQjuGVAU
xV3PbaPSns2vhdn/2x4zxUgg/bBNUnB4sP/c6Z51chLgS2igUZKsVeeY1ovh4xS56hovPHKFzlXn
xNtclA5sMm+Y8qepQV697sIJ1ofRlTUhDzydIamzI21HfWQakno4kXcJisUzPQpDjzNV7dIHboK0
iEDKedipQD1v3/Jaemn4JT7UAYdLsRMHsI2Jm68ndc01A74T2Ht/nHkyHMNcc7CjKX9OQYwMvLnq
MGp+ZKo65uOG258bsbkRUrtRuNYkaaES0hIFUjSSvk/aGoQ5or5kDoU5i107WKaCrT7iQODhBKHU
WHYZYipmDk4Pqrwuc22jcpGqiXjopcRFspcyCredVfzGgXrkbu49OHLQP+aPDs1ZYQ3yXGh9NBOv
egw2xjiwd4Vg7fUqmCMQNpLlINjk3P0R7GpmCwoYxUiAmvQZI8umphVus8sG/JrDfboZA0XEDHmW
1P/EpspG0G//EpIe3DL8a7jLhKFn8nwzckdmbMLqI0t7GBtKABDfJdoNcNGXjK5npuTZ5xOeuXFI
nZnj5ipcCORRljCvEkWvHZWrADPhICXCkIcgNrHrX44jAGKPmRTwUMQkFAVm6xVtVkBnuX0IJ8ji
L4f1Wz+2WbpaKB8qOTNVnrOfjUPGF2IYT6Tr94drZnM4HyuHCldyedbFb3WS6Hekkyk7CCLTwI20
0HQuAc7tHn35q91ZtE7yRDczFZz+B3q1U1Jv5I7UpC+y0+lmmitFBLDMkaur/2aE+moEW8omF9s8
u97yj0T9Ct8KmLmYGoHkhzk1f4LJ9vLLGa1H5VoiHTiWRGsii48byFm6ykdAiP1/YIBG5m7riiJq
2ey47y38fOLWsUcr2Lv8VtCOtYpqPl9k7m7O/oaM0jOSpDqn7fRtfgUbH2OZV0y/wmRAM3a4X/I/
UdGGoD7WlGhnGW16NZ5FRbYCSpb1e0d2t0lTxveW7UgGUuhN6Ozlko3ux6EcfTxYxaaPSQtYGlmX
7ni/xXLfssSqq5EYGtEMrH812kVfdQzoP9kHYbKtoZ4KL5d93H2ecV16tuvZUqw3RsFV9ZNVY7wq
RwVcte8sfXxCHbaegfPpIxu6pkQpNOt1kvtaz/rl4OadKn9DIU1tzafOeCfxtZsEO5AAyDAhrzMI
eSQMMmzRGMw2XOtccQD71X6hK9/fPyf4Yt+x0dB/1PT65ROHQiGP/egsxErKu0MC/bjgHgNyYHW8
S2uGnYTStGw8SEzdyWS/jZvFNagPVFipd/6elisT6H/uGzIFeki1cfzT61l5tw7iLNwA8Kph8J5/
3vImu+25oEr1a6ZqHeGhoCaWV895gAHss+RdFmbnB7nJjMfI23qpUJntCvUw5K27Fau8SDwutIOc
vL5DGoPnp5EuaWicTNV7yb9FCVmVClTHidcb0B2/NvMvZsmHaCiFBVqdmmPkA9V5cmaT7OFhUMfs
X69Fek2ue35eVnoCrVNc428W5YYDb7/EpjNiyXgZX9YhcS5h7p2mgI21BGaykt3H79qeffWCvPxs
uPCTYTY5dKDaMk6Cy9Pk9s1rrsmI3WE3z5s91Wqdp3pl5I5WgTj9OVrgewCKVnZHR4sS/Tgfb9fq
B4IboCr6YfNWTNtwAYl3Wl+2Iw1xsAT5kaD+1bKLAZfYs63DyOVw2rEHES0zFaOzGDSyABk9CDGU
+EhvUjdGPV7gXXaql5OyRTC5tEKJZafZAfdyGveaHYBQqPe2Rmw/uRmRDuMSXxYMUks690rMzx+F
Jt4HDysuota1kgRru3BHN+89lhDHu5DVxD28BSc8yZY5XfVO9MmNEx1fxinZdhokkXyayBGbvWqm
TgcdzaKc2BNWZFHU9+ypWUjy8ywthnfT44FccymxIfC1jFibiJqHfivkP2T9Pah2BD5P/ysES55/
PQdbbzPNfg8NjnxGXXoDdgDFgkCvBQ59mzceiuN3rHkQy2kzgzT95c+zVXA4nprR159mwetcj42p
sTD3vCYdob+TR9s5jxni5OblvsVPzcCP2FukHTpmcRCIsfryLe3Gt+pnkmse4RpfCWRcRZjYZelM
JM7wrEQNAZq8kS44jugeYiO8kicUddJNTkkGr3dZQe3NWNXlMDC/NdIm3Xil4CxHmtjKCRjrjCTJ
6cqAYmO8SAaCWKSUKOEH7wE6Zo7xL+7JcJMKhT/yN31ihpOWRvM8mjEtUidoMuZb4P1s0s2E/23P
yTupfbniXn/dw0SBaT04lZsU6Rr3OkJIchLimfQEUcI/7ktNBnzZEWYIcwgan9G1U/13LW7S+DjK
liv9Z83vYgBzUBv/LjQF16XziyAcNGXK/6JVkso/Y2+MPP0LzYs8wJbNlIO6G0TlhUFf8llQsX/L
Sg4uajTjHpThS8a0EZRAOPj++a1hDyANcT5pQNCBHDA7FrccCcoAGnwRYLmdmzdrEshIbE8VtfmV
7czyFb/CoK8j9dkrafDnQio8bebQenc0VYBzHJDcAY3DukW5/Q9dzLbKJeaAs3GB7hQodj1fgQIb
FSrM+QMOfowHPmokR5MP0R+tga3XqUL8gIvBOOErxHzeNOK2daDi4h+n+Ooi7OOYoAe0XKrSeuTM
Z1cFRjk8rhHx5A5iiDO6HVW6RqMnXlgKNiLkhlDI2bQvnGtO5gU+S6Pte0cKviVqXG0bTfDU5/oy
PWFVjcn+hX2KW1Eu2e3YtKMK71ox+eRYKyisUYbHMC+cFysz8BCz62QK2WWEDNR+iNrz2lUsDea1
OX8JlPunUHddziaQIUdVzkSF7aD0v7RLifVgKrOhkT9XD/971uBftVniy/4yaSbL6DOkY+wwwXN1
mLT3GL8tqAg/9jd0QtL18CqaSqtSTADQtrgXUUIlOy/hSU4Sz1PHA9NeMxEADVaxJBWyFKCFl87N
zC+AtuqL4QoPNcAAdRrlCrh/+2ZG0XqA1FCWeFHf8xeLWCu+iWAGW/kDqzF7pqDjgcWBvVlMhDMO
64CSTiLvEY65A0hBlt4TkiR4pcJp1LQj27QpQjNVN+qcN9MhR19qgNbvUF0m1whwVuCq2UNqHXT0
ujMoCJ7wZdsD0cnk96ekL9WG6R4eOjJr4zxAJawF33rH3lPCJDrOcYeOkC+eL85E62PMFBQuzBdb
1Yq5S6jnVNY2uI13q4FW9TJ4ehDKrC/9LfBVLfnXIduqMBiWG6rGHz1rkqh46iXgForwWPWzDgvf
JazEZhR40vQgKPECMYwYn4zyogMLpZQWscUx4gSmvqBk8JClT5eyMTar/oKcUdLBqZr+oXg7nsu2
cJ1OHWCHRWOurybeLmT+0qQ34VDd4NCerYCMcX1zLEOUicMbkrkNEmlKRQkVZpnMKRd2GETL7Y5P
xlR3tMrCTYazlV6C+TjvzdDHf0SxE4Bme1q8IgSZa7NqfXRFeAL4DBDxDMdAFNuvuRnk1pPsSg1r
+ABLwqt1jsUxkedSwGJoF1KSBBiu1DSbqUMg4pBSWffGdfBSyoUWTG2NBXIUcFZRE9XF2g1+gY8a
Y+K5s8ZzVYhyRGTLNMnwHYGIUD3OMZBd7wpcraNR1hOFMTKKzXvkD1zmfD0JUtil/Sm+eA2+YV8F
sz3Wy7efmClJ3agniYTrKaJXfUYEqfAwhqq5130UxnuxlmPO+tYg+vF51x9kWMLKHyC8cuKPH2B8
4LB687il0zDnUQTJzatfz0WUU6Kb6pCp7zUrSWPx8NURjaz/RgzllemR0vyDqS63mB9oV1Ud6LwO
JQa+qNVXxpyeiaEW0r5z56ZRzZD2RX5QdX1SdzFNDH9rAXaHHacQvuxjZMmMbcIxdZZ8mUrsxASp
ryDBK16OFNer96wJLr7Sp8qLrS4uvCDupQbO1KRLjVlzgYPYxJ4WT20fEgVsXRRSMTgtm+HHlArF
Q4o0/5PJYMw/c60uUftDNgk10fx7Gov5n7JFi9soqEhOWZJvKxFzTzfVmkOqfGplsLsnlFOMHsuk
TDop09AJ7BKLxgy8U73Ctv604ZA42O1gU5bdAohEnPr3JJ9ST4PUbGtUmp6nWJkjXujpL3qwzXha
v68Jl+hu0u0uKlq78z0aKcsJL2ukTHJKZHLFHhTINO+Tuqeqw10WVQFyk6Y6f05WejpjANRfIwBU
PiEKegcA1uQEE8XJtX5T4YUjs0nrePQbc7VAtPxEJrTXhWcNeZbfZ1pq0V+HlEajP3ACWKm/0+wP
dI+PvhDdqheW4UY000uUir9nKPKjPIJLzYf5zNdwD6qswGyZA2cFixJNyRBJvvALftOgH4JZXgfn
mWAEC9gy3O5B0DVBqbxFlRrNlYjk1prXtefN73fmYJJjln7u7keMrZKhG7VPb0HXR+eD/CcEQFnw
dZJSeJChUQ5yY93fJSnm4M+jtk9TBpyXF4sRimXWNKBnFsHv2/ySV5VFbG6gVLolFwCiySVFzdsv
BFKmU7yh1YkBHCtqYYsClQgXmww3FJU1Ao5TGgakQzwQGeMtnmH4wmIvXTFlOri6sZsF9cyD9nal
8wBG3RoUZhTnwsD8BMiI8fIj29NtL8gVWm6UxzfcMaH7+qYv3zJ8vteJl+xHTrsKz/RojiTUUloA
dW4zgMVFoy4s+IfiQansmyQauqpZiSvTDlFE1mEWC6mJYwNQNV3jTCYAopV40K1ntQP2uLR96fRk
DlN5Zqyu0FUsEfZBG4d+Ly59eb8SlpUBuWRMDkoLlxCkJB5eO57iJoZa8lM6e0d9JGhCRbAgPzuP
XXhhlFkPHdicHkN0LFpXQlJ0jqvJyBlIdA3bcM5Stt2GxSR1KbOsaV6u6rWXvfuF1Htd4Hb+JN2o
X7kaD0KYA2R591n+5A71v8LsXO0q7Gr6vIlkEGzZIYsUMOoJXsMQ0JEaslT7mqV0T+oMtMOsWk4Y
Vgc0Hr+RDRfLXgyuWGy2EDCNTUgVCZ7F/SQnSPsbjNsLVPOeA6ZHZpLgc5i+KMdD7WJb0Uzsu5X0
Wkrzz6fzPn11hFXX7zp2qxLx1JQhIiUegcvNFk3Sgxm5i6jl7CxgmDWyGTla8meAlkuwjQtAAeIa
wr3hk25x1gmH0cmd5SJOce85hgExOMOkYQ1TCjNdihWKbrWXDWxPc6GUpRppwELK5GuO20q8jsfQ
lhaw12lN4dKZa7XY/YbWFUaQ6Axgz76wcSCNXN4xWRdCZX5orBtZS20ZjswZbNsZi44EV7yQ+v47
Z9D1sqVSvQRapqk47d6D5IMwufSSS50KaMq8avbXJa0jHnqW5ozn1jNXog07oaBlHhBvqa5hfXhT
eiREntZu+Kt+mgGVVSBhi6V+gtvI9y1kbkauhoIa2PHce3dn/97PolDcJ+Q8O9FhnuhIL5/IHrUm
TErF189n0En6boWEhTYrcLvIZ6UTpcemmrMVTAPumUNgXcbLyaiu8wuisJSB9IQkFz++YBaHxEw2
ZKcJqzts+XCQxRshTLF1ywndmuBlBBObkV6O4KrwhiUUvBC+AhPa5YlsrPbTc9KVNRpSTMoBhuhC
Ir0NbsKg3gXgibPUb41pkND6GyCoMeDYSANlUg55zPQkWpGaCBaxokg6LjGLlNcCvkTwijnwZjPS
N0zZ6GIFSscudOGCnUh/V087AUR44ZDGDwZeqoWMIyZJTMaR2B0dOSt/wjeca3Hum5pkFD/yJTw6
wpu0sPI8BoUy+N+bzZJTdTZtJXap0rWVoLR4I0tec4gvD3vyZk+c2fciv2E29gXvHefHwgcdySxg
1cW3Y2LEczzBYq9QC7FYDtYDNeE3NrxL70O9CXThqtb+4UkgP/5Rcsb2kB8aN+/fDuRuG1NQEtdP
+HOT1vnIlBZA4yDmW+ovAdb5t+MvIgF93ts8nf/ke7VXqzUEXHV5aB9TpfNpCHHTGzHlaieM3qu1
Wcari8Bssp9r4TQhVgPI3NqeXXou8SBatAb4OeE0oHrgPHkvTYoyO3XmRugRTa6B0UYVtOCSIuKP
AyGvnLqitN3NMtpnZgQrBkjo51tM9QM/RG74NqbrnFRmcrVam6BDMQSxeWH3Pj361VYq9OduB9Y2
jkP+3RCRuqycP6mhHJe8LuRywtBAegQBJBDk5/u3ks2m7VnLs//R2oBM+rQFqxA/2E4ATJw+8rDR
QnF7pwh0amv9fmNnJYAJGiPQwuN8fW+uefQKp9y5mMflmT4AajVDq3mYC9DtA9gCG3qneaBFDm7e
TaOW/SwA4D5wsW1cxzHkpHZ8yEmOWpXdhZU/vT4/pZmhv3bOVw7BCK4pHB4qQN2XbJpakwrcvV/i
xpgwgZd1jrSDVARwcF/Mia4xp5jWKRJSxYTU2h3hi8Qj50m+gJKxFESn8HX+xfhFBKAuUBRureyL
Rz8QDzn0Bf8bmdkv4xk8Z0M6sgWjZYXytulSK/W8RJBXOoqpqPeHSweXnl9Wet8IZnIUBI12sfMA
XYs6AqPowEc/KD14RaJthwY0nEZFCLeqoHU1qW4cMTiJJMmZsWrhpc2pCOd4ipLowIvHqDhg+rCg
upgSsJSBwoLvUins/607LjvHNM3ykXEtZMNxbcimvDFqx3aC9mA0ViN8bUSVLSOb3bapSeOb66ej
1PRL+fYxmfELbwjsWCQ2jAmQrtULyVAtB/LVIzzYmbpOX5FbHEEVp40yU84k13/hEQapwp1ECjhc
sJ+T5R3knKKrRyBTirl1+0uT7pO2ls2FYVA4MRkr983nml9Bt6O4Jr1/cn6jqKE+UCQYgOAg/KzD
YTnKjaOR5MppPkOOcPTFcYGDvpJrtCYqoByhRn3YzMhOeCC+hxmrgxq3prxk0OtVFbBlBq9iBHoU
19QkA1Bd9SWzWiaFY4nldHQ+9+xNKp5NpbLSos4LbW14UNVx2/JcLivxfsPiVUaanyFw2PHYoGtW
ljZfG8A1t0lExANFMD7vvVQ2xuc8ozJPTAuLiYmUzlGx9zXzJgrCLwiIbWopgT7nhkJDenwptGEM
CZf1ffetlNs9331D01mN2Vsp4TxBwe0oZpU7waMinL1R1XVGHP/fYlhvm2L+gmmEE8DQHV9ZhXwk
fXxfn28C1mIEOqrGvxzmWBbNX9UCWyfgDiqF9u6z6GQjcFwb1vkTCn2B2vvlPeNzPQgfjrx7bIbL
akpXu0CrbldXcpyyyKycmJCVIagld2plgrYxHYk+BQ8RUv1qxP7q7tEH6EhSKu7CdGjVxNByEY7d
3eD/D89Gv+tC7BEovAzKlYvFTCwFcTneo9Wo8jy7EWaPzMfjNUPftW2pF2fC/vyAnC9v2iZKGZsA
6DNUYJHE0+8A8IHGiS78pqsTKCxeMZtqRrI5XO6YmAgAhpUCwJJPkZFvVllkwC2OUyLJKJyN5kiv
sD5kB35gnLVdLRqnpajj5NQ2zWoTSVpXqRBbAgoKxAcLX1m8LCZ3XSUyFYWVvBgc3ciKRpp8wYGJ
Ywq7uzq93qT2ftfb31IFZU7w1RN1BnjJJkY6HQqAC6haEsI1SEanH0UZ2OUL7f/YWC0+zDK/D354
YNTvxNbJIM/NXRoMDPTg0b+oNDa+eitfRO5utoaSlZyTvW2GzbqWcCQomvyuIXeRePA3uBivAgD2
ocx9WG6XI9RJHUabKb5yvKkVDQoIVW56wMFS0clOKr4yCJO1YkH0kJHG33sycbWMNzQ4Q6HPIeUS
dcL+6xFNcX2jssOKybz0T62rrqrzSacXayDxvMZIHxdtsB0sjS7X+Xc3LR2sRthoElVsOzgHoeYD
0PCRh+4xz39y4DRCgSgT3a0GdVeg937RNlmRsAdTwqCZfi3RTGhJpfggYaZ/xIsWi7TFrYOqpr/R
JEoHZj1Zs+sLG8Me8EH7XYg/4ILHDsPU0iP7blxL3ce+OHWeIcOFSfL5TILulUoo2LUKGqMinoDU
tiOGcT8hXq94SsYBiMWMU2TuplT5irXGIjMPQkmBBOIWIy6T440Hp+T4OlQwK03sC3SGH2/jLd5p
cSEff3ubFfAlRMjdQa8N/VCCdwUmf91rffOxS+M8GGKrEO8wLLr59t56baluuKEI85xk5MR2HWOD
+VaXXumBx4QkbJk8FUstJd23TJIDkxwOw/LiA8OAIVaQhoEHONwEVcKs2qF/COHyIoqbkzgXDYBw
set/9iNI3deN0mowCViYUhJ2W3Oy6w6aMxY0C8hFc3XlO0OJg1PLCIwgDlKLSFJZ+AkED/XzLzXJ
1mSu6itPxrs3Q3qpYJ6jtYlntivDaioaAK/zOuuA0LcQtpaundrzwrnKnIIYqKMGwJmGabmYeCUc
pFkugopbwHcZ6ve6VCrEQssR2KBCFo6pbk/njSCg1cVHXT7GPI2u9+bQEg/hW8lq4mexsZQk3Pgc
vMYkg5Y1LKCf4jVscKQLlK5YKbs5vRCdU8AHYTeAdeH3aNarXyt/ATQa423Bm3IZHDOiM40x4ivJ
yMjlZlg+TPLb+2oSG8icYVmopCJQot2AhtZeIWEGWOXiDqW7ZanNWPwF1frSQyyGu8j2d23/P2IW
9bAQbU+d5+aZ5OVlG5FJrkPjKWeh/X6QFfeeBTuicLgoVa+EcMum04viwPDQcCnOC7wZgWDn/6EV
d5zrkZsGTRO9O1MnqDkqvhfWYSO6R1Ba0V6oSpHw3tGGzikzpyzEWCJt+84R9lmfs7O+IjWs79eS
wXoZYGzBpfhIkPcAwgCmVAG5j22jOCTSYLMTpNl1sK3gfU+J8TK8pF5AzDVtrleOskCogSp30fk2
uOnitQWeIkC0RRenGsHWrmKNtF1X83z1nukmaaodEsfUqzOhdmQ3p5J9o4ha5iN/z80QH7WgaytL
s3eMgG4vGBfOt0XF9EvcmNBk/IyEcY9WspcUSXOE/kHDTtqzbjuRw71BJNXbtn4Jc/jap+IjRYza
wamSSoQqztX0QuktMF942yGvTnmF3CtTvdJgvSluA+zk55nZ59JAe6l9REwUYZ/kRR1RsN9/o1wY
1pAHIE8ZY1FouYJ+YSbedEvgHFsIJIhWvI6Lp3POcD/rtckHnKS7zszGetNYg9CyJ29ZPH4hf7Zg
ltCVoOPp0FIWRr78VkVNj+HJKPZFaVAjtBqrq7ONmnguHmVqvPZvsSBzQy9arfwKAHxOIi+sZaCA
4L8bDe1ZEwj4UET+OrH3FJuaSbljiUUX+dwZKV7vSawHUOxEmmizPZ+BN+5OHXq+BdApyIgXDUK9
9I0XxmwlrJkKfaH+kExJ8zU+hHvU0MOGed3ANPUo3tqrWy6ed7F9swiRHVyWQfkhbea5avKae4Ne
PDhgKmMLLursr8IXIedt2OXHKDo9y/x+YFZlS9QMRG8e5/jVRxNdRRI/XXZ/uZ0mobwPm6gRJ0Dy
3/byc8OI//pjwcpimABPDQNDAnIvHpURBv1xaA/669Se8w6WITmZHvwgbUs4WHrZwUbwfUd7QhHf
9rebJydvislOSahcyB8zBRyrF7RXAZIAJmBw2g097ZntZI3TYU9lX1IxFHZW5oC/M6+dBMHDB+/F
LqKT9yxKBJ+bxrweWQxyHvKuwwmAdOxJ7JLsxP620HvMKcedS4Vd0nnew3eWKAHRg6DRBLWMC4PH
y3nVX7IKG3gt4xmKlw3YyJDz/Nrq0yEwmjQ5P7FZDF4QEyZMdNI5dWkGERWVJpAED/5enrZjbvza
fWiR8mwBkV7Q/Hcvm9pU07f0Lk/4hAkpf62euv8Cg//e2SSRvx5cC4uqtMauCZs54w9nfozIfdfr
yH4DojinMMd5Un6ZiJhetHq0P8pv14LbTwJUgJNcU5O+GK3KKJ9Vv0qV+aE5m6+1oZ8EjowfvQP1
pVSA+08BcuVC1YlZA0FiJRj464vqGH0dvwokylOJN6g2WR92e2HuzOPNyJMvXupAKpym0vmNuWZk
OUJKQYTrwKAxKPYKT7alTQ2kgQJ0EElsrF43mTESn+W3vu83sbYLL1kROj13Jrd6sqMWpoWcZ0Fz
bfrep0AJO8baZfl3dAb9960c0UxeVH0P0r9EWci0XXLRMLpwk9iJHs6PZ0WobqRmfq//YXBCxdVt
bn0NyqVjFbEBqYTX/93Z7Ca6pmd04xCDAPYbdZvbHoTABMjyQNQe0GQSzWD4EUxUrfshvHB3lcGZ
+oFhVuI3gHkeYbve2F24DOQ5C9rRZ1kBuqNalILjJ5KTm7MydKY7uFQaMqyhoZ3zUR8JCzW+aJJP
uid2iZzs08OTpcH5BK+c9wwsxlkwunyCORg58EDXsWxnmeOKbkoOp8ilzP1QmX+J8hxc5Eh6yycs
eLoOUCcGmkUldp/qKvHPJkc4K1KoxvB7VtPAZQOezE1MhWATlj9jeM9t4XTF8urh3/hVXneZWfEc
dqcfunUeIec0nUqfPXIX4SaAyhmcttguMlsArDNlJrI1WUpMlIAbizfZgdV2sWNau3SaOYuAnIpf
YKDTlog7g+GaD+j5moVPIpcOV7w+ZaIsKP1uLtPOkXQqbsWCbZt85ky28OJQsuPX+PBc/Wq1Apx1
g2vjSTkrR+clIV+R1WV6EN5DBJMj7VrwsLWzaMV9MO/jh4HxRCFO28lsl7+buqaXzZDHQ4I2iSAz
Ggr+0EezlgGIBn19gKbgC2qeOBhK84Yqn0WksJHkE7xZnjtl5e0kaXldiSfMLeb4BeTxSiBevNos
cNGvWcJRwPsy17oogocd7w5FX61ijFT+Pc4oxF1pJrYhHGNeR7DzR1ukYR8iI3qN4sEsf/S6VlfT
TFkAGs9lGDZJdnMmahaU7KW+8g8g6JCGo/1EOCUJR++N5I7ooJ+ixCzkFnx4SxCIRnVYDLGJsceS
RdkMV+/Tsrzfowyn/6OfAFlYLWYz3JufxRZJRQQCff2Bav7vrLe98jRf++sVBtjXAIyQH/qun/09
QeLB7LfXQATaf2WTPznXPUWy/vhPHC2xf1TtEzKzjIOy0mC+7UR2zRMLqZWE5j9SGnnjU/he3aZJ
qEQFVEpK/2CWvezPq92/9MYL66EBBdWUFyw5FIx2Jil0/7SFa8PAwCjmekxrr79o4lmYhIqm681z
fGUYJSLOtuL+RnguhcYYqHsPnrRr0vSsIOLdFwU1/lP/K90Wfm71zITxEQJxGtlE0+1hHIbBV6td
s74D3bY9QkgeSd8kepIngSUAvVrLXEbFU1tx/naeWPq/MFQydOO0YMvj+TqG/9awz2NlLbUwYEjB
Gy/tAj2ilHqFO02eNEhPWWnJ8XqQeIou4UMq0GOTqW452hzfMBkmxHlNmDOGhbJEhc7WPahzdApE
zqFO0pv8etdSip5yNuUgl/7coGT+Z+NMx7GZ/r6H5jMo4US3vBoJAOiTs1dCg1zGT8Ty0tBcsVLo
orGMyITNPSoXr7q1fOS8YglTvuVDlInrlTWtrBfBmUUj0heDlZHu3DBfU6B19e4Fz1pBQc3jUjez
H14LW1Xd4bCCKHL3qu1Xbm58dfMUQwXKLRXenJiyffpZY/KnPNIreDWfbtOBzN2/iDfLfH+QTP++
xR6PHn9RUuxJ4KLAfWG7vAZFwXDIItOcrbezod53L24XUkrtvYj3uSydZnHAURRusQN+MUzkiBxk
8iZXYPTJN9Kop9RJPujnJT01PzHRSDESPdo4AGumsS0N0gHKr6f7AslSboG+TGlQyObg6j+WwYfl
XydvZiCmMfnz2hKpS0dmL14nSrz64U6SZhBBPGhr26VZR5lTwKrN0Vk4MmaqOXMW7ITUg/bWFTW5
dwD/+LqhEV61Q4zyDL1bPfzOcPxY3L96pbS2eb+pFJWjbzEkkweTq7dNYJJHvqV8rJEk5odAHxxo
YcEdVpubvZh+aUWKz5qjfYraugjSanGJOTCX1opMw91JgJPW3Q+zqjhjcVex4icmUMIDoRIpuLvU
7gxazD/1DKDgdv45TLniQ9Dq3TThYxOKWYy8QI+IxQgRCp8C9VTSYxO1bguQ5KFXF1d8P7aSaQJ8
D3Uapgqt6CyoMKCmHtIKI2SCG7ZPULWBSmcvDnpOxKYjTAurKwSg6Zq5/eGniaUHN2FoOd0MlVZA
eZSI4Cbh5/Ibm6yp6ofuiU9GiSb9l9Pnd4KTx9dhLFPgl9ZtXtc+I3Hqy5o/KBnPcPPArrglG23x
f1bUdAQ8YwpmLxHufyM3bKm0NkazreaUYcqU1cSmF6PipceYzXE090xZq7LTu4FplGSrI4ZywvQX
JKzAK4Qox+SCz/upUUg4FYGbtodNvcRKi+uu11ETtJWlfr6yZ5tCCjK34GtBImvdo1Fi0ja8mG30
b03lAZ1NduiyACcIRSWIFjmIhH/irYvXWM3t5VKTDEbxpqclv+ZZs9j+aYxA7M8kxmMvjJJEdbU3
M4I23aGPbw5x0mR8WiTgSTHsa3Nmwp1JkXJMC1TksiAYGe/Btx5iaadSg4H+/7wu3ay29q4vBx9S
rNKNZYZlAurgkk6BxMBQgi39dHrCg1QHnRPlY0MEYamLgUS/uNB8w4sobgTPa2p8D+bW/VG1GTbY
q0QQWQREyy6lEd7QpAvKw2Nub2i+h149lvWtBpo4F3z6gVziGH30sZI4dJxnbEKPW4IIqYi1qF3t
+dk9B6C4vnjCJQwlFg6//iy9QfUKyKhFNjlduKp8JZTh4iy5gd13i/LZp9JFC/S3JWQhnhlgNv+e
WaDYTlAj5bJh4Y17QtuaY41QsujpueHjoYLv3d8VoD2tsDJGmn1mPKWbkiBLA/fRDZcnQauapeQi
QogRXPP057JLQXWqzFFYsrG2df3DC9KG61M0TXjHG20t1T+64wj/AzndV49f4Ij3W2e2vBtQbQ61
Hgi3tFVzR8I+rkiiBPId4JvJmbyAbaDrVRDFjAyA/o+LG7aLIcGzYl4nIcrA02DdmpKL5mHwbWqR
YzZqy6k22fb2LD7tr0b/QuZ2KZChXcecNObsbplHAX5SJEUMLAFkc49vbcseBpmNbTBzK6FZ3OyY
Gu/XIh9TssPvP8Cl+nWwLVP8ENQ2pR/CWwK314KFqdhTtv5r4pqmgpx5mmwyvoT6SArqYGc/jgsc
i+FMTfion4u6JUEeSuaAH9SPjS6qJsOCXCBtjwvBOdJ9lXWo21D8Gn0AvSxTdORdiTX/Y1e4anGF
iklH9MC9/Y2AfkZe7cYwGUbs5uRUdLyPUJlbaw6aeBJeBzAXhws83fkOhrsNl8BeLDzY1dl/9ODk
I52xztvfSiU9pp6NtOP0YImQqjnCehbwfTE+8JBy8uV21elw7zHu7+BzHb6MjcOO4XsPant1BkL7
xwrEeMYXJMFn5Y64JgK+b3bjHMjQEZ5RApELy/c8s1Mu0AOusCUZSuR1B1ogaptnw9XjNgAPAbpZ
wM6UtKdcHyKGzO/PtcKdm2D9jt3nmszYbBlMwgjIyrUW2L34ODiApTmsWG4nxMJg8eZ6M/7EkMax
ZnpogNpIhgrcK+ougCEFgHiVWLo2D19y0Aig4rI0tviTdqVwmuHqMggu8RrAhGnTqluTwby6sA5h
p9lxVYPhKTzEc2JtcwDzjRbMSclrmmQep7iQZIGH9XS2BUMJSTvAQVr/fODpkTzc9yt2bcspAHFl
8P2RVmZsix5+gEOV6Eo3Mgawtf3s/oXcmrLrKV1dbhc1vhSe/9njpVfZgRJld3+iE8R1/Xi2K9gc
HUjdJsuBCryEPbSgvdfeMNLKZsbhHUHB8XcrL+ccK0F1AW7hAwwYVOogWa9XxGdv2//TR18PAhEw
XfVJRytFenYoyG+4ljGoXpXXKxeu/pD7TaTndU/Of8QoBPRM38kAPhe/bdo/MmAYRQ5TtzjMBTlF
GmKtG8H6CVPohdBtTM/WjKxoRHMjtG5+Y2WHMa1e0M8K+dMDxk1h/sYiWdijZE09z7eM3mg734MH
cSdPKEWjL279/2BTEzuOLLN8QXJslGuGk/yfUIO4+jXnw7xXfMcLLhG9HZrcdxFI9PtWBu3vx3TE
kdJRYu9tfjlDtOCFMe+0lPMUSoc8HxugGRT5y6L2+kB06Tmqmkqqcta1mOrOXr+/Im5FzmZIKbyg
XrDBX2PjZFtdz+76VMeE1p09xh/jz2+zpdhD5/yeoClHKmBAd10GYksWbH12XvHgY7+/tywiZ2dV
UvJzT2LJAHt0ECpYghYpEQVyrRBlOex862eaCCpi4CROxUQimt3HTlnnl+KCukcOHU0ZnVb+iHxI
7wgzOv6opNGfqQLTfS3Mbw5Nj7p6/7MCorwMTysDeqzgwIdcpw2EYnvSZXjciFEAeU1/V/e+SCbk
zWqmfFo/Ou7Sg1HItwqJeJgVfwJuzeGcqu77ovpDybFzxm8mzJBXmTcMorVwYkOhY01I8zn5rzGY
fhTt+JD3EQ6UFC2f1uFsHlVFJejX1egG8RyAyuqE0G9wX0rTFlgfd94EQs5KxSqjhuvcF2MXHJ1u
2gyowE0DSb2YKfuHfCHj4oxahgB+0tRfi+MWB7QhxS3ZWExTycrps1mqdqQUUVknF7Dv/ctl5Gol
H44+gBOCqxSaIl/H59dhaKLVq6P2EQuC6w+geZ9ldJCe8zXX/b8OaL7eLxiGzK7pSCtzZKz0z2Ls
VLI4DWEHDmfg0zv/AnnuerM2/TTPVGLJpYZx6/oT0RZFdjWQmxAKaA8sJUI9A8h1JfBgTBcntrd6
ExPai0fS/LdRXTUPQntLvFNC5UIiPh3LvjDoXcwPRLzoUrsi07K4Wx+55XPrqhX1fnqQM8OTju3U
fSfFAG58Dw/eKzRYQUKzVoOafiU3gzMOqSHhysVBWUyUUsJAafNnmYPrg+hjqeMLenH1m4wc0t2v
jn/+9NVIvsK12MOiIZW85/mVilAwaR257WfG1GuDddXeakVlrcVn/MlvxvfFqst2890c0nEH5SEb
MO5pOhJk6P15KA76cMsS3h72NTClYNdxL+aOH3u3rJcpKUNr/fJM1TelE8TrO5Wou2K3D6Al+9Kw
xbp2MJWqd50d+40JTFAiBfI6zD8RNd2HP9iBS8qS3YtUN3zHS4H1ykk+UH/98Vf1T45nkJ2mX/5v
mENov71CuT6H9yCaHY7A8X6fdOgjTkFTM5mNPIRVTpCNXTWSvKsM2CDth/oFKizpLxCicu1zm0X2
kvFFHsSz8NdfYjoY32Tldi7pnBI1mV5FiEpQsfazQvUzEy4YuTErLYM0bykm5/lqlAHHcmnDNECY
iuRR0fX3qhuZCtw1I994ixYCWV6mEr5fn/CR6nhH0tOar+Bod7SC6lH7BqeAdVNwz37EAbJte6nc
uInwWU4RXyruIoqXUYpfPimZB+0waLXqHVGCHT0e33GXyRxUUZxb3LLJP5Isuvo6fh5gBWbnLCcp
tRBcKJU3n0LESP2erVyr3pH2V0ttcziU+h4D4trh9uxf8vEUqxEihuudMGeATpBLgEagiqbb8NT1
LscmDPhkOWF+91MsF5gLNesLDNaylTXpHjqkbEJaEWIguuQWqvRtXTbS3Eh29g//TzOBahOQDpLr
ADQiV+8BXCie6ZcUVrntHOlvxedTvWJ7350eDLgSomnNC0akxtNlrapFkqx3d/rB7T3inM8/2X8s
2vNPih/QgfeHTR1k8afRJpZtFF5jXbu0ub3jtYX9t+/CVT/gJFNIBG08GqpOGCxt+IXvBQoz6qAY
g7QExZLQ/dNzJWfQbE6LLGPxONbDbbeSvhfomofnDc6U9wMUAOOr+jB1aRjm6X58fzlP40n7A1Fg
kzbiNjbXQILiszWQqsivUs/F+OWqjcYtGpyloB/K4XA5MfAScdufsrDEHrAgFC7D4WBZSjKsaReC
OeyfFPfyY5C1KZvof/tby6RlnVCDQzAP/xHgVrlvgCaBeDroiCA131b7yM476Nm7C7kcrnjCeR09
gOVcxnxZUyyOVF1dZ60nY/Nts/yN+p8ae95+aHiYuvzETGiQPJwR64RQ17VjAyx3C9jwKnboCm/B
s/d6vn3ZFLpXu3FoQdVpr5ohgWSdnaQPJJEGWt0W4LUyzbuJQnOLD6M1TN5iPKlBuI/sMIixqMMA
HXoFCy81r1qO53l82NawYuKy4F/76/pVcJgZTupImOLGxd9YRCN5LEIpn+iig+4jvxkx7/IkFP1w
JnjHlxiiDuST1IRCKdpYJfYjIvBpOehm8l//3RZ0HrKZWJBz+yqB6qBF06cQ3HrLbd9eT5nXb8bN
UIsbk1KxH3IKu8dh6E1nJ5wh0YrxmQP7OLr/jOT7vc1O4JjsQh6RsIUep2R33ebbhBKtxjbAi5Mu
9WgsyBZLrGFLIsHG77o/m2WMPfeBW2VZ+rk57DYR0P8ODG14yLCHWxrUgssbicvsCQpuWa2kl4ga
gZFWMQgt2RXN/VnzN/0GM2GQcdd55TR56Uw0HkhlvPGNrD19LBUkeh2J16UyPM4Ljfa0n+fdaZsV
iXrfXmocLuWrE5XyHQVp46VoZjTCHVme7TrKVJlwdbt7YBHV6ETtQDXwgqBlZrMTrLwMyMFsgyml
0j8WM1NoUfShXfJFGf7twpf8FD7/6mdbHxqqA1rEfn9YrTl9hBOsvpNirexIb3j63ObXHd8incjp
rAgFTlbWBbVgsaR+sm6NmwCd2mVwlE/k5SMJ0+b34MoSzklBB6r3hIVLJk4ec8lGwLQjDc2qIDDh
lrIhTHqndZ/UzPh+vVwgR/yyqs12R/r737dzLupL4jPYNh9+kKFMxalTQsqaHy/3KpUUOJxq4XGn
Hy4YyDkQ7vLFY9VLxYPccDy1DiG89eInhBynnBjJFlgKbZSYuRiKkW+BJMRQKdy4FlguwHVtAsaW
62X2N1NRY1q/fYGfJlJf/A4hFsO8PEYi6aN68tDUCHXRLEsD+N/VL/Gr3DrkWxUlRySCn3USxYH8
2oyKMgt26cYEzF7h6eRt7r5LAsUmAS+m19Sa8E1isegfC8lzzJuxtRMG5hPkharD4qk/7P9lP+mL
RbIzPCgVQEd+R2tdYKNW/Dg4J0gxA2hrlXn7W8F9ltw0gkyenmwYLxJMrM443RJh0v19gnfQXS/e
cE9BgxEe+h76+wxNIzvE1fpMIwKoYJCXaj2qFjONGELoottbzpuuCKc41YNMx9y82TFp2sGND1zh
dkf7TeebzbSr/m6+TbF3FnW17+gleVVDtHAGspJr+AqXn6c4hb8pVspc+WQJ9Y/QcEnVWyoSCYf6
bUlW5PKzhxFgRdKvtbO6damOjorYE7JnYFDOM9BX24VdB1FkNlXYDGSnBgXA58dlhKqXIPT+wr6Q
8T89msIIYL345i/y4516V1jqUajuN58oNPBd/BfTCKuPpE3MtEJIfl9qaU0I0tEfdnYSdE4MCevJ
nG6pn7x+9U0zHMWYEuKY8X9MAimyzd5sqFVz5qZAuf2VMfJTw+fRDQOuFARdaathxgKV4/pj7W3g
oxAPveeTVDFCPj6RKU/SQYtMEhvKxq1ypMfR6YhIoolKBRhjcYsH3N1V2F5CqbwNveHPmUY6DT0x
xfhFhkxYqCG7e6dqzl5CNAkYCi04UxR7X7JgY+d8Cih85F90nBMnNdt6B2RkZMYJNYrCkaVBwbPr
3jKjku67w3BqJlnbSwH56K86AE+LeGd5hS33QGvJiPWAbKbbGMb+7zoFqohG2pFJuoepJ0hcvTY0
wy7lKidrdjL+bx/jq3nVkST07Toatk74IQ6hsXg1CwmrXBfxn7txnmua4VRPBcPo8V8AKqTNbjGq
L7mSyMhFAlDUkLuZ8p8SPuiqlS4X46o1IGPxlA7OU9HVPLfPiq7M9hNrFcaem7hdY7R2AOBEGe0W
6M9K4qXBcYR2vZSrbvH2vJg4DGwJ63N1rIurafy+4/hrQVnMfeM1nhRf9gD1fiyy4CdGuN+AYybZ
qwSYWo9XhG7GS0uSr7tD5qSdferXuHXqWMiVXQVCN5Ob80vfnoTEMunJbwmb0qrE4b34lD2CgHBG
hpJhBSdtW+0C4mbbn4qWmqlt1aaFnkvhjDXey/6dEopELVoglbUEg4sdiflXXKjWSM+zYymMa+bh
4AnoKl4bw5iDEdXLLUv4z1vuNzopnZtdXxFU+bRyhQET2S5LeYP4cHkUNQTQfB4gxVb2t+ecpY4a
8TJFX1lP58hvyKPxewEEu368ND8qsxqzQs6sPmVRl/wRyhrVC+olJxcieMq5U+as7zhITXFQiY+4
ZPnp5FtwfVDvRAG1Rkh358izHZDIo9smPrhWLwcxpG6lo5cCNFlw/wPYGcsO7nNoVKUjfc+7FLd2
YopXX4ngVBRiLJiXA1m2nRJ4P64SMPIZZJXeDx5AYnTMXVk2vpg/+eS/wu0eRKMPYHw5BqTQWXEC
Me1HwZpuDzFnEf9f7qmmf24n827FOHlHPnWK6VnOoFHQd2oMW1EnqhaaX/0PUFn7gu1cZO8c2uWB
k7H8+6vfZLFmUqtEwT7YSKP4XB4pQ9DTiqS7yImQZEcTFKa80q2TYrGohshRoka2xH11GEhYGsKU
f5yWB2lux2ZQOBivsDkdo52w5voBVxwaD2zzjR2E4GJFYyuhW76afk6l620j8UevhuNbrkKL/+Ch
0szHifwNP9TiMvUtNLg9pI2yx1qKrnCdGzBNrWRXghmmHgmyHIYZEiF9i2EI3tzbBZX3DkxFEgGr
4/yai9XYrzh8bypirE7ig6DWKJXTyDqvEOQ0v7w/lO2N6FVYwHAR7YL4SZ8+g57Qo4cTprOq4x6/
x3NHsP/lc/b/tejG0T9qXd6oH3rRXr20N446GlzB6W2ldbzsJKI4kmk+k+LmrVKBHJw5cPRf9E0c
ow6JPANZyygu8N8hcCEjG4AX+bHsCyjqavBKUjZy5ofG0hK3SCa2PoOmJLI9XNYlO+C9jfXcZQ6Q
sOVdHmoNuHUFd7d41MYG8HNxHM9rdD76+n4+vDL3tCHfCGy0OrSIazIlSsGTX/1YLK7NnWaxMiFw
Nc7h0/iw/DGSPxddo9vY7vhO4z8XRXFOtHCeIIEVbGqrlOY7WCxs7Ibt5YsRoBGsTX4iPg6v+uw3
U1+j80Ivo8bmtKhIrESbfLvDI5QZfbBkmbllIyyBd1Cezq/gd0vuePCYxLp0QoY3d92ByoagpC5m
it3q59Kevd3CPcjKrV2UwGky8R1kYL1htVp845x5wJuJ+Q8sKzehpsSFyNROqKWTqGFy16esVtPF
MQ0fJjw3JLPXYbfKh5a6v18jte/Q9d1BCUkWIyqQMzoscaGvFGUXNT4gN7xuBFhlzQB5eCNb2uoY
oU+XwzaJtsjEKAa7l4K7IRWbrPexFIiUFEAlMmKzPx4P4PuFZjiOgpVPY4dAnxiSrJXzLYOTMFKL
9whiBzVgJ9RTtUuehQqUm4Xl7xBPOK127iZqH0hyPJPejIrZWu1z5FF1ARDg9E/pBgIZqNvSShsC
uRMv4s560X61taJZqp+S5zIqTuuc3fxhBlOUeCS5lnYkFOa4oRpGZv3UJRfr8lTU8OLIgurlQ6O5
U7rKOfaot8vWCVZNLqsZshzyeiKzV0TyzLj727RCh+ubMxgO52/ympkgmzs3vB6TzcC83amwIg7u
k0IVR27+y96m0xiHoFYjklowTRh0IxswZLvu73TMG7EvP+cezMxk//mWbPycVhEGsr7wRKLSfFIh
5sHimLmUxDmBhxPTHFv3SkZ4P6Rgq7/lXjbHlsjiSUo6SlkJX8H6HlyF0ogYUd33Q0R19NYEFyF4
ss7a/6olQbdfz7dFKAXKTADzAtUauXIhdp0yVb8fTCcct6De6EWqDXNEzCEbaJ4zgxLeHOPv8BnL
caS7VUBVr7Zzez3Qi7WVVlN/SprJIUrNSBwhT45kG67x4WX2q7WPAEgpKloaWYUX+bXQpgkk7rZN
PwfKZlNoIblAFx0nvUM4l4L2FczKnvUSPO0z6zakUsZCrC+Rf+Wc/IiV3zhm21J50uM+WUxhVSuW
3LuazA+pNViRWQD1izbaExfiQbbgVE8Yt05oaS6JxwWE0X3pBfdYQD87gBtGJdS9TigATLJYtLJo
W2hvRzQblDnyWV2DLZJhWrYsyN8FU//9FmGG+NBZXGbV7mcWo+IDRP/Mv1piuVG0fm5AttROFv0r
/7VuIBJ7a+jQr7E6nX7D8F4S+0He2oyG4DFwSqiA1rHiEx9VXdoxcpC3XWJQ6mYy+IA36trY2qP2
kT+tE1xRSQdWzsu0VGzOWIgBmTHPzqprty2cB6x0kmbfMkt6CSfJ6TXXCTPpDxMzU+kh4mRI0xBn
NVF+aMs+nwo7YdQgeZHh9LlAHb+O+Ltdg2+WZ610WCcrqZwbb9GTW8/8GYRw4RRdUEazF/SBC2c0
BoFhHjWTRCHlkR/gAcwTSoTHh5ccrN3C5yxNI/tW1kgovot9kL8RgTCRyh4MbpDDItDsQhUBZdf3
I5HIxf+pL8gK7pRFIfQ43dBpB1HDYv37neov823TSwMptpAN2a1A25GVe6mm55vSdTwjp4Cv5it2
sdTe74mD7BVxKy6yEWdApLv45jQ79zF6NTN15lsKvpAqZIHrtukbtskZPfHLhLG7/0X3TNWdFOiz
kx6vGirV8iN2/nkjCtmPcFHGDNx2W55bI4meVqkD2j4OFQsQHV4ULn43pNEikZK3M1x4mq18CMhw
BnNI1xalimRpE5kijBovmqanci+nkerrDaxlEST6hG4jOJx+UXwJMcZ9/QWz/RM4Tkk4m18d3EhM
oso2akpLcKmd7CPzXB7UMwQMfSkSNjFYQgaYttCRk0VI2S/6yU1BxVgOQHkpiI0Y4TaorSuQg960
geVKqzz1wAZ1W/O8DG7rEyg8U5r507waFTtCNe5qrEICerf/smu3aIo7DuxMlrzGxSU2F2CSVUHG
v3TI2+thtHak6iCWNEe9zag5pPnSY/7Eh5NLxKQZHotaRc1y6HOmQopScCnoHaVjvp8JNN4rq+99
e6dLWGvf/SRxnYKfnZfEgeYQ+d+saCCZ1tbseWJdSOTIQA60vbodyRiYmxp74gm+xC8Zvle4c47X
o89h8ZtULAAL4GSeAx8TDdkmcXgyZWOQd+7uQ8L1Ijv5NQPJmkFfQCKThUtQWh79BJ5xl+hB95cF
XDKFSpuKxMxFXbKZaspckIBKzzN1g72j5OSf0fyrtpvIruOw+ItLGGid2AUshkf0zjOnkdov6jHU
d97twoOf3j2yNhJUbuA/nfugEcMym5OTqCWksJT4D5SIvELtfzPj1Q2H42T480+YL9GQjoRIZIBB
y+wQ/9KLJQEdSm5m+RWRN3cCoyW+Yuplb+HvqiX+wVfCeY38MhT9ppYzZ+PfUyuhFUpvBYo3566S
PupbedTFwsYkZEpZ0jQvhdsse4SRxnYBXh3dZU4XcguFawxavhxfSZFT/WxRATyr67iMYo1GHFiK
5k8ywjBTtzTVXs/GnQwRVAafywCGdUaTP7DHR1IVkHqErH/jTbGBy6W7sCkZqinMMxQZ/8d0rVpR
mX8pbAJQbpgwP6g2d8sobjJRYVMMSPMLRG4lfwpphWAYFYCWQzOjIqWkswSzDVF9SeSr5JEa95V2
IOgQ9dxP2MIcNRTZmUQiClOGPHSUhIPCs9QjxJtTKvMoABNgvBornlpbwLQZKO1tCR2vnJwOTJxX
TY+VtXqVl2IgZdx98rzxJJl+WpLKFPhCmIidzxXTdfcgFCQYU2vFR1K0YS8SlIg5kAIQl6j3Syq2
6mkfjHjOWJdQiGznRP3vUYsFsZKdQLcGnhgjYM6r5Fnu/IXT4SYTT2zb9IXAdTlVB338dOsspLUh
CQcPL6MeqOqrfeu+36tsRYRsnrSOddRODoXNH1r5P3n1crqsxc59o8obN8jOE6xVwfP23J9bLJA1
7gTcqoz32CCsi7qbxJfKoejEF1Xz+CuU+4gZ/3NzmcfhkFdGsYBdUgxx/qkMMVYo0QVXEa//btvZ
+L2bEevG14BLzeZjB7hUOkro572PnyJGP/GQcIj7PYIgK6va/sJZfihN53rBiYuRGUKTFJZ99e2L
ufg756CPZAhKWc9QwcpF59AT6oUPnb3iyeKyEzlrDiye1FkeV97s3sbtL0e2uWDCI4iQduq5hMhK
zj2Y8C552pbYsPyCI1L3gPxliJe/K5DKauvtys+9Ioxa2ZEpq6hNW334//PcS51nXg9oph/zOB1K
LaBShcKHxznTjEc8kQAtlZBwYPRNBDgUFkDvL9PP0X8R4tlUP3LoHj9Yv35b96nzupVVdz20yOiM
Yd9BSoyW2d57fWMFCBjJZ8HeJ5iQggE8YDwtwf9aa5u83iyK0GX8cqdr3emLK+0qQ71KW532VBAM
2zUUUMaxoh1SfAQdZ4kf/SEHNU52Y3DAYBi1NOpfsdC5qVGMn4bXw//Sn30NMoKuRdcDiZYUz4Al
hQjj55TX7XRHhtOHUDlXoHJDT6hBHL9DE1+7ez/k8DhP+33MaYjqPVZJvCRetPRQ9T5JdkgM11ax
UB6Yv4HQUEilXeA/0HdaiVVj09xx8XVWVBYXuqF+wKW/lMO1JlPEE4+S7O0Z6UVb6FG09nBzA+bc
rMPTYDTKd+YBUROyj4Aa0uqu2Ct7DBBoIpcNH8Dud+bMP0JrnPTY58fNVpb9Vvfzvg8TpuWNIP86
osqQ53fZRo704bs/8+eWGUbg0RMKMl0vW3pKFrfrUID4k8S4HTIUVRzOfXn0/Ei4WZuH62P+RRhP
Wh9RAHgchhXptYshtxsmxtW34jvifHld1WhnqR4jj/AJ9QWZGErJF3T27KephWRdvQooM9uwd8rm
ztLWvCuAl6bs3gv+qGZ292s8CVmXmdaTPSedSK9X30rZkgBKblAe5pxndFYEzNG5h2pGwOlSvGiL
E8RkndGpHw2IwL06clair1qer1wKFnudVYXsCm41r1d5XOoJhpDobJLh8orXHipCKbAAeC2Ayrq+
Ukv5PMSbJcpJG4s4qGS4hUldhRobpN8CVUIwsZRgExuP7+daX1mzvXF8jmf01O/JpVqid9zda8NW
F5ufg5EtIXluk8ADIxeHj572rhC/ncUO9/9C8La1GX9Z8Pd6ubM1t/0hiM6n29e0W5k7orGTUXf0
YoX7jpRRks6oyeRzwb31XcPbut1+1Qy3++CNKL0cVlMivertvaVfWcziLAnCpgz0Pji6fBg56DD4
qKuQOnxAq4LWqhSAUxpecaaIA+kmVWPkwokPy4/NeHBuDir9h408ddefERsLLmXFSs1v4hww2i0t
0DXrrASHR5bpd/pJXxDzjgK0A6xTtn5rpO76pURlSBButmQVYj6HSg/w1kO70NKDtFrBoWdjgxwp
sXxr4JT8csLs21mE0wf93vH/zEP0b7jU69lK8xLYfYm0ZDATPkHitiPZw8PWKfW+jYRmpPSYTtg0
gxhlwcMjVsZ+3sG8iQfxPuRMw0zlsp5hBmNbIyDw2RsJsUMFwgISZ3eqBXS4RzzdAyaHFpPVc6eu
eoPX0XNBfirCmHyJbSL2QcTHmUnqPSFbUQ+C7wHU+WLqRyP4Ui2rZEiB47jMiVrj0vQw5pdERDZ9
lbxr41ryggU1dSNMxmG/rIPSCoM1DdDlILD6aTPIvn6Q0ELylA9nIFpHfzeHZIymPLdpNeso0LKp
Jk8m+6hoUNFvWeYHg1e4cRkBQED4/qru6rdoC0JxTGkcGnNwzhGC0GMFz+zRBX0Lz5BLJQypthcV
vbZUPy1bbak8Eka8ihC4SFd1+QWRVQ4ejBywjRaCSiytYYNjYovYpyqK4GSp80nyQ55W4QnrzZAQ
g64D4WK0YAF3Bu7e4glkzZNDkGuHlCJBSqWHWZgQeLMTYcJqkgQ32HTHX4TO/iaFCqkuPwI//HT7
WFL93UFhdZ/OU+pZtRmR28ADaNVEK1lRCLg5WXQgwlQydxoEWiEsOqwO7UqC7mksHDh8KOx1yTUs
OlQSPzw4OtO6n+U5wit/oeaJ3QiVNxdrFXAUeNzNz61+VFgs23ugiQ76KDl/w8tXkDUoxcDlXD3o
5kflBt+4H5AovPOBsDT+J0TveunxyYgDzdOyh2JI+6mruzxtFTaT5ap0+Y4erQy4fHyF2LNxbUmt
AgsTetaxprS785WK1IQwlmfLaJq9pXy9ctJGQ4XZGEs6kVpujOe1mycAVORyup1T0H1A+HcqsHoM
gibJjKMqLM8dcLfqUlA4xo8kTqEf5jv+fx6bnSl4PNhosvici8KxpQeuUhtSnUMIV9x7V3/hV9HC
NuNEItC3FOHvN5f18VDI+4lIInQW/v+LrJ/Cqmsz9eeh5z2GPGAXqzHZzNvxuofINhuk5JChnOVH
Gk3xTzrnOn3CmvzT6X5CEgj/fK5gj6IYu1zPwv/ABMvO0Fd42k9uAq47QF67X0mAZMFQaz4bAo4G
2fMF+9mmWZB3h39WTzGv915Wkz+W00rixdJ/FXcr0I6azS+nllPOSgW3CWIwRsTck5FZpUU8zmnv
F8R4NK7LVf2dPPZOp7sCG4trCTVo/nRbzFEVC48q+gud3QuVNl/2PE4HCYPCjit8dLAJbfSCP/XD
q6HLmdoklQ9zsXF2YVZq0hUVbYrPzYnBVWxuMC+qmzFaCFT/+qb00Hobb7FhD4xfpp+ofPqBztoh
gKQp+IGZmWTkSrL8G1/JVT6h+S977dFFe1mMKmutLKL8+j0xb3I51Ret/owg3Rk7+BRxoVKQzdG6
ztH2hePy/K0NQ4zeICxkgUB+/Bt3ExzrNX0fI4TFLJ4OzdgXYkUwTDnTYSxXJfLtPcOzHLRR1w78
jYHAY/BjwSD6sYjd7Hize5UXOPfdnAsCV1YoZt9iACQxwSnGFIUEzVcGhQwGvfSSUsegazhBozne
YSbmU+XRqFLNfCTWe2hjAW9+SPOpqILchyAJPbUKK9S5C7ZtsfvO0057xrSKZsY5Gsi6kUYAjBXZ
DVr77Ys0pU8y/wqsOaj3tyyXZunVX/nDON9WeMyMQSbDu/qPrzcgguSQyF/WfvNeSEbC2vGnSNk3
CXgYdG5SGv110Uq4NSAekbPuFDfNAwjhG9evCVJLnmT1/tsagZ9UIK8FdUXDxAvmXOJKGKromrX4
zno1i6Ry+UusDdz4kKUmY+ajVdZRrHuQ++ZjqP7vCmEnYYgrAw8QaeVp7wJonLHYqPcflX2oq5CF
M7JZUncLq4QS9wb3M0kncX1+JLHJzbCnvhBIE7QdjBNFbzYW/OlIMMo7la990VeYFTkjRcyoLvK6
6f8EnBa1lUkUyCWDBK2H+T3583PuNa/Iol/NWWnfJINHF6MldLC3KAqjn/1+hU5jjJQ7ENOd3DRa
SPT+bfkZC08CxKOiPqTkox90AX58Or3wGXqzLLLFlKFlsLGTLpboh2WWgHEr0pSG/XsPiJTamzTj
PlEhrtZFLS4YcrC+9tKY9LTtvvZO3D3pHDYkl6z8xe+VMcCtybLMbFHdh5H8Q0mDExPbDN0BQFgY
EbueCW8+nMaQSU7d/RLUG9/HcPqD25prGSNhKKnoe39fXag4iVxnUygZjDU9hU7eJKdrt37eCbNH
GvMR509sS0pZWRPfFDwMLHKD14j7nwsQELIZz/FY96NQopPYD8v/dIM8Q8PrgL3AVpz7GA9hayrl
EtdfVhAXIoeQDFXxDKgNLgRuTzyEUOXFzT/9UN1/tk6blwfiqWegx5UpM6qRq6dM47vDGMvrT60w
Sx/RK5lNoJKMEP4adsnG513idiI7Mdywnem5V/2dBjgTveVUHitRDOHJPZee0pjrqZZvq5bfpt8P
8NYqcJj62+T9/7pYn4fqGw23fiTW+BGuhN7rwofuLh2R2x5KwJWVs20GyNIfet76uz5wHwajNsS1
q/8CFGlH1EpuuSxVW8BvQMxL0KMx3uK9i341NCexjWRz2bfoaKsVjsBx1dD0qojev3OOXUr3uGva
OvdKzwz7mkG0uIYqyU4LFXc6TZsCakYqiZHQCYiTDXiGMO/jYljImuXiAPKWVUjSmbJFcaCCmRyi
F+y5Q7hDRRmIbP4tcQAZtHeaIaT9ALo7d826zuuIUDN/mh03EYGxLooAyUaPdo6Vqimu1byHtGd4
sOu1MmIzVrzOT4rRWdeOvucFMBgwsUykS0kFY7QJQzDp+HXoae8YmNZ7qiEeVC/ZSKSyIMt0aYqX
tNcD2rCiffYn46LRHtx/DlqmpuviKFuZBj6vvKDrutpbldh4RHWTbQH/F5oe3rkC8uRaaG2lbNfs
xFAS/kZKZlfZVNBw5ygqVJEmatDz5QIXbiwVAt48TveZcmgnlS1FuIMk+muGYl47pstCPpt4VX99
tXxAYHHtdf4Uu+N5GYw8rC37CSpMSIqe++kjFGdppXLxwnXRXUi6aLcPKIlUo4AmPHJ4Ns2IQAdX
WZWrpL4iVKYiHJj461evELak/ykDsmmIGu0Kz6XYJP2dRhTgJbKFYUXEMzb6JohZVToG0lsFoF0B
LerHDJIL/Q04VZrdXlzL9r+Aznx6U9f8IHddEJMXcJ0eqW71tUBzaxf0FhuoXqtKby+a/EdLS4Zg
L1S+fqkOSQ/m3Tm7G/7sQA1EL7mAi028ltlC4fdlAXabu6L2oMjdtMLe5QlbVwjuxlrg20afFo+C
/xnT4UTFb1HDC3s1V3+T2tFc5p/xx4Y2GXZMm/hp8wWp1jUdfJS1mWRIY5iviDtz/72YzUQiN0d2
Jl0bdReMmXR5JLUSZnEOxD1y0bal49LTnnjePQEG3wOju0xuqE2PAtovI8ah/DWKTGxFSDPn2VdO
zBnxiuqwwxkYD87Woa0p4RLjyFU1dYcGwKxO4civFPXZNsunrHS0/ANP1aBwIvBnD83BfkNigHj1
/gFjLRaO0H6OevFtlR95Wa1kWqP6jejI1G6A8zeOdSNUUMoAJHy/b8AE3qCRsVL4OXa53PRlpWio
O4jttxx5q8Loc5Rpn2iVG0wSq1/JTss9Gap++rJTRN/0U7DGFFAzBo+bTRvIIW/MqabLUZ/7nGaX
oPjBhLA9JtuB1ER47Xozo9qiEQSfSVfE0oenEfIh+6mV2DCkagURkq+F3YT3yr+249en1k2vOKxe
FvDYpU/eIaHwIfOgC3AK+TN4ifiqQDwz5CWETMofp3G3VStyVNsw+hk9ntk6CE/voP26+50F6cys
y+pUTQ7B9guCCTzC1ZrhRYMeV2RX6EOTDjGvx8OL9memXxeMk3IUdcgZuuIXSQAgvSBlUbN7ErYj
sV+F39O7cTG7ebToNABS/UmbhAFkab2jKZLcVhCnXY2W/7n1omYjonyQmnyEL0YECxAqIzAvJDAf
jLOBfPh3G0U2/srEC2O7NYZgsVfcsfeYEtWcUq7vorsEAnGYKfJ43KMtLHzPOPFmpJvNdQIYa4Ci
0dELLhFuveHgjOBfE4iyz3SzltmOlGeQ/a6Ay4dc+5lzdQ1uSdAYXvUwxA99U8LPMFRDQFmdPqA5
mC93r9hMXogth+ieF7Zz541g6D9ecpI/dO7v0Edw5dLfr+NAFApaEsqyibxM7R5aHnEgugHEBFKJ
7N8seZ3KG4XpCvPWcS0Z5khmBpblXTRMED5U+ohX/8orezFnCLuaz/L0r5COvgA2YSrRDW74UorQ
Seot9izjyTHuLLZqh+tO2C5iij56woweykva/U0040U0Up0s4OxXZRre+cluv8rUzORQmVGgDG6x
2RfyY5gXOdee1jAl10vkwX6OWDP959HXjKGck8B51xxRMsrzZWxn1syU7tjpacOd74WwkQ7G3EsQ
GeC6D9DTGgdhQIzjbMXDVHESmSYPpITpc/KRrgVHVJRI+eVYwTpqtpiEOt7loL1rPcH+wh8cz76f
R1H7H/NqCi7/TnGwAllYQr6u4nG9ANVlUVTRrW2FJs1n+yOxlLHgV2QmFc9n0hyQnoEh9XQ3reci
+7ZoCz5AarHdOi7QOCUlUYa8bVPe4Z4sBw488e/FphJSrKijfz9kjJegw5Nb7V/gaEu8xF6mYxKS
8gyP/c+0sNfzXl/OWmGrMd2cBw1ovsqZl/WBtgXZ7uw0Rx9QL1fxcgXha0Lpe04RMpoHF+eAaSQ4
u1yjGkfXZ5IX/JF2fDIa0N7gUAX4aauxpdKuUqyeRFHAjr8mGaaDmxbaaJCSr566RABDzhslDrMO
ePmMH/Wn1Uft7XNgO6E4pmZQpAXYtjRSyVpxg+y0riy+5AJ4Bh/y0mzDewKrw6Ir931baMi12WiX
+R/SiiKgmoI6SkjHOcCg5A6n/UmN5ai6abT87xFgzDccUkYelNucORfTq1HujoHH/dB8IZnsJcbC
X0RJ6QLMarFgy8BFSFnsSQtIJKTaqyh6sHM6n3pq5URmDjthX0oTyEIVFXkHEHg/1om8dtMa0/yc
ErIQdd25UeXjD9fNazzNdufRHdkGUOBiiWa9lAtjTchwoxO6Le2MX06xM5xlkO+iL4J6kI2k330V
sR+BCjPuUqkobnPlsAe2EzMIc2BJOik5LGPLBcDyWCvWVnM7eSsKXzfbzsS4ZJQB9zLekKQvIkDW
kFMXWNw6e4/KEPVG97HEkqjsK8PPQokhNzselBntH8M9bJ1avRBqBYun1SVUjs/v8vJgxG7BvO9X
Or942qL+eyjJGoGl485hg/DEVskrJAkLzgU85bU45AgN+4W3um2EwbFtATnjlxGvOy/wAgQuLNpt
uif3imXwh1iW/4XMX37vH4a79voxx8RRiwi2ZMsLTU9qfDzBdAA9HqDJloLwIl55gxJaSYiPZFHh
IQ7uyhGSyuzdOcfzgbc6k3gYUONDunNdoxOhUDpDgKXExecbTsBzw32nVOalHV3CG2uv7L6HNEgf
zexz3oU8ROyzvB5kN4x41KZJHLW/JEtscE3lO6zlACoSGggGNXxvvY66ckIpdQrZxsd/Mvs+Pbu+
xf7SP6JcSV+3IXXV4aVFcWCV8WKaGdyMrak0Kz/eGsNa4H3BZy9Q4xx/HB37Gq1G2BuX/P+TcNa3
f6N3lPE8hQl0qFLYBmxBaWa7YUSaAvaRFDaApwBay+4z1Q9ORme+AsNPGL0T+1csqlRAhip7Bltd
HLyUCLbLt5QaRlvvCHvcd3muq/o5bIgACjFB8H8D6iZEY2gVCOh5/fGZ1hEVq7MxI87Bd2FR9FMP
QOkzi/fPGi9R81ooUYdv8vY06kxBLgRFAsqnGBFvBU5mzsjokYsBTboH4euFLV7w7x78TuxhYmBs
reTkZSh4CI/b0f9Zdmus8Xzk9mDHOt3UvCJitBif0FpLoHlLFsBdoW8+ItYeh4/QNS8yL8/mD6HQ
QzCYFLNIZMRKbL0BXp7pTf/CPsH12VoOusIyEbrnXWaAFZBD/o2pjztgMFIlLqrnY2agrklzLHQP
iAyDoPHThGBrA9t6GhBc3kf5m3VxgTBgFpVLbdDaokkLzZVukaJJDFw14YH7RclezXOUr6xBKs1n
MpskqZyCbp2gJIa4xEBaZ7xnN8QIc9WfxDkbUFjOOAAXflK/EGCQkv3mVS94tC0yA6OmDHyAarom
ZQbpLEKYszTTRmYkfVYwQHgm9G96qz754DCYQyvHZ1dIUZu4xIXNKp3xySOJ9uual/R83Mk78b/M
wel2tyYxGHoJtzVsjzAYpTng2HXNHH7CbBoOWvHwahKbk4gXVzCIT/dh0sgb+M7xl9rYnKaQDKKn
rNqHDpzg9/AMTisaMASPo1g2DraVHOVHw6AOaBd2PgVPeRZHsGHoB170YN0M2xSKosFmpP0SMUtg
YAHwtAR9nD/myNTXNQPbo7kBQdyFlJ0+MSYX372MUKvdbU3HcG2DTFUIHW3oVXJFmZq+LKY5D2hy
TI5k94n4tFrOZshb701xCSwEIa2P2KsA+C0v0qB2kKNYLrhgdQ85wFmuApTN4MkuofwQMTbfLQlg
f4lLNDr/RY+fMY4IK7n68O+TG41Dd1MfDgO9BJjsOsUR1dfvXpHcOExb4lkR6Tsmh/0nU4EINDnF
uHPOLWEY7HnEGovkRkrZd6bkrnNUXuLH4P5Q8Pdo2iQe5s3XGJQl5c9+GEmMAelZlWB9o3Tb+NnI
qs8ymLqPG/Q61So6h6sCkRobt0KwfqJ+tq2d4WUVKyTucuHteDqcWKJ9rGlMwYgWDir0HtICI/1O
Mejb9iRCBqCC/2soPil6xuHNva/sm86lexb13PvBufxiGq+V7UQ3Q5S9np/wcDdAdR+6fXOZgEgB
EMAdSUnKQP3MapYLVkA5ZS7hyDZ3HmWZGifiMHUZjx6WfhgYupC+Vw8pswX+4n5r9s8rWghEAsNy
hnyYKe25FvVQFzHnLoJHCCA8NwFRrIBsdOKMeWK6/xdBhiUkI5/XmWp2WaYmMYNSEhGAbkSkLNoF
2ix3BAbcM/IorAzQpKglraGMZbkiX5c6qDiXHk+hAX4bjgCOCcZFCQuUVUlrvqeZvdwU7RETQQSv
wHSH4nS9CrPnklUSWnnm1gUCPgHkL6dQbBe7lK2XML0DHMLQ55sXBahqLGZiuuXJKTw33U7C/YlY
C5GhvNl+sKTmaWBWAtTRT2dEzztZ2TxQ/KvpH1oeARJE2wPfJVmkXGxyrEfMpC0JulDNhDKtZ6xl
eJH+LgQAhE0ElZvxqpbQCXtVcdtCDx4DvJghT+GaQzq2Qb12W54DraQYljf2AIMsU9b+YioToX30
tFD1aZgFLt+GWD+aM5WDdzkcWntVAlPDyBZLP0lHFc9TBbx2u4Q9pd47aJap+FMdKqEF3zTxeI+9
3VS4KnHlO/1Cq7SecJrr7wireUQkBCE/3Y4H8u+iLxSILYACpRbJNjprzbYoFmLZ2TIQQtHhpsQg
5R5HK6agTTn4ZGjjj0hob+t9YEO6KsofGtHK5buCRfHPcYLOq9BSuta+SkxDaVlRNltFvBU+c3Jt
ZSdsGFVwKJ+eIBkp6oQOLqJ99Npk4mGPHJlfGfOBE7d9+0/P24k4JNHL+SV/cKgDKOV/CbbIcpeK
yMtoQGSRdlgB9Wx/FS6OJfpk04I3cj9dnlycCe9LI9RWIhhhokGn6HKti+odCyT50r9hmMKoixrP
5JUvtPcjA/UKS/kDGfMZOxEfwweSBXgBz8tG/g7ivHwaXHg4Pq4KP9zl1Mt7O1ijIpg/mo6V7YQ2
URcEwmjBKMp3yC1dubiLX1qXhE8b4gxvfYTXO2yAh+ZsumySXPKpwO3GX9pi78uu1TmGIO07Jwhs
IKOz/cB/fOKS/b9zpTGEVZn6mRsnU7tMc/tFgnQIzR8mVKseleWfQgPpI9BGtGjMi00oOrc0syCq
Ihe8lSVPURM2OnNGM4r6ehmxFdDMtcuF9Cd2DXG39bXOHQ1ddv1SsKL64txOJo9baWvw++KqWGK9
LVhoMY2Bu8U5MJ4yQEMnQp0bYWjCq0U/2LPW+iKmM83AsB17jogNeh0wdLCy3Pv1ZERYmDKAQVhs
6UqOXFZNm4XJWSJRb/liFvJgCJZgP9XD6kgErYTi7f9v04g3Y1YbIIziNmAuEKJqOegSFc6KeRsb
uG5VbNVWMdpUfOF2Dzb/9D6OvQ3i5Orqju0rk7neZ1MmVJULyYROT4AY5wSE16wYhpdKevi9UIq8
+tLojKQuvX+axZy47dHyRU1QXSHeNL3qc/2iaPhLVJ7u7vb76G4cJWZLdhHQ1dReITJGkpSiUBr5
jVhMOJ8tnT6qQvuxKYynKK1+zAV08QU76t6h4vJ9fMgHHqCGD7zwLqPUwjZ3AVOOws3gKJb4kp3b
B9fKGgP09jRL22B2aVoR80cCMByA3dUhCBGjOx849+tnzW5IezWzUqqZALhucYiuPW6OnJyiksVe
ir5O1szJY2zFa08t/yNXpeA6qTsSCFfW+XHRC5tIs9SMowqxVs7D1tYRR946HU0+uTX40TD7vIIT
KZlN+y23goWbGWGGQPQheYqXdNyZGAbQHqy/DGP1nyl8qo7tB1pXkKsGZDukes2Tv+lo04vCvoCY
r/Xw7m3dUUEXt3BCki1GdYTDls3lIMZH7zyYdFsebXt/xwSK/bJUdYyIXOGHyhO3/A2s2omJa31Q
q2M6jvjrJxDC6p6MPdoJdRsLklrOje8hUXteox3zH8dZjpHsVcN+fGl2ahrqYHFwsGhdSnL0hP2a
82Hy/UKHvzsjb2QEag8rynMTS28GXwF0C31DyyRcmRGRYTWwyWZcTxpsGyyZVurQQsyPnUY9MXMr
1o6rPv/R/PCNtpv6GNNpTUeeDGBI7zS0rJTOR6BIT95di4VoAFJ35pfG2JKnBneu+uYol3E1M0LX
9b5ObwHdbVT2NOnJvMSM5IVu1TYTNBAoaRwTXYuRLbnhg5kekPQMsIloow1QSsaCJpWjRUNXimVm
s+68Thex4guNTuF4NKF7PwpLodPEOR27lBsJraIhFKW9ILNM05CrJSQF29AM8IdDnoi1Dz4jFYX0
Dg2xmIdHqi3ZCdkCod6mFhBsbM2SY2YB1apmf1raCoPsuIiNNOBsD46FlCLwAmT0GlXFXTE5J/Qm
niDlvmfgctjgjizjVqCxsIjn/Ndr9J6log4dX4UVNN4Y/YpVerf0qKco6/sOnn6Yuq8c5LIrScW+
MqXAXZ6DhVca9X+9PufBYkapHGyHoIm8nzPyNAdS4Zy17tBMR0ZrbvpClGqyPmM5lllnxNnC9SCp
8jaQq6onMYAUK786c/1ut6uyu2rhDj6/1hJQqxGYeYI/bX1yVLopBB08aOfGUKj+HhoaYQhvjpQR
xrgIczM7L8Byb3skHsMqk0o59OSLh9rHgPuORnGXCXr6LywCnp92/MCHDUqTox3ehbRbK677CgTS
TfYiyFnmGjFVfkHBfnFrdTUvojgwiIIlLEuLNkeHPvvWdJ69o0J3co6P6XG1SzpnvnhJjc35bN8w
yK2L8DDZEe5IlnABPwg8IPLiWV63Y9Ptg0g8YToDnczpc8f6d0/412xUroMTCgRRYMMQ+MyXiclj
SLdoCYABpU+EFKCkAn2e4X0r3OKt5Ul59bcmLiX/EWTLpcF0Z5vu6XDVGjtU0sZ2Db0F/zcSb88L
29cKnvg21JHLPgcOav1z/zU7p7Uic+o3aB3bX7QGOCcXMrZ9KD2lk20MQRaVVTEbIj+dXPd85t7H
3uYh9rNoDD/Q+xAfAhyDd0qjlMUbniZP/BP925Oi5+0EgY1eGtzjeof/lqdNy6lNSzpEC9t7yeOW
x9PFRIoi3leHUh/VXx5paOT50J1v1/25Lu8sPb7MC968CXAlra66+B35ledyBIkzf0FhcxTazz96
sqOgcQMrLXgGYo//07PEZvWCaY0a/lBGyDG1J+rp5e8nA67GvWCpZRsQfopSbUc3bjsSCOPR5vxp
f2UB30cfeSjdO+xpjWsFtaHf1u/LJjr1elWuCjiTpVb/EY6hEEh2ATAuVvL+S2ly5tZiiS5eyHoV
TpGeOpJOYVbbddFBkAHhp7mSbj8EZAWKfX8Dc542Ty32fo7ejjxUQ753f4Ht8rveu2FbfFvgnC+s
Pk71z7R9EJKXn+QTyIGGwW8gXVgyjwoSeyFmyswET0GMOQoxcnjQyNdP9v77KjQ9HibnhhoxYs1f
EXOCQMrdLCzAxFkac4KHNUa8zNGRZ+bUNu+8FnJaUIOt/YdjCetUj/UcGODE2IKg4P2rUP10UoWQ
WKdeK1gAkrcke1JITktQvBT+58ISjwSZ7Y1A9ZFwYWgG8rXHEU4P+esPVwtSKnt3l/BI0n+JS58k
6TxEJwxjHWDIj5XaQFLHpfW7sloWnLpSBio4MUrZbqlobJsQtzRo9xDwP2bIUye1UgUrgc41VCq1
SF4vxliPDkc+uH64MkMvoTuN8DSYTkljQtKYKY3Pq+xjP44zW3wKV4wBHicQg7O4pQd5U5IdOqu/
NqrOAH9dyA3s9XGLffuH8HxuM+Tuj+/1ZURMm4TA9eBe26k/Jaohwjox5OIx0LTbQgD1tE9jDlE/
aEUoJgD+PnZPfHWtTeU26hwY5kdcgwP4Ho24y+OXOCKlK9H8JUgDl+2VJjePQ8MVoQ1I09QwUhDQ
/SqEgy/DF57Y2+KM3bi2jD65w/4Y4sVT/I/Jw06NLpHbl0toeljZtkyLW9kRjToRwDsf6KkZBH+o
VySpWMn1EJ9peE+bfAcxCDGiqSFEISsLUQbOjUGUcDPUD5wmREwY/ebwKdUdqD3JtYcuTHfOVNJo
Fr2yDsI5FPXg3iI+2YNOkWos3+rt09ckBgbjHiRp1AbtCO3HQCwH39ke9xoajmJIfd8MbUyoDaYL
SayWmx4Tw5p0FMCKiKloBTkG/bEG8q9qneTZe22f4GiJzQhKqy8UOlS0eiCENdyto4vI7SgCtLmO
92FKtcsI81ZbgbFZiAJhMnO69lC2VfVnHWcAUSiANzcyth7i4QS8ouSkUw55dTlg1R362H2ICPAN
irvoc2/5ffOlvvt9QaPlFjyObFwVeY4CmA4roh8aOAzQ16udFb+jpaDZ01uo8V5Lz/mjBX9EKNGg
5l7BX/3Fbx26BTMD3gpK2CrCE5+hftOpjszZvVq24vsiKiNBk8EC1R9M7Y1PHU3WSztEAlrwU7R+
sRadS8fhbFv2FTzFtrzCKOaaDRUos7INphsV0zHRLXspNJ675jhrHSG5wBuljSOrIsJN1ByLlmdo
Xx4YPHx7OB5gFdndlHhRQUzyajB61UMUjVLYJv+3CuJ9e/aqFCJKhDMb5qN39M/EvWuFI2/7D61h
HvVWXgmeZJGyTMIerjzmSe7uKh+afUD/CQoEuDKudkwkVm6wjsXQjfgC3A+Od4QhbjedIS0KttMa
iiFrarttthzXD++UcfHadejcu2rvtkYfVAWX9tYE9FMglZ2z4037LAkv6ZQw4d8s3xqm2ujH4ZVJ
GAnZvjE/EhI/iWsLPb9RS+FvHclZNLv/WLBhDgsqqDEBUhZSliF0a4A3xBlRgwRJJOdF33f9Np/X
xoTHJiLqxPMjhlcPmnfl+IAKxKEhZuL9MqGWQyxQl6A88NWwJgUIS+d9Nd0ioxRRDKD9T3xvBxB7
OgHJRf+lOTaw86RkIXYTofXrbkvij/LxjeovP8nDxZexOl1QV+rX+/IY30STx21k1GvloLrlNoRV
oBRdNYd7EwenR1KGuPX5A2Trc2sEJ+N6cZSSlL9fmNio3WyLZuEgrn3N78+LuI+9dc2/eec23HhH
HLwLFusfS3rvSgAUsV/ZTgDwLWm5Vj2h5dw9qPdHgHv5JqYe7lljxJ31751l+svD+SMiKFAd9EFw
fCv8M1PxWnoixPOHEEsuFqcl6LURLoc87a2CkAClS/uqpb9cJajP2rtXq0aSvgkNsGL1mymKvpIH
U6fP7fD0TcnevzhNvBqBnXBTqU5KgoienLs3pY9gm3uqwCOd5gv2IIEyL1zIxi3dEtXly2jWlZUU
PhaXYWnl5ze1UVfvDz37Zkv+x7ts9eyFYsK2LpTGSMWmazfjHfImR5ji0/lU6v6xTN6CRUkXgsAL
lqVywrXSCxk/a9vH97soqSsE3zLyTa6/y0ift4Zo6YDBytK9jxzrFensllFZu8FpHv5BVvpK8KUP
x7cyXSULnl1wJWqlqdzQsO5UCV4YbxALbVRVO9ZNuIsAI9usGole/fcTOEnEGFS8/+qwlCNdXzBS
mE9mLLP5fdqxI6+WRH09QRdgkZpiNmxIKOC+132SiTFZXotDZgwS6feohvbOtsRAtbKKzlBnIewO
LF0nb2oz9LlMJjDaCy1cxUwu11CUAfSxSq9HkUpG+xAIc2iu65Sk3CZrkrCSyP8QPjVN70rg206J
6eQcT9keeF3RK+yHU7RoYuzap8p6SFcxuoRBZ5iNgnqnK1arvWZi3hNRX/RfX1uBOYnnyyVLHFYi
QLYHIu1j8n+UL2VLQnRKD/BNZSW++dn54e4XXLhU5YaYfTpY8ukPxZMrzxtflYbMkoaqEz+hir0h
eTrvgHe5zN6o/Qr4BwSZc+VB9ltaEA+l0HBN+3u/2bXDk3LVI6arbiydWfSkbr9WGn/Nt45yze1X
8wGQQzWTfEJ0XZ+c4YQX9fGi6KdotTL97pErnu7+rQEaZyLK5MdiyDXvAMO/gwogWpnToMbfb2l1
nn9ataHlzMDzACCmqYCjNc5m1JY7CwmnvJjTvLRHDL+I+dCmaRyv1Ai88ShNWfgYlckGhO/gu3p0
1MTdyitKJ9KtkmtyU3zaxtV9kTkwmvMmF3QlnziLsv8tCqRieTbKW9y/tdoRviRcicQ8PQGpKgKW
qqbvrCNdDuvk6ThLr91g4pkRbhlNOsZF6c035nphS0gWondmT9NoO9ImtES/DXPgQS1c+2Aok4Rn
gvN/ePWiV6wUekX2B0St6HikbzYhditvIe8z7MkTABZ3yfnnbcPFtnQzUnYAs72qqzRmyKbVrc19
A7E1GD4fQ0PWNthzZI2H+9iY9LMEOjEhKpJoycOT4LnN3btUw5tLqdchr+WV37VBQ6Sox7Ew+YDd
BbsMyJ7aBiDHNNdrbCcrIImZ6RMXOcFHKblvwVPFDM2oETC4OboM+KeLObCa6Agya8t7kqQ9FLyg
Xfgf/UQ6p49G0zlxzUpsO0FTF7bSjTpUFME+Lnvd1SHc5B863YZN2vIOVih4VhB3GRouHJY3F65v
N29eyIp9I4nqLKeFX+ozU3fnt8ied+GexKKuALWRwGzVlQrVrY2NlR//LZ1yxjsIa6RlYDP7tAcH
j8K5kl0g9vTPoKYxoXKCSNW+ZdwU2uyF1RWEZCfxBlM1fUMVPE1MTMuRB9uCNJzH2GKxEaVnJxjm
uFnGcIWytoxJO8hP7J7J/eINnNI9+WU8HIDqyR2/DFQ9rYyHoKLUxQjD8D8d4ORW1+adJ5oKAeEo
XJsCoTJzJbSLK8cH6PBeQ30rrYUs77i0Xdm0GI689y25GzjAApxxsZL39Ptf/L1LWX9MhY0BAJbV
q97qrsNOpPqCZLM1w9qaBsPr1ohICeZzXmwYpVSoHokSrI1tpHbIFNCBJQCoA4b+YwS9VJ6pMRze
DuBlPj+T3o49XfcOqJfCls1UHOnsED4UH+sgyjEQ7F3Cuk8bXTIzLY/HELuV66m+aiTUXzngtrIr
aGgC7B7SqXTONDhhQTMh14YISGebe8tgGAalEZwsQzszEpD5+I11l0IYlt7BhdjqQmHodkMXQGDC
02fR4X3EVF6tnzreZq4fIgpjDONjnnfV6pz7yI7XVBLTJYfTtwFjaTFALA6wbsYU5QKpY5idm50p
THjN8nvNxPqnZuA2tLNli3VFVG9zwFDPZC46McHfJqu1WkjqtittvndXxRp31Y0U8cot0+5gAp8A
gUOVFJ4piFIkvj+UP1ddnki24NvOkSoEekRWCtApzudfGATKsPJrrbVYXo3ppR58Oqknh5Ex6nnO
faqK9CGGESW2x8UK42SLx/vxHEXrEVPOd6zCYR0fcdF+CVAgwvL76PbrWd/5GDiOb3IWB6u6sTBD
TGmq4XdOLIGo5bDPSqS1/aOPI5zu5U9HCfISHfNMpF1WHGytiKN8FsMYqMp39enkysKJO+5+80qX
UVDewijbEc2g1TvZQO/M3ZOxef4Amw3ZDUEDw731bDjAUc2gV9KDDmDdIB4eIuV6iFWAAZmDl/rL
12hxO1iMROCB0P/6u1zvLM63fdVYzxGXD587iKQrpEVfld2YXQ8VfO00Ujx8abDC9mAGd3DNLDO1
ZWsGYkVeNytn3Q5Oh60z5aI3QqYnB/gbzvm43NX8Z0bQj8xwzvw2ppQ0BdnNuGI6DzxN/hw9UGSG
pmKooEuGMQM+HRuMH+X7UxsauTJA3a5008Md+X8bv9o25jv3N01XdeFnGqdlFeNFOwyqkokbpSHy
B0M70uy+Rxwj4VRTYB2Z647DtZAOZcqACAsYR9tiEL5IMHzT8mC1BW4KINe1EuBH6cf15BXHEDCA
8eDuLfaNCFedHWaU3FRZ1YBOHiTUCvFSR7zVMxdigWsmUDxNIk3KYxHZwqx64eGvG6lGciFuWeC3
fXauoe3SUHhWlnVALxz/6utlYlpQyieucKbMBahsRUaEhq1e5oDsJT39ydF6PFHqkZZf9N22/UWQ
li6V83PNmzey4KvLGC6hHIqV6SAvWLQisH2oNtLCnsDjXasdbtaxrJ325Fwd0SAoNeMgSVLH7RHQ
glV6Ms10LVWuMwppjZLBrP8tn6mcQ2cYeFSFe48rfwec3i+g3uKGuveSs/l3WPAqg0qcb47tBQDf
p55CISA0EIjoXlNUGP+8ypmPG3fCWN46Q2S0+2Q8Q2u4ZgNy4eW6qmfsjzFg5NoGDOVLd1VamWZC
Cils+lImoPbvrFW/8aAk+zCORMRyPw9RinoRpO8ixO4LP2pcSUrGv7PrEfLjTlNscBMRD/PauZLG
ngtzDKtiF2EEaUx5Q0/qC8NyUx+h8+yEZLeCeglM4ExIZiCZcPOgXhl3GapHqgdYu8jSBFNx678a
YmrAZ8T4Vb8iYxYFfRj21uXwCDr6Kz918vKmLMXRcgYb3co83G0bGrspc2rZqSDymhirmV0GTyVp
MnCc6GM6P9YhVnkhCzXPESZ98QxEBxlgEfbLstMez4Y/yPqcV2xrExk0rpkjZAmrLENOC9pUIxrx
6qrKftsECna3cOYep3GrIfZyexflzCxxzbagyintC/2j1zDbJecwSJTUqRK92+joPD/qzG7WJLY7
6aZhSxHVn18u0R4msWVb7kOImU/YYMbtZTgfLNjcTyv7X3j1hyDtvoCoVLLiPCwRomLEp85BDa3A
Ko4yjOTRE5hPmaBbfBl1CZyqGhcQofjqRGUAeNoVNnJ7P3jyB5yCV0ab4jmwiP4tYFWzA2LCnqOd
QtBGH80oOG0vD7wI5vumd2NsiR/dhxCHA5VeQEEk3n1WzP2DkUEQ8eU/lFqyGL6/sNoaLZAbjCqD
yVZmPH3Bm3W8oWWxDZ7qHOiRl1mFH3b8xsD8ndXRm+F0XE9EhErCW4bGgy16yPicAkkr/9Z9viEe
UztSfytTTA24Z1EuyzAShMKzh3kspe3f1L4byhMDhlebgpQH45jFfNj6j5dXkzZeKRpAYyY+6IPh
Rc6ec61Y8t04CroueBdX18qIuXazLiXleSJN5v0cCZmYfMnVgZrzVkgGvvs6mzvGNTPv6no/Mgym
XawjU2/FSM1TR4j21ApotDcGCNM64MigwiPBPptHTuOkNpK/yCqQumWwb9/pkBxX98ZJdEwmF0nY
gcZhe2WeNapy4+g950WPCsCmKCOYk9edne0OdO4Gw2X8HYGeC+1sYB1EqB6lIBlqI7/nF93td+ut
/uyeqLe2P/qSAE+s1RUWxwgDrl3goAhL5/B7ilqldMYVQsowqs/rpilI/Cf4iKcsIzVgLZK/LVQE
yOVsHTE0QAeEe/KFzlLs/qPXVPoC6Jy3jH7EHY7awDnoo9WTZSfq5uBCZ0nz2mIJ24tozMiGQrIX
huRJGVe7xpM2KMjHC6Sd8NmjjMEU+14RZTHW+FZdw4VwaqDyZoY725sV4J3xKwocByVuZYG6koFQ
ZUPvZI3NULGU0QtQuOgOrkD2nBbamlychT136HH7oyJE6Qtej3cAOZBBn/aNmqcJx9HrUTNuo5Pq
BhPmUV3cibr0kr7yb35/LC/4lODVWAr6SWT/rI4gI68XC6ShVZdTMm4J8B0/mkDbM2p4r+Ka9sBM
sZSqnRXYTU2+XwoOpZMDxuTB1i71chc5J+aeqMl3lpYcgtjIVD2jkLwoTpF07cK9zB3titldZdAP
n+FMOvGNxUZvr70tHtofLwQVkAK5WwZgZND36AYw1PjxY1UwxaPNE3DeJU4Wb9QjxBYJuD3k3S3H
/FMnuLtJTdPWz0NpRGLRxqx4T/WBxzSRl2qd3FcvWYagSpZIDghD6jssul+sGDcRiGI+osdYWOST
+4UHFwULgmxU0IjEOKeTMSjBmLeYnNz7tNDsH43uiFA4yMnFJSarxFZyKzbcdjojqgowV1KC89p2
ObKtk7B+miS6BoR35C9S16rLPX3ComDRjTpIVRQCMz3gvmdpY4f0YMU9Sr0S8R4akLb5l2XTwjEI
cAESroHTIvOM/IbfLGrBd3T6EZKIHA0dRXcczwX2kw5K1gmsrsvd31UtioDzpl9sr01WiTjzH+pc
0eBq+m2Z9ByGoy4i8VmFl+wMrZhurtSnK9yO6N3Nt9yt4MN5wFrUx6asTPeJI89B1/6tEkw34IBT
ZTNe1rl/kHkPQJkQ+6eESGgPPzpK0JrmjnUvEnQXCKXhEhVsOK+S8PQcgMN3uMqEBuIGrYjiH9pE
8FJEl3rmg57mMQzmn5o/K0U++2SwgIVsptRPIZEbNLPo9GWuW4OftjmNK/6If0xdsQ/5btkVYwiX
pSz57rA/1MuUSDMcXA79S49+YcbyWfjdkHjeWBe9/9/YegpOxSSWdCOk3Pzo0SZybgFVwnrMUB9Q
pk4q1bOlOr8g75EHLCSTnzMzkYOfMbhQXhPyBBIlIgl2lOIzOSE0HU8CYWuHhEM4Fd9VfME8zt2X
DxrOQn4geyisa2E4vaD3797n26wo1h+a41OXEerIyUBkDZFCdTBsYebhKkdKcFQShPdUC38QGl9u
HYGbCumdAs5/oyB7ASl3mQuqsyjo0JzYoYDY2Qfq6mTxolihKXyCt5v0KwSSQg+wiNFvwPAYBoz+
V0lAVykzx4q06ht1cyZ8vIWAwHxYUKuH6A0GkVUMqcwxPV0+mEFc5J/kP9SBYckWRkPfDbGjTD0u
FvwsEkiUjKDQdnwFmI37w5wOy8E6uXyS6Fwr69x1Xeb+r/nwqchU5z/feG/3/58vWtGfGAn08uUl
kI2fRfUTKfGIyT8H8gWDriOTPWG4+ZZBCBBqwr/zXdfV4CBk/Weig4RwcV5JUbKjqlx7RtZUOACw
roht9MRINNReiryaTSHIWNsf9GWRAIu07Rc27O5JHeWLpIMqWAes1HU0AamvPXdaMq+RvOkL+Yrg
7VHf+nhlIX6jWrD5zNqEBbmvjPXPvufevrRxQcGLDLvZx6M3saRmVuzL9tGAeQ87lj6aAuc6uvKa
/1Gm81ZTP2wcVWGmAMIb+SaN9tXX//IFNWlCsLJLYbpCZIcbFet4Dfd79Hgcm90ZhXh3GegM5BEG
xrbacIYJ0cI6LbsEXZmoASouxub772KuD79mA+AtXq/1rPsfma7JvSwsfmtz6MD0vUmQA3LTuPd9
ZrlEUEOQ83wqHWjnjI2mOKF67my6TFD4tM5Q06eu5f88XGFxzPnfJpuBgpKHDkKtjtDVvGewBd+z
ABhiC3GS5k03uvDq4b2EpguR54vwA7x72ssKVfNIZLy3kNq+JkdJphl/yPeZFWOmcANYHr331c2X
y1sK2ydl0UT6vb/lZYPVQJzm4p0pdkRCTH2Hp0NF5ZdrrPnVjHiwZD6Ch4+7YMxyC/0287eh3udx
j2yWwF2yw1hmHgncixlXkZvJUkpG0SVZJOC7cemBya4DJEEIIQ0CmQH+xOJ/c8ZzxpvZo9PUEgOg
cmphOxPK5f49JM1ufMXsyTz+8qv63CEF8BxGFLNmJC49oezhLe0di3udXQRZRwuYa/XTjc4vwY7H
wfUvJPyHIHWq3AsIr9f0RrNQdovPp4ijdW7+R238UfbtQtwuVYsMfB/H7rCth3A27iLI++/IUVrn
PiJgErkOrQ0+T+h6oPyDjBz2eaaCb+BSjDb+uCNIu9aQAFpnRDpNIP7qjKpYY69ZxXj3YMy5LlBO
149O+upL2AY0txdFhX6nHkN+XLAO/QFJTb7C8jGHUkOocpV257PTgw1MCFrfNnQGFUoUQoXL61ky
bzW0xMc7PsRzzT7bLtjHJ53GgQ4sFzMyS1rbxv3D4nrOlCEy+hL0ahNm23uZwFMUt8rxUDb7zu90
PlP0cdff2kyti9IOM5qz3jZ8hghB5u6wSiV3IfdPxymZdOvZBvJrIrkqHPdNBVLBqdH5e80q3/g0
0cIVcRheb+YkRzaBgpyHeyJm1d7w9btHqIT79hoLQaD4k4AL9V+ll+VRKkgMmvoyPoqEacwP1WUK
2jBpyFYnc50+NXAoq+CTkOyXVFrdKNOTK78gHbaLXqT1k+y38IfxgVNEjrocjJgd9A7x+k/mOaGc
R+0JxiaFRrRSbXYhR2NRwhykZQkFA4XvdgrHt6L8IWA19vbR/z0n/IhkIc5x+1hy0nepIsKuXgIq
GTOdIzR1SDolXdNIvIfIeVvNaHOJt7if+DZSl0xkygjja11m9MR5H6pLJOD/qsUP7HlkYthD7SPF
CA37+rib2yQU8OwYU7hwZPMaYSCnMDx1FtWYnGhjBcvs69uBUqELa1dcJNBAK7wm+y/YJThURrPQ
Pe7bnJLwLW8pFg9ueiBraiQcD/1WbbFYn35s02QJX3gxArw50pjXkQFIRW4qD8QgcUXF16VlqvhG
gAOcqaEy5VbI2H7YPLgOTgIQUmU6SEH/UZdYuGYKj/dyPsCRPMxZYHczJrzjtP+aoyGd0nx1Feko
t6fv07KXRfeDldzR8fKcpAGooyJz3/+3JPFXElS5ieHfmo2zeNC+xVkk6TMKbIuxuvrKhbUksq6j
L/fKLAEAlApaL4Pq7kOlgCWYALvRnC7C8CMAz7ZXTrYl8tbG6RRH+ll2K/tIzPH889xO7A05p0Xk
TFbFk7XhRHafgaU6u3SLkkbFGcT1OW5Yze/OT2BU4oLlJYkybjRB0dMdz9EKYBWXYI5PYlhzhJ92
iHWFHH5zNJnewStjLVOHuCm0DG0ZRt7Vk9ljMSB2XGWRnZcH6f/bLV24ordaTjJAWHPbrOgGgbls
v40OIw0aI31OuHQAfX8EB9sE++jZrWyYORIFhos+vj/9f7lM8rtgW2CD93nRk0Swdn/KyWNR4hZb
yFvDJpcfq/W/lIAISg91AWEqRrUhSYDbCWuukhH7JRMbb+m8/VfHkiK99CvSiLO9gn2teihMR50f
uflHBSollark3tgKsqEQhy5qRev2mJ0Av2TXP84mI22A/ZTqugieBPNuFiS8jJDILsxiwIGqXbhW
2aflxVtoZLxm9xtpWReNlXRhRzJvXY0/IaVpje94fhgeOV39Ez6REJlp1AH3/0nzXMMaX8CdHDag
SePOB50Jx1cjCsI65G+Ec+EJXxVJlcP1VBY4i1pIMH1GUUAd/73+jeQLF+f5DcOsSD4q4W6JxUyU
Bhv+PQXefzfeFcuC/BKgjd9fXv2l6sR+1iFwEzN6WJRt+zxECS4+V3Ji4V/gv4xnNUSL6LR4s+dP
KwUZG1uECy8oLEVYyCyoZSJ8tWX4HlYkJ1bVj4outpwbo17BAK/4fS6lkrsW5kRbQmHLNjWHcPcN
OYzMKSXXRLzx1wfGFRR8m7KD3v4QMRGSkA4YV2gBf2A7Cajw5EzxQtA+y2XlkpzaQVFmoL7rPTLH
3sTEAbTCXYjvsS4NfIkMox1GDq04MPJf37XymFAXCAnFMwEz5F3v8/CsQUJGs4e6wVurlLZkkDpf
tU0Yb3O7MiryEbWO0FC/SzrDYbfy13tWoAdNqn7aSGzXerNs5xxCV57OD7vJNEmqJrrXjKfod+bW
oZ1V5WXHZbM9G8Pm491tZhwwgnJsZpwBdUXq+0TL8hSG9s8r1CAdqJhhKGbg96SLY3lG6Y64mCR8
jLkhc2zyiENETxixgyep/Mq371cuQgzrUtr4MspsGOjGEjvo+4igdwxmvz3Jj1e53y2cXMiUsibY
D4qMMtiA9Onf82i2OzdC9sjKlM64NdaeNFX+u6y2gMo8qLnAIKNebq1WjVVhbbYi1+aLXv4zVhxQ
YLLL7Hp0PjAFO5n6Sw6PP7c3NW3hgz2CZ6eqGtBAUEvSJZXW/AJlRuSOITXZdjWotccPt+7Xk8j5
cqXOcZ9ApgSzC0NYKS4F8TtwL1JUJtFRKkdQv2nSF/X3x2PlNbB3jxffGMF05tkvgRIeBE1v8IEH
8jcFFxc/H55KXsO304HpftutmCPRpg4tHm4xxaz09qwRBqzddyBGGmk52K/DABrBdcJ5lwBSAWm2
rNac+Rr6ST78ELif2bvDRhWli4nlHvxZup50A+0AO2l5Mzz+ocrTBtDwl3D4icOL+At3+dhMovN6
FKDYTw8W7L2AVr4Qc26ChDaivvSCWf/OFwnk+Cshb8YZBBoN/EU29m0VGHjcozOilYVUQnyGleNC
j+JdgkzTtWdFKtDd8nFU6q4XjT2Y2uxN5C8ghZWz1JsPStLi+epzMSPQILlgLN8/Bb3upsm/tHqq
OwD+SSr8Wowj9MxOrsydu3Bn2Nml5IL5Mr4keR8JP4c9vrpViuIk6ofiSP2YypD5wf5kPiIE9A/x
vlvI6QaeqUy0YADvZ6L12DIVcybrOeRDBwtXzngqc0cHgbi5t+7d+0gb4Li7bnrqCrQMFD6To32v
yf59UDpl5FZOEVk97pMcnPYMXsohtpoQzlk7iFwPaOidm43PV0fw6lihOh3skDf18EWKnyT722Rt
1LCz9gQv1hR3dfbKtubmx9v68VWIAZxTgLCqLiYvq3sOlS/Nl4hcHwSfDUgMClWX2C63XTS+41Gr
QY+Z3P5BYVvfxc9e5R/Ci204HiikZ0ODco2ZvKbj7AiSsWRNAuA0Ef6IQHvnANwsPOgPuX1VXjJJ
WEukQtqiqPAkmGXOe/EhFKzR1V3rB58PRF5l68XIHnHeqqvvflZPohYpIGKga8QbHFiJY3vDJX8Z
c1GA6nI/j592ppOHYtjqe9gn/VRz22r7csd8z8NpOOwcVAV4TFucugKjSU0ybN0O+xrW6bHvRthS
H8H14iwIagHQXS08VlUCFNWSjFma3c1n3PncP2eAnDEJTHBcMatfIoB5aXWOqNto78ovN5V47cVy
wkYHOVtn8fvNy4RAXuZCOmGFRk85O5pAxM8shls+CKl8XtJxerfUeWBsFGIFY2MSmIGPXfHDRMAa
/XnCIOhiuETeCPihZm0D8IaG4QuAoCnptYew9lEJov7Xyn9zEqwF1GIFoxWf8zuFOeeF0QXKfJCk
b46SAYICFOJOjpKo7L1URX+s5Jnc3fyDNfO6D6RXmkt10/rJ2AGRcBWZBZ7BKKYR23CIO/UgrI+W
5pPApOWWWysxFuWjLvPlXD9hFkrbhgPQANnkA6AyWYO0yoA/x7VxsV0CpPU4jhcC4fFL1aoOk0Jy
S0QoikEbUc62JYkqBHXt0Pdak5R9Yoom9KM6qAuKMcbfHETJw1Jl/nAjGlTPuWPIJaVPZBUynunC
SMheORiMtcZL6NPBf5DNpRuJPpLDp53qIoJG9y/TLvVis2QFPMEYy/Hagb7bOi9AL1NJbod4G0Cs
4gRm8AEG7S8p8/ZKrYB9qOLtlkjqJv074raK4/MLr+nY3TlszlKzB/A3AKHntIb3t7BxmH1u+xaE
H7dJBngXlifvgDJdFXfIpcMHP/7/8U55AwWZ2sCwQ93UFR9/dLVFRde5iu/ywHZT7tQCAEItxtGV
KWJpxVqBF0cQx6OIvg3OMARK34ZdO2E8BHqFlt92dop0Og4U0rgG7p1rr0PCdXEr0OVOuH4+K0Q8
EZ+dB4dy0asp3kR8gpq/Q2vApUuFFwT5Ui6LWzUur3qZ53dl8VYuzC3cBzm3O/vmFZJ/+vss/amo
TmCodi2KE0nnAB07Wadqtp/BCWKmZzw6h6YPCxIivXtHbFi20BulRtcsHT/Ui1zHhfsbZt9xIa1t
dYJ6E5ec+1CRZK3HAgUTDGmT7TTsKvO9AePho7ZAZK2BmFNzzMKMkBpQ2loiMwvEiCjDEoFdzdZV
WhDlqQZooJpHNuk5YvMJOmeyivHTcZjbiNePehinjudyA62LwwJIHQW6XC8rohlSSGz314HG+JX6
1s2FUmWRUH9tQByCY8GuPeEhcaLao1ENqv4ie4mft/ymJpsucxytKTcBFVP8b5snTNQNKg4jStTb
J3l8caZHR5VjLkUuqPiqTSLc514Q2Rx6zlWIoaYmtTmGirnYYs+kQpAcPDyCr9osk3O8LM2g5GEi
+TB+CrHVCUhomhZc/Mo+HSSHyS0ofYWr5wcbbyfTpWWgd7PcBawtYWGwgDOTY7CDuSd4UiRdCGFu
eas5XV6z2pRu97ijkg4zw89e92EpPAyXvH4mjzRXsmtivE2OBMCiLvwt6p1w7TtxEz0GKtRuAYAG
AcBwf1019tKY/0wVeDw6pPAZUgqZulYt4IKDJHnIpvntFtWU+Nb6EnRjxNYrUsN2uTvqOZqp+9m7
wgTacD8igAywmm7wI/1SNX23ps4J4bNyJnICcMIGrpJDDDcM35LNcRsBQeCWU9H7b/JWdaYCuWcv
dCVHoD4JzceiExtCAa3vk5yYqmSi94RuScTXJpL13Osor2/nzoOjTtuAz1kFxVRqyca7FCFc0HkR
SUgCa2r9kpQ3c29RwThyf6BJ6IdPbvZ7AIrFOs8FuNk7XCZARoroQfWSVDjkeJEX19a7citKCJz1
S/6zJRzaA//ZvwEts6KYgJH5Fm4wW4TLVjkOaN4bJ377uLf1FimsvvETxW0WpQJhTl114ltcgIFT
85le5HG1ZLDW7bWT3qYTqIDv0p1CkIPjYPKbRYUwW0KmVGVsHAz8zTpi20qvcMm9Q+z1G24Poo4g
RDWbRBXtsX0EIUC5gT7eXDUJHGqJMwPCOcAX1nMYoz+I74HN1FnY3bvVLAGysL3E1FEdk96/4bop
2tT8tkU5TPxBCC1cmor8xE8m+RPWh6M9uXuVl72MjOoSIenCGhIJ1ReyF8aBEUxwLCNXnxuuPGax
DGuJTeJSveK2eXJ9YFwav+SxLv962BBIUGNxYQxix3g8zCe7CR6wPquXWj0ORrzcl40PZDQEFWgG
AqpUmSQjfNAX5NkkiJPPYxyt49UcWRQXwHLeEqRws11THjgW5beNNE8mWxsluq5E7pLDevqk31ts
MeIrjz8M3iWvC6sBI5duENsTfRPUMNFp+KHFA1uWppfmKBAyvRCHEEzEcVyVZRpnztQKqyIPbKt3
ssvDQ8YbMembbDmaevtvULmOCkaW0Drnrb7COI5A3fedi7lzYSoo1jrKYSQkwEe7udkDcrM+M5BO
i+5eX20YjMRa9q8je+LXfKGAbXuY7BfhpfYyTS9c9r+Ue05tPHMD4JnSPPy8+iq1+0N1u7mODiAe
gV7U1azUsjARTMyjWNCB/ikWR4QB7ndNyyOMzDuA6LgrvzY5bRv2pHahLqpDg932sNhy9zLDNoQw
Oq0LNEzKfFAoQQNpPfI5t4IvdNveSSFY+W7ROXNpvRaxodhGNK89DShmLBXCusjct4TkadanQb3V
qdoRR90qSLQ0m0kraRXURxdRVt8WQEKfb7lx+kAVd0SOQznxFWu7snbeiHXetxATXQxabzKlYG/I
PRXfmUSGqaOE5bCUlAwUndN9LByNnchWGic1FrqRfB0rlXk59ZS86dHrqOQgWftfFfEgLjBhHUNg
j4Tce+96N7T8J1wnRIgUm28GXl2cl9gxrjCAtFZECRVTRLExpQiPETTrvgE6whH+igSn5cy2Mm0y
SgNFfKUZfxQeRcRr/h3hBJ9I8vGyznYXijQth/Srw45P8PVpHf/SEYwcfduucl10kUWPwo0n6WI2
HzLMjVPBHnb7sNZPqN7/oVK5Q5K+Oa+72MSb6dFaCtid8GyqEs/1L11cl6FYj8p5p13ni+c0XM7F
TBsBdMQ2smTAtzrIo7VS63ybllzcmvnkDFqcX/RBrPBi5u3UlsCqTVm1vFY9LFL10b7FA6LeEb70
SMlD5U4AEue1CsR3DEfhxtmpIchGfmMqLHJS/AIku82kVO9kNzASToUvXUp1nEEGwsoeGuE1tdpT
vwqX+0T7MG6TdmnUprtmw528nToZ7inGpGf1GK5yyWlVI13bhupXQSX9mkEvWqAIB9/KqGULsDaw
+ZaSE7zi1yyYD7GElEU4Ghdd6BBJZYPkYsivMVg3Um2s3TKLay5a8ETurUbCzNZWoplVuQ4rvNUs
PNM1+wylKzmAruRFiSXDW7L16pOkMOF9T1tM5cO6hA3PNceBrteGDszij1U9yq3jPcw+WrG/Ya7X
0yMnHA1OiOA7lqGrApX/6Ei28KV0sWKniJO4QIe+N4nWTMWhI1FJ7M5+/lUY8vWA9WtjfzzJ2iLq
emMcuDhbrzFISCUm+ENSolp036ssg4jhiQir7t/yiR3OD2jxBg0YMeQEgQCYWTnkGftweCV+FOPP
CY31nlzHk9r2anVGqJeGiGP9HYSRNOXgdfOu9UyRT6u3VXdMram7Z53ukoIDGCYLQqc9ogfjg2tU
KcjpIboRt3wIGY4s3YNQ5OoSdzVoyIP2dt9GMbDOjj4tDAgeV1F0EVCNg1DrZZZ/9/bMThJ2I8Q5
lxmcHeNdSUnQsiMHOBfOZSoMvsqB5mbKAaMs0LkGhCixvWG5TcSd+XyEP6g/0e2uiwpga9oeKtFG
6ZthTJt9BkBKC4AQVu+P7lWRoGNcjJ0aUFhHPm/uCLRgVbuhwSRRBZgxGZGNltlBJEoIB6ciqA8Y
NGZzg142Q4g/NgF8UvN2vvt3hzoTx5AeB3xi1kgHPb6cxI5+b98LQ9ACHh5huEKfan93ohrC44v8
QxqFtGJKNP6zalhQYH7ngcdHw2Bngza7bnAsRZGJvYB4DU8MnifJdwNOvB3NH4dql+DIa7sZuZJZ
8Nyk5oLFGfDL4VOMKVVP06A+QsRNgUm7RzUMjgO3X4ICorYEQ4/58CsL2z7j2OD0vPHSdeiJwOZB
hRsX8/Z4Svvojrrfsu5ciOooJj9ziDEpdnCm5zAFw3608DftnMhefFidCeK9bK0QJxxgUXMjARIh
NTrUBH+eRZJUK8exA4lTlQh+LR0ntfU+R3SDJ8nZn4kqs1eqkFT1JAzBZpenX4/6OrxUf4nODn1f
QOWejIcMLegm7yQip186eh1lbD5inByQqXIDV1hoduoz4WEHfud/Gia2rIOAhETCUEoIiVXpHNQY
kv0HfteOlB5/nzd5vYLThkbCU7rVDQL7Yy6g75DVnUnsmvIoubcEWjkRZPcpXAVezLez67TDxpMg
FncxGuQCysnNsElrHRXxUsqBifLlCPFE7+j9zUzQZIS+hDD/qT6Pcm1O47l3fnTAxGgkOznyLodg
u6S8KvBrJg2NVvZAl+VD/V757sNDveRkHNy7/jds7+KplWJxGvbUiTgk29iYf587+A53LKmWz7lo
swHSl75QRTyLoiPhPhyNMpjXfROGGV3UHPkwR+PqNe6nWR72QekXqi5nPMC7u6nUBCEpCYAP6X11
BpVSf6a6zVsxnCxla/uP3OE39PQb5rnPFigHX8x75VF2c+LiQBlte1UuZAQ50RaLgEc4DxQvsK6l
+LAP+13trVwjv45SVYShzCafDi2hy8HR4I/U72j8Yx3VxFwT2DQL1Wf4BKkBJj6FaZ8i84PO8ruL
ZDdU8AoWX7uQvo5pFRv6JTfIuSi6/JqxKaH8c1ZNvUwE0zilxZN3vHcDkr7Rv47SDn+VH2wY0u/Q
CLMmFIwtVG9/ldDmjHYg72whsBmoJQH6/8xCtjPadiqNv2T2HExEYUzxV02rF84QOpKw3m+mYlIO
+rZgDYQH6tHc0kduXtTOwAqUU/xQ+wPvVLSVmXO0WIPBjonU9C6fmL/bHKRa15fH77msflUDZ8pU
2VJIruh3pJwjmkWDRa4S9J38ZidA1Y7C0BsSt6RSbMTneAT2SGIjgvRCmL4/Jg6X3RG/XkaN0qIl
iPVaxQUNvqco0Tu2HuLI3vQ5fxvfApdQ9ltSYB7heCqvSgXortO2e+QaEyDcxhc8s9oJN7yaFGZN
Et72p+yyPEzWIQFGAEGeOElYxA6ziKYmY/eigbqvUF4xOrz9A/6fyiriqK1PPrhtVFlLbk97wg7w
/bjtHLon52tffgR7aoeXKq8qRhuJfio8+X64KQlXwkF/3XEOZTLskoHwse5LXSOdc0WlEgaHQ+Cd
ZdsW/ADmG3NeomKbJxQ3CLabJXRtGiugtffSWWB1xz8XjqKWij2pROlWimkqkDEXvTl9VpAHw+yU
s8sLPQf5p44AjbuXWxOx1Xtu6lIZ+uOXSrzzore/h4QiEYJ/CkHkJCcGwO5Rt7QvCgVYDMAh/MSD
OO0dHr04uWjzolHjEO7GxaoDwX/tp2TJXExQ8CMCpmaU5TPCK3vaCmLc7DqjEzQUYWMAoyTQa4oj
QjPtA6KiR1iQSdAyjR7H+nF7sgS2Ho580bwsXo/vnfvZ9fuDI9xhqnnpki5u3NncDzJVrxW75tvu
NxknhERMx2OCvst6LZYOnAXQXuxKsmOHhvFTURioR5FctJOaR2ZLhDw7kUcQx03fHEQhTpMVKYxj
5edpYfW+xFCo+h3+Yl7j+ow6CHI7//nZ15ZIjEM9uwQURXhMHWs40O+xcVon0MWfSxcPPDJXe34J
9nzhQMs9oMMrrF8kWlazbSN14cUuv+wPfw0muq7B335O7q5suNrbvklET4Kh1gpUvgPzyZo8E1rB
0bOPGE4hrl7tEPXiP2PsT91VNn5Kow7KGlMv9079BUVSdSACh1d7B6FiAdN9//APBDjK/30byikG
VrAduqXIi0wQ5KMHD73WhAPzC/laqCxcRaSuYVmxI3qg1F6WQ1of77tGwDeGZtH26ui/7QmlpAAf
VAIyS4kcUAZMqOtlmHezjo2uEsV9ZFLhSQwUPvoGY9AYDvKUtHnwTmUKbILTXjR3yOGD0K+uTNyO
W0j2KV9lRsv5AHcO1987UgIPsz1SIlq6HQL7VDQ1mb+lvx9MAffs4PrB5ZlddhbZrsojjlphMB9D
Hgs1aOtGQWPQ3NNwifkswZaX8Vcpps6XH012Eial+ZjvdgSgd/iaF+qSyxZpQLLZf3PWtgs3XIfD
Tay5ZhYa9vc7WywcgzGK87WHALc8DLK9h2TKZeSylSkAMmHRUwaYoOKj11lS8TXuaCffYVNixsbr
OBoazxx7x0NLcV0GCtN3ACVLbNK0IcWjLJDlAU9LEbKEte7T2KCMuE2YPx6S9cW9vX/GnCtgMih7
iXfq9pfUdtE1kaDE8DjC1EvhYaB04L6YKwvbXrWLup9Te6lzgAJbjAAQlcaMDxXogfsVD42DrXI9
K+WCVzDF6DhoqgbTsW/YkEsQMkf2g1sD0mylhNK4onRY7gn078RGobvDbbTFuDbl8N6jUVCZCSPK
GxuNzuwaGqzTl0iX3xUaiYq+4jS6Gjgt5YlWBJhM27LMygbZgbCIn918XjGGRIJTZlRk30WSghlI
w+SX45sA1FUqoueWTyNDIT1reZJvUdq4x7MLbzPggsyoQX0+fgFCqaRvVy3QLSGH1IhqK6S38ygL
yEYZNuw2AtGalR3O0jc7mJzMawBtssAmXs7QGsBtBIMFySreeBfWKcu+JAm/0A6hWET06L1UNzLB
WfrszSEeaRsUtHLbyDf6fxETeV9U6YML3w4UE1UwmSdKWXLq0sKxhdPr/kzm7InsG3FqG/av2AEd
Nd/xA1j7AnnlrqG2+KbxrzXsmajUN+eTeqcRyyxKIoxwKodORqLyAtu2BWbxtezZl6FV6rjINsqX
5HYiYCJr5SL/YAQPFPwQPpUip8UHh+z6C9DRpEZinhZ2y4sJu9PSdT0a5zO0kHH0HzTW2r+F1eyV
ok6xxBfCZvpfQ50NZEy1zXGII15DYhE7OQa2cNHs2ZG6jq24r8jFNPShde9OOj2Q28krvrCsST/m
XzsrAaUdjbtjEKcHqa3k0/sIiBIrIZIERlYHDuYwjtOyuL2JGMfgoiTYxPVzHdLivd+enXLHK3A+
aV3+fKCJXGtxc7lRZEwyDM82WLDe63/tq4WgzOkif1ih0hjHMZvn5p7uoGtSRaYzALQqjX3bI9Ln
V84ZlrEWWhkHfhxGAw4w+2ghoU4O0XaAU/kukMMcCUvv4kuawJ7e3Zs3/M/uSFM0bRIbEyCBAX4g
ZbaSnjtt1gRAEtXW3hqNl5RJmHfwMt/5K0mS8j/bxJr19ndp8AWp5UUOvkS617uCSVAOiaDGjIYw
pZtJOvBUh7MMsTPK8rs2EXew580ZjulhytgYpYoYmixxKpQfU3PVOh+SA8PfjqLTCNad4ITr3TdP
X+i56PGRKPXJOvIXUVEusCmpCRsZ9VcpwT0QKCwRyV8onaPJykDIwAChYoFrLcCCiQJAJB34Yzv0
b7IN8FyJA97ULjMyA0O1pcVtGW41wy/g/MPlDaUGDWjwFEC2j0eb/HcCSSdFss/tlXwOwbVoKcma
ecVtx/W6Fc1YTkg0e924s+vkEDIJivCVMnE5n4fIlYcyscM8dxM6YfOL5S3qPhbPg+J0hLeAhsDq
qs4DWNNuapkm19D1s2sOVOS6k2yQQ00qBusDl/sKIIRkpxaX0lNr5rxIr+4RUgLn218/7vzrKopr
xAZX4koPs1mUyCR9/CrAVPfRnSkig/YZ4SRqqhDW7MRalro3lrNoDPXM6qLT9OHVwktAkq+eSx+Z
NXj+PEbNmbKYwq3zACk6va86SZisjlN7P2qFXOVdZgbkrgRnPqPbFTFuDglMulSAecCpJygKtWLw
tGqsc7WA2KRbkMouQd8zNRp9T4CtmVtUdlwy/tBUnUbvlUnPUR5Mk3YE59qKyYeyR6c8MHPzw7q0
dcDKmxj8lGNHMOM1haRXtLj3FejGnc2rFcdyYSriNFZ0PdeU7Jm4SMDSH/Hx96esVozfpMbzsAZD
ho+4PWT2EuOZDmsNvkYxUwMRvJExF/1B3Tiz03hH4FOo0tauSOIXKEJhLM3VjiAWqxlPmHNVT/oA
Yw9EcphdgTRo649K9JFD4hc7sIPyvDdMIaT5dVWP+DVF3qT3ci2LT02vAM+9GM+4WNmEnnM/+lXV
oKhR0mugXFGJZ1s6VFfopZl1MaxEQghu8/DPCZU9iK3QH9y163D25/hGw6Of5qs6rvN8W0lB6bTz
ODr1rid6wcI0MIMyAZJAXeR9kr8uPPIAx2NKQFW3Vgt/A31wWf95NNDygNsquWf6tAnO3glcyhgb
uERY36AphwYMb7po5jn0vJrjaKuTGH49DvVApyoC+tMCAkQNmDXi/RluIEelNq6HAOr6F4KW78h+
FzM+YxIlR+Erx30Cn/+UMy/othQWTWzkd6cuPAseyKv9/Xaw17V/d0EvPSyGrnSGbwdGYE1MYJ5D
MWIbuRfuFIryjJAR2CkhfKe3mZcj1UWh2n131zyBJMyqoi5fN/FhxyDmzsa6A20DK0NwP4LZgczH
bjzbFvtVM8PTXS07rmEWliACYhHP5ZB4O7HdJF1ILscLLd2XqJP/WcSSByAlSzBWFXb+BClSMfbK
CD3RK55txr8dloAoHz5BK/4eIzIKUybYXp3zEmB92G1aUi3uFHQC8iqQgpiqbX2ivnogZyusqadi
Qx02HSlm3U9ibC/FM3vDRC1PJUzpHLDVClnEJdZY0xzutpV4LqsdGAUSWozV9FgYzRPqJFlQuOnt
g7QM8BrNd5tUZJZKOyeQfb/vPxJxGmfwLIuIjrMmPpz2qXEaUgkOQ2cd/xHKlNG17141SybsHCyt
ZdxdeUvTkQqxTglvc46nseRxaUXhbdxA4c1RgngjZcsDcPSRfnrFxwWrxc0G8sXdHXOfBwgDVuPr
QmgKOy2mHX9t8aBmo4AofVlcUHDEurEtB+0D4HCl288OGQAZb7FjrDfWosDGymOlGMTP8sUZz9mO
h+/EKcghvZB8jlJXw5fKEW9zpXG87655wAaJueD4ST5jSsOTkP7DSlFGAKG7j6gMDf/GLrhzqT7O
bgIEqvQAlhB2ZIM3Q57MphsEDcEWWv/TYsZgngb2rEmpzooEVS3LYNtb0oqWWLEf5O6kl9wQKLzU
PgbVy1rpin1CLvta+IB/tPch06T7EgoFl65w/+yt+ykCIRTwIo88Oc+XGsSnH45ONRttVk5vNetV
aesEoMJ7Sd3M89hta3OLO4CG2e3aqvyvcMPHW6LE7XWKXslgfXTiwIqUtLfgTGncrUdPjzQZBOgq
ESHNaPpAvXaUNlFk54Zokr72DsH0gOBVMW7mthmMNpV+IiPQa9Byty+0VJ0SqjaXEvy9uAgZhqHf
+jqrOahBHX62FN4LL4XAETaKWb3ovV58cWPi60TZnrOOL5vPT9EngmfxzMV5vmlr2a+XnecG7ZVa
XSvZ3U3JZgeON8SYXDdHPQMpWJQ5FNZwz+mTyuRIUFPi+pOdjrFoffRFMpa2ZiK5bXwP8mKrzRRh
fDLsYoBK1E3p+77KqYu94/SJu9DE4mqfkJJ99ZGXkO26B+ENl4k/a0iV33VPYOirpzWbtusgk1fz
WwlBcs+wZg7kPEpCdnETEVGONA3CQHZPWbsqH1viWDxhX63SWrLPbje+u5hP4/dfcoErZbkXyHkS
CsCy8G9bEI3As9FfQjO74MS3ruOCM7WlBUDFXHQjKdt/ykxjjBJESlKce1DK3sae7nwkjnxPy85A
68hMTkXXjMrg7q/yP6Su86BNxKP3lx23Tam2dNSLC2PDRf93SDeafwfBGjRtti0Q95h3MCtURTNR
qgQf3l+D8rgqJ3KWPmfdazHvG97bu8kOjYKQeOrnGy3JoH/y6jqqFYzO/6cK7bzrNv51lEZ7zFmC
OXNj7GQ/ROYAa3iBulIJPazxotioDn8TKp42mOjiUlt+w5zxC9+nYX6C824XabGbnorcvz6m5crN
Z/c7WjM3bNrO54NSW2mwdbLD2t9UEgi7Zjhu5/8E9u3pY86J94zZ/7uIR9itL1EbQN63duN24Kdz
VCHw0l8/Skr0ZigaeW0fue2y3sKUfDOtY3UKUcia+d3wkJGxrZZ5L/msmJKomAXYwECb7LtgjylI
LaftjaGsHVpmaojrJZQqEM1nbXtBBeMNkho9nMFADm3BswsptnR4ZIa7qaShgGaqFJvqqtZtf/mf
EjtPuu5gQ/I4J25li8F9vSEjz5UcWiwMPxxJ3BF5BkSIyZzisNfJ6mRyUy/iXpuljJiRgXaiekKc
nV8JJUfczN4t7p950UOFC+ePsw5sEDYSenpLx6D2RtaOOxG/3kLoMB2tr7Dqf1OMDsGTLQKWm9H0
sHYP4oKBzt06OwoDtNuy5jhRx6z6mA3it8d20KGyP2+cFO/7sIbseyxFuwnJxGrBbeOUg+CX5vBQ
IPr4KvAtCDuxWdYwG2vlAj51htGXNBv4C3qTyJCIBaAd/UB7M5cgJO6ktVQWbZZCzYQQgAAQ+W+V
FJP4BrP/yyQVuP+reheA95EThI+h6LJNX++ekWubmwCLyeS68cBgicJdo5EAK7f49UF4/c5Za+sB
iJSM5BnOpSSaRJx/iKdUIr5YxGjjNR/n/Jl8PzvzFw74cPpgWSurEdHFNiK/hgoBo+FX4EKiOn9+
Za8Aqu48DTda4fja6+di3FASdaRG8QrzRUqsVkffknvkMpeCt6T5J1p1c8wKGN2iqV147ou15qvu
jgTdA8W9cFNUk5kROU050JA2F4j0HxA4c5/8SPEyWsjY1nWsw+lM+lC5UeZ/Eqni3rSiaYUa+k8p
4U2JbjYtjNJg6Gt2GjADUUuJnEnWNbsbQj56oYHyMlG6lkvk8Y3K0iZnkG4J53pCIjJr/B5ef6Ur
fgJ79IUe6MvTLqPOtd8qPubQTBZ3tGArFerMM63ncGgDkus3tmm215uD7Sb8ky+f94Eh59RIsP1q
rpraMzxlO4bCk8utnnPcBVkHKKFOQAySNMe2ch67pD/V4IXSn2S4vl77KzaQXA6GRSWpmukJDQy/
wt0fGtvvnAho8nTFb/e1nmlJ6xVLssSta4WOKxPI1FdlHMqYw8Hy52ud2Zc6IWobExYap2la9NVx
P7UxzjTSk0P5BKmME9octB+XyDYaeyzI9dAwi4rpjzzTja4i4ivEJ/ML3RLgUxjKeXsWEYQWlSYh
J59j0zYE9agcrVzO+vwVwAlCnfJEuLs17XrTGn+rQ8t49fFLcOL24MqQBYSOzzAid/afAxr7w5vj
GmlfjYhCBtI57tgQjvyxfGQttxaRds7ScKb+9dxXGxzjGuQwuTqPGRKVPbC8NLQdOuXlOtv91Cw4
AmxpThu5T5glIv8cXKKWeftTHGMWRB4wR4Vj2NOOqkFzkcvbjhuCjYuinPsD09InKTkmr0/hgY1F
pAjkD7Ust96gAC+e87DBcLzvoIuflCLvO30/qdHPNb/9a+IyFp+aABVPQYrEYFZ10OCAN0jSQ4M1
U4x+Elj0ZdfRQpCteMoF5RTmDF9AjDYgi8v+EZ2zV5f9A4qqORNpnHAiEg+4G1dgp7ddIZc+g0N4
OSYMmeSL05RhdBwXElmvVqbILTMMvxrAOMAeezyMfKxG6S+ubdLUq8jHZN2tZNRAtk5QEGyDfDVp
n4UJZ8iUIk8Q5eRP2T/1g3av1CtZhs8RhmZaXccUPDRg4EqIcHKc+vYcDkI8eYOQSSwf2j21L5bJ
z/EbvpwIf6pGuUtBm/4SZEdh4TEkQRBehTcLEtjyQWkXVM4TyadcBde/52s4VO475Mn5rdytOPKH
7rwy5/IBvRlhJTb9jysCmmWr09q7Je2UojfRKNApIM5iu0K9KU1qej33ufgua/LAvoJP+FUBEvr1
BFnjzkYc1S0A62huOEcQQ9hUWUr+fY8/vzvsmE10CbeGylOLBU/XOXTv4ncMpsFmEKw2Olv89Vrg
ejMowyTGtfPXH/r2hG97wm8V5W/pQiak0eSrpBjW1XNCoNcJ5jg8JudgqytJsJ9GO5ANgfk3l9HO
h/ruLCOB9VVZOKHY6H5qQohjAhWu1PtfWErf9B0aD+WC/juPVmlTfqei+duekLH26sLEMtJS76Zb
7xDkkKgLj0bEQkz0kwfMFJ7/CDVw2tXG0dWjnTC3JhondmS4fufG0l+Wwmkf5HMXeuxQ+t5NNJ27
0dNGXcjHQDvjIu3vjIFgcK0igfbMg0TsgHViNcEX0nU3SLTDXalJlhi14AxMAPwcaSkJ9C9Nr1jV
JBB57sTVxxd0/1C7SpNhJh3EK0J1wdc6bbHYxeeI3cv/FCoWiTQMaxJDWWq9+BYDr6BhFUbYB2QQ
eYibfHswiOvb95mfB0l4eiHlKLOoIdi0+WwjuriRTxj+Xcr80C31U2E7EnwgprlaNu9xzzrs1cEo
A9Z5b2VB+/b/NIAPBKbl6OfBWYwPow7T1HFu5qnLvSXg2LCUnhyWgDLmtvisBJHi698JDrpvEy6T
n4stkI+uZZ2fVF9SvzGvQ53jeNkqeN5EbOmTGeuljzg4QNiI7VM9MSFzZqG/IiRQALTMw6DkBKpJ
vKTizVVaYxMjPH0GFOoJ7D2CDL8q6d+EKfi6T26YTpMQGH6LhH9qhmec3v6ejHN7AIfLbnWuz6dU
bKpzf76MehC4EeYJq0I0A2+lHg9PtuKzMfzVRonRpAjRKZCUjY89xUBAnZ4cEvQntBrlIvlgweBt
v5Bb0ku8442u3cbqSnTo6irC46rJcFi38Lm1g5ZtsGzqDbvuNw2NzlP68cC+ZMTSNdsfOcdFNHQ/
1eivkG1o3ERZJ9sW2rpSDpf8UA0TS1cLy4ukUQUB1H3oAs72MD9cBSLU2cvKHbDEgXVeHp3sWax7
cDkvzPNxQs7ACGvrAx4QvmlNkk51+2ZM8G3wiz6NoVIlCgfXITS1GyQZlT/bjYbGJogFdIhQTyy3
xov2J/Wo+u2ArjBHW1ISfAiNbBvjKBZg9eCLG0B+JsDPmQZDwyQtSDwsudCEEJmZaBWk6/ndRjEA
JiZpUkwn/eZHB1QwZP/VKA9a8uupUOMltZQxqwyLh0bK6F5KZ5tkvSi6qctekAN0aj+r9oMdsHaF
XRhVD/f9hxiqxdbCe8ZDJQjD0U6vshQYyGcxxbiQtrV+p684V/wD7rgZ0/16l/q1U8RXXxsZ9WaF
44JjphFCYOiyBJOIjXIFUnuQTCOmXp8QihWgnGiq6QTU1ms93dLwW5gGJD3QhczMXui0ApjPnDS/
0InsLfkCg780pi4sbHjQDLU0FoJyvBrGqc7HdGonQN3qL0XEaNkSKaTAUpxRX9iNXQWl0DfH91SM
OfqSCPDRmuT1BKaEgufpVJ6j4PSDXh2WgqEyNTtoZESCD7dtEVM5U+hQCApvVmhI6UVbrTbmjUMq
D5kNlPpZlD2KQa++q240ds16huSKAbqpqnnHCE3FEnuI6oCpUPLLNh0p9ocmYCswYBpT+hYDDEaa
5Sg4ACMnp4AbgKury9r3mloRIMvsSqBePGgD56nekvlmTuZ3QMRCtX7QzuVVpP5z4ifM9DH2yAV6
WGinDdNzrNrbTv8djVWCM1pwXiYXwh5YShbB59HIzqX5nvyr/dOmYgncdnTv30RkUFtfj8/KFxUV
jq97uijvim479Q9jXJjXNax8qqA7s8KkpXXxQPMH0EyZ20Ob/gt0VNenppqWeV+j9XROxde9pcYi
o93L6XzCj1PP4fnwKsDsk26Zm+M5HwEpSVmFmZF8p8vrlWTkEemvkfCV8+fjnPSbIVVl1LXWeY06
+mBNLt+X5MnBIu4W9Xhl2xn/zBV0HC7+jnXC0hUb/MI9pSbvskn9QhxTUSgMmFWUhZEEO/i1nEM5
svreSTrpULrA2+/+XoeHfr8PH/nXGv49aK6YLsh+yJhVobJWycxpXQBZ1TQHiuwRBM46uQEEPAPh
twEyYShmBYRZP+7Zgpw9LiaYKcK8lwwbApNDAa22VD6b22jQ3zTD74ioKmazIXam0mwnTtolN44y
bby6sqB+H5WvbntLtTDRL0Kz6kG34MICfU0ReQ6pfM/3WRQAvAzgsfFfyteOiQ7mA9VpD8i5TDRK
ZuRLEoeL1bpxyrEIoUBqqyGRfSjI4n3Mhnls8D3AfxjaIIod5q+/z2h6K1NZF8rYsAvRvsgDNZcc
bwVtZMyTP3ok3a7GGY8vqhfN5J4rAR8OrW4cUQcxiDWCPN4YZMEhZqdX9qTlOPOdkaMl5Edl6W4L
li3I/LNj13UKxhZYFJjzVsmksTJDPCX0+fuOBfYdBtxoSPOankOCe7ntrLSVwntDqsm+SQzNLzFd
uIC5xw46QWhMFCb5oraC0tdPtnbjNBLEebyhTGTj/Da4cb8KkN6m7O0gknstS80CKLwkZvmzL/1U
/ZDgOv2coEVqeMlrVAh4bfF/ndF6+nXiEIUuII9/xKV5t8FNLxm3Zh0DZzB50Tp6gAUOefgtD+ax
lGrcmcz+24hX7oAlySbfiuMuD8KvwzFHIxIfhgf931wefowhshfGvwQg7eevnJylusObwNztTeVm
85OITJg0axF9Vay6JYcqj83q2EdOD+1BRXdglIV8mavvOD27DOFxrDiCnHL1otTTh3/JXPKecC90
IqYG+1oHfy26LutPiuGsdrWWJKBi3URkmrsRGuEXS9t1+g2qnu2KpyiZiMSv+mTGQF4RDdK5RVKQ
68zCV3DJnlHm6izhDLHALUn+7NZyQ/qN6grnCHJnGdqKBD3Pbc+1junmjmg67r8UhwrLcJM9w4y8
7RB280nK6UQT6MnFRlS2ROHQMp0bcJI/GH3Tix1KOQsobCE6kEhq7xakjhu//+iIP+7p/BT5HMAJ
DLh0jOohLDj4rKzl0w3q/aMeSHoR3Yb4mSX2sedDzYNdEdvUymZZnrGgJh1NXFHNKebnrAoGlLuO
uxX8qxKU4ugF3wH8WzNAAbQBQbsNDbKyjfSdwbgMU/YXqvLuijH7VxR7Z4ubHbWGzqqxLNp6f45H
6kTnDC08J03/vGk2Bo95sGfecae7z31Cx2s/6bim3TKLSsf1vM4/HAZWUk5DPe2kfy91TuJAJHVo
ZNprAR1glT49Tu23hkLDN6JqQaelcNd5FxFLnzu1ysSAWv1mt22aQUmfhTnRJAf59QUgz/cx9VNw
hv28Ef9C2VmsHHZPYneGbfCvtO4rb4rdVAvip3ngMwSBffhiMmcgzYPpDR+LWwYXESFnU10mpJez
Ddo9u/5q8PsUdX2wZBSjT9dmKrAwoe7WyyoaYCT5HJNlAT5mmwEf0Vycw/RLPTMRIRgBkSkU7vgP
AlRNfYmjcOI5H8tU9h09tMBsVsAxW3+34BKdjxZ4D220Kj72pAVm0Wzb9Avy+7Z3ZYO75DROUDNR
w7xw4GftwSCoLT3Ut5wejlrhM3sSo1epeyG4OUflTNts2ABCM5tpm8ITN7Jwg84Yo+wE/iTJ74JK
8+omf5BB5o/xPbicHc4ibcHmNZgEognTwggXeg2wKRoZNU2pf63HsGQd57ZylIV3C2aYdnt+udWy
FB2Vdmp7LGwvpKByHB47L52tHVqO582yET7mGCYvdsp6nWpSy7o/q8tniMq5vPDwtd2YSQwQRlVb
YsTm0poT5RzGqfkHKO9jv1DWLNbc0ShK25PD5skZrsJa0PrS6pm+nuGYARfABj+Cbhhm4o9d9f3e
xeix1MvRqPK8MQ1kuxuIxvUSoZqihQfDRyfjRxv4q/PYTY/yJ+kSmJ9XKtY3Ddagi8+mehvIfouk
7WsETB0vvwgYdg1KQAJdFmJP4ZOfw2cYJ7E+/P+y0m8pBTihhCgxXVY13Hn4gT5QWA7MqOYXMzF7
fZTj5shjcccLfKvMFbAe4XrBQPKdbumJ3Ldh7TZxuRKhkjc/7lrcYxybhSPkONp9L7FkXVeuz/Cj
dJgdOEv3Ke5+MKkdcJBWJtvKF6ztvMvo7rvSAzPMj4i1YU/je7yTQiDUidSeDswhDNk4uK17SN8h
yo+CjWi6n3sjKiTEgGDhoCupmYBNED3BEjaiTJ23Q4ULASQF/pasFt51bBqf+shrYOBEokoCN4Ko
DIeJXl5XneFe0AQUQm6+2yJq2nwKnqMK9iAG8eglPuEOYERYjVrfR9oxsWNiGbug3X0Um2T/JTn5
NvziAtcwq/HUGttN9nyZDnnu9XqrcS2mbcvLU+n4t2S/JRa6DeskUTf29pa6kNk+TZ4Cdo3qc+kQ
o1cWX1dqQZNbWEp63IPxWHesXGNPr3pu6l/5F4Sm8lv0gkGZtcg6j897/3yBpm+Q0Xfxkia24GCa
6t+92UCC/WGu6XYtPBwPQ08H5ZLrIJvWeENaRWI4PUQNtCMx5z0aAmMLaMDhlgKGb/SrxDsXx35J
k5d4W7GEYnzhkOi6CxjsUO7P8sAcEhvuFzUwfOyKLZ/kDrXnHf9ksUBTxsTsalsOssFy6IhdOVF1
+HO5zHkPAkg733WEjfrQqKufUg30JtmqAuX5v9MbnTPjb3EX6WMw1OoQjNpUxT1SoERLFbMp90re
0vE0jdwHlVzjwv1TcKbBq6jWGvgd41QMCCLYEAXSxqUSrc/muV+/uFj6dSy93LCVN7Z/mdpuc8sn
po2C52nKlVhguyutIBSgSqgLFVrEJQZopejVomL27lWEbLA+Y/23Q6WKVlmtKUjjS0Z1o5hvbY+4
22W58bGTjpqvkWjtYYiZEMeOlEvTubD8KPQbsBu+Oe8WpZDwALI7KIMhFCHuQHa3MyzQWL1Ydwii
RkZX6CO2XF2NrKPl77PkThh/gmc5a/JyV1ljzaZGI2lIh712OTzfcHz7HUaNcUoY2HCNgzTrRAlV
plfxBlY+tlkXLQqlr3E+uCuS7A6DsQW79ywFBIyKqagzyLO23gMVvAjIepO5IfgbQpgYha+rY3q5
Pyrj5GSPMi9qSkrUqfHXyap9LPg++Arln+28UFC6fFVkhGejH3Vimu+lnYoihMJgvziPryl03Kjm
hQz6rcs3cKJ6u0jphDR0lNT1J6mrQCsaECfXmhpkaqmbzqo5A76ni1XoqNr/SU0E7ZIeuatedpWV
ixM4zrDKHWWAXcxAykCeIHqmFC7UwB9nv0D2pQAHLDtRmmhqL6UdpdbsIv9armAuj8o8Q+XjY/8k
Isvw+4Rkdmf1WiNdh7ag9Iy74teNxQ0rTv4EqdMMENpsioTVm8VL3jZtcbRlXzMfz/UdmDZDSKZA
a/NNfAHmlcTR8z2BTIQctkGXediIzL0xgQWKEts4Z10jnHWPxy5aESGsNj6ZeT714aEcgKSvrCVI
IJUgw15GWjI82u423BCmbRnRAt6soR+NVrihf8jd2UXr3oz0TE5+r7Aco3P8fktG+0ZAjA6JVh7A
z8ClfWc6sTNWQqs11j9UuYgk1dtVat7RTKvqleKC7Ty3dWexegfByAsaxfiAc3IsrcEa1Nrc+mRw
prZf1/sUewZmv0YXzoVZE+alUCPGGf5hdz5zO7SecZruGFQxi6mVOhvI2Ya0SKpVe/lhJ5lFtbUI
JicIpbLjejklCe1GbfO1Tk8C77CLR1eB433EGPlvgMK2vfXsGmV/m3G9One+ME7m5KwGp/DyHVNJ
+uXH0VjSYkJVghGk51mwHvdZKBz11IPoKoZ8Pf6yHVzdmvRNTjURLpTZB5bDHfojyeImhRUJogkj
VQb1x8AJIu2IjcafTaxPhmfjlTRJKESyMkQloOKYzc7nDuWGgMkZtleAMAN/2SM+OlK4dSj/UktP
p6z/Jyym8d0h2Nara2HYEX85BFNOFU/7VuQt8gpEMbgh904TJRGtWDoNlPLjiOWTeW4QgBPwN4gf
/U9OGKtYMo55WKM+nbwy64R4x6yIbJ79mWhnl40cEmZjLlDYEX81cYTEyc1+3eO8doCk2/HYxroD
o+jsnWhXFKWetviI6eVk9rd2mTLNgzMysB8x4FjnLT4QUEa3z6Yqq2VSemwSsGRMP3cF2Mz5/BSR
wqkMc7ZaCumByG8xxTkJ3QAlY7VgfsEfWGiTERECUriMginSkNMnSAzqxdaRTs3+KJiizftVEbxl
C+m8UTkr1knyUXsVCmLDibF/nw7LlR/EzRZwt7a/alYjVcNcgZbUMSetUPAu1tssO7kwaFQlzaiT
FxcjKv4lxdSTyxZM9U/EDerizhBDPGTRcGFFKCK3KsjeSX9CKYsR9xj4YQzpKfXqmYXIGEHh3Oj9
uVfXMaq2WvdwESNkJvg7ILMKks8wxFlqs2CYyC+4TDmzgQJaYvnbYNx43OllRmHvqEIXG8A7A2XW
v8RRUt6NdAXRRjvfA0hY1N3ZJFtUfR52RlnGSFY1IRF+WxADawIoCtO/zcKuQ4f53ISKwSCmCJgt
tM9Qn6rkeAzO+dqqAFAu/kllq+p9hxgVZ373nC+2I++BEXmyCunWx6SODDgUauCBOmYuLtaI186r
xW1wEmr/9K0Ufi673IpMTo76ae+NinvyhYkxlF4uq2C1a6jbDIJBu58rLKBTSjbts/bNMC1DkaqH
+72DpSK4b553AJNZk+eo/LPvFX/pP9n9CRuVeUQ0Npx8KeOL58qfFYRqHAGwZlMMZSKfcnEUIrnJ
F13Dxv4rsQ9vKVo7yjR17a0vK19hqS1dQs52XUB2d/Nj5T4V4foaVr+bR+xKQapiAiSWBaPgEBVU
hQk6pGErO8e/p1rJfSoPQFmV0x3KAAzRiSo5DFh3zs2yRSHMgwDFn+SSQHjSexqdH+F9mFKz3SZv
/1VLNZmcWjIw1OmS6gXX0XkKc0Lk2lYZN0Xt0moZR3SBswgSANe0l07jmsHD9PskAh4M5eBZm+us
QHkN2+F1pmU6NYRUqkn3Ph+6oUwdxGArxPX25MdeBI3zC/ydZJs2S0YDfPtmyWuHGKANMdDXtG/z
3F4S3oNY/V8EGfLTjAuNwnHIPKJNLCBcPaP5f9R6FXkXWSWX2xOQrY5PKxeBmakAbSzGaGu6kjwZ
4qzJlA3sjX9dVGuc8yhmzlarDtZLEvf2RCO28DjDjmPHZtPnhaQGt9LSXpxxivlemcLaKuBjplYu
hSIpZrqAbU3kNoKdxxa0hI2gcKv7J80GOom83KEbcjWQHZTxSDhbnTKlVrhSyk4DSl0BtZQhSVAu
7O4THm3EBk8vtIAZch50sMz82YKT/lSEd9Uybu18GvdYD9D5v11J9MIB5zaFrIvKktdjslnxlEZY
HOzyhdTyUQSsEApHkjqa5MxJltd8PaCsn4QO1x7f21gA/coxXD8bjFOYzYTDqKdZq86t2P0u0E97
e+ESeW4tMJMoI57smHw65HzFKJ/D7IbShPe6V/+MM9Yad3odP4Hw7G/HGOP1x3ON75cQ59wLKfyz
I2aqmTiEjTb4KyevLEO2CWQtiasF+Ph5NNhSHWOmN17lGzx3Eo0lRCAoVi9yvrCz6Umywynf779o
ueqtxkxgXFjb39M81069yMS5Rd42BqZTJTeUxB8fS5jwYG94Ty1Bex67wC6G+CF0zT3y+oKWA4pD
at6UP1M2Zks6x6g+iZrccGdjFBXMwQumVd8mquQNEWpZU+oVxCr1ytHL0rr+CZpFTzFCqaQ3VkK1
1nNUJnceLohZiUlaChJWCSZy37xTWJCg+YjMpJbqV3pVkB2bGUOgLLm6DlrMQZ6X8gE6Lw+YT5mK
VKreEcQPldG9lHAzmYoC5ypbr79mNn312qReVOAWMPsrk43I6p54qfnnF0b4cSME8wDxwpOepJQn
SxWBIvegLMgxYmPomvshUmk2nfjtYqw2NrVkQcU0VWN26rEngC4HW2WCqdZrkWa33Uef7xEU/tcq
8XBZrtbTshLs9ahuQnYX6QAyuC12lRtAgLLaNe6yTtAwKfHTAC6SB52kVZ9ukJrqyJx253fE9Pg9
R6OFg8VZuC0PV7l+B5hOcQz87AFAOcdkRQSTErC2ujVXsoZMMFOdpTiSc60LLe0YtAlg5O5SIWYu
q5iv3U9dVj/xMHwNeb2HZNgvMB56+T/3byYayR02Hz29EisdVsFawZ/3s94p6TxKrXrR+5reBU5N
Jr9IK+z0tFnfh9sNPo6mD/BIavRIQ3wxAw1Pdqg/O3wc3JRkVf96eonotTOksI9JYyNZDbqfTbMF
eu22dq7cAXzV4p5zTVCkRaW7G7qY8UqgYjMxThexgE1Ej0O2eXNyWb6hXWEE+oTrpgGr+sa7mF8V
1mY2Eyf6bCXtP3oN8G4kO18n6ZGZRCNc4wxSSPckvL1u5jW4XD26ted84N69Jx+Ib0sU/4/JLWHr
4CyaAphYFxGbEVob4dtEnjozynlrnhKaZ8fkgP0+5K+Q7QcHWAOciQhyGxYDL4G5AAZ+beHxd/p5
oUieFllkRJjGz5QFl06J0bDX5vb05+cnJpEf7ghlVsdX32AGKnj+yhZQqkNgTjuYPJ0x5JXBjJCe
/qhpzJZl6RwCwEbG/QuVRKp8/qxKDC0EgzvNkRKeGMZHPMAXnMgbBE6qStyXvofqXc9BeysQ2X9w
65HtljUCjUPvnf+Jl0HpmC53Vd6RX751LVKj1SUegVPtk0rArB3Pw5/SdQo0oVQLA3aiEAZPpHNT
Jbe7WFNIXg6agVE9HA1RYzHOSnxLQk16k0O4IYnBAFzRP2oQzk1qKQj9in0h0xVZdW7FMPm2q7tr
VomE95fIasQdrI2Ua7m8cNGQMgbKFD0RgxGIIrmQxEB5VlPHmPRvcCjeUqLjBBAA5FxV8ZODPtrv
z3ZxO8LL995LZNCocaU6JmPhbjldjAJaTJsfuhly4nKM1j/lwZdLLw+61nVPE/L65bnbosho9p1j
lBptj6bMJ+8w19+rCm+S4USEI+Nz9oznbM8W3ki3DyYkLgnkkTUVEm2ebVS3chl2Z28mgLgsWTSg
CIYedh54jVoJ2+pvoeZ4nlCrZPKxLfQYY6Wbpnh5brbrN/qcQuJXD6UBO9x+R6bsAo8d3htq8gdt
EBATMxgsrTcYXHX78anbMDWHTjZ/yRA2qbXvo5mGvC5DjsG1vYa33mJKEOhDTyusKVjJ+X7jFocr
B2eL85Z7V/1yRT9f5tQkPKGC+ulknKc5vme3SK8TZEzVZj1WTu6+lV7OkLrune1DobJ5DjovlATy
eIW4tF11zty+pf8RY/AevokeVj4VzZ1EjhNsi/qs8DVKP2TtwrIwe7CkaPfjdjE4KDAbE6sWchZE
qYTkJrwiyeYvWwPSHciP5dXRPhb1o/h3A8iZnMykvrTM6MDfDsSSA8KiN/AsLdzolS+i4PBNdoHU
3nnxo3/TXvoQj7hHBM67RUPJhsUu0bLL5yhgCQf29qxXLnI+z9D+MXBxzrnrrWFftIuiY0LgqxYs
cE7x14zCJ5rkQxr1G8Ftcag5sD2kA/HJ/eA7x8iWe7LCxvizIsRoRWhEa638DGwBbh0t8db/2lrS
PgsjzJPTdXVoowkC1dEy42mRdPegrCZK3IG7X+Py0yf+in0UqtPNLqzNaUGZJNkZrFIbdV7v4fva
9eYpatGGCr0PxIDoTgqvby4DLmW8O8MbleEX7q+68rgGLOv2O/1FphUxmaqEhw1ObmpPDIFLpt7N
VTLVmkx7nxqrXn9FrKwPqWrIJEJJd29p4mk38WYqIUuJwN8pnVpIowjf+jmN8wgClNGry6Ptf3fT
CMiSzw1luW7fcL7aKs85nXC3CblTPrJ+FiSrM5rRbz6mNe1GqeeVSxEzyUobbulc8bmpWrp9iO5I
UjBxBYGYrfrSTovDIqefNlkRwW5VWpPjpLn5JDR2KfhTQuOXILPApoG+vHkjdppWHXtpOKEv2rQz
GZKcMSFPisqjiDvH0Tr1raXe5+sdEmjMdD5aJe3lnMz9Brbb74QL4lhyUVFwyrFC361V+pQzB2lx
hn5JY5Zzu4DHjyzYoPyXeO6YOnw3Gz4AHkqkbuE/wu5EMNb0cJhpasrgEEuaGJtOPmASa2U0X56Z
4Fm/Oke/Pn31fQzKZZNVSs9DODDaWWz2vHbcRmxcvWFbG1PHNJaDD04VIminJzSj3rqebgZUiZh8
6qaud5nAYzzfbxLCQWlQxs6H+1KQZH4ZnTUnxAK964/35k5xQobwp6LjagLJ8PW5QecCMU+UwCDU
HbCnb4xKxHiUyEgPsKm4h+G2gl34njSYkEN7tjCsnVsbi6JMlFJz+mElAsJJrw866kP5FHUf5+32
pENdS5urNvPrzA1rVXGLWA5Gr/0eXjeGwAHjqWVbpRfrIfqMMk1rOpGKE+1iVaxwN+cvI2gCm3Fe
HpksdRImvYpOmQmzO7VETRnlfBZQV+qWzjESkERSMk5S9gYSGHmWiwSmKi/wy2dRcW27tnwsdqZ9
OwVnoMF9hv216/7OXWAnKXV7l0fGG6Hnca44ifidKy4Mcgy7Qd9Ik83d/BRGSqMtzbimzpbhc0EI
kL2bQQKiYOFz56sxcyJNrr2yLUPBwZBUDaHyE5tCh0dnw4zLA6liY/3Dv9r+zpDtHf7HlUxrYDtF
ge56584dF8nvAXMcKH3s2D7PF0M/sPHnDvrZYl1u4Sa39DsuexESg2FxQoDMD70uZPlP5R//rr9K
zq6etXZ6/yzlG/rHZu0U+EMAO88GDf0q1zcvL3C0Q3S5kcx7s84NOHb6WwQlMcMn341bBy4DuUtD
/TrcM5oIzOZ5BIexrml2kwiCId5j+WNX6fKGOBVxbk0dq/7HKumABvKVeZ3yH4QvX2nhcLofxg/Z
jlmn4utmx7l0Le15/2vz1T628OioVyMqHJU57EAooSDLTgy75t0u+6+HkQkG2UJq+Hg6JjjP5Mf2
rafBylZmeQpDfitVnu7njV4uqJ7dYPsgRSvzUOHiM4nFsWuLZ7gSeEiTlAvakoesz8xTHHSqtkMc
gY/ioVOU94R9OA33R4ajfSrMJcBkIyOriW2vfj5TVwS36AJ6SQCb3Fk/ZNyo6zixXueuhbDszesY
t7ceMvrE73K5lnvxXSabgPBMEW0LZS4nWXUJ3io76wCTSZphRtWIk/0ILEVc33U+3ee/ZHTj3AFR
jkVjt4nPk/EAgI7uQUwaJFaXrk8JvcO/7BV7xe/t4efU2lrKyGH/rqf9uNIk6Nu0PhYOuMQ6o8ZK
Vpa0dvs6QuXDPC9+us8lfE37dgSrWqSnIYrQ2XrnAzokNT/6j/rVNjpaK+JFLnyPd8gM7udBzlB+
qspcvY7tj48sGPKI02efhfhXrelIb7csapQFojS7+qZhbxw5TUMAnii5yDYuIju7Y+A2FJwwFVnA
Ro9utM3RnHPsWhvAIPtCvyO72C1xjHbdHqBFHtbNLBwJuey2ntyBlzl46TeCmgKo+S9MjogwkGrC
8LDwglzZ3d5piVn8Eteuw6BnGYpE8209j8qDhzrA4eN7KttaOlHj6435XPa/lWtqbymNFb+1UZd+
5ebKPzZi/z3X7xH58iIulZ0HUxD6Ue81/YcOmt8y4bY6N0wO8k0PyQSM6UheQDYfnALK4ciYElsf
g/vY9r6BBjcCl3RsTdiQMCg1Jirp4rvPRi0NRHr8jTE5vaaR9unZxCIjyFwoSDgOvT81ed6PG4KV
dTyC9l/DjZAF3uWcGynr2XunM/bklh0LM0aU4idarGhKZq0d3FXpOm7q/nuMcos4uv3XeoFrqK5g
axKfkFk/cjRxuVU/r85g2J79zG4f7lzqO4rpmWvFT9yvrxt+VPo1p8i+kLYwY11ncFAHAJICsawX
AywzdE27UZELFXGCQoOSuRrbppR1aC/MF/0HbWw9nz4hmqSBGoWm1f2Z+3KSeDfgpWgbBKtHhA1w
DUoEGmXMxc1quoV7moRinuyRDhqCuo/LTKG0RpBiOBs/TM6dRke3bWlulazpQ+s9JfRBHz9TDtYo
8uFERdnqe+6Yoow2aehf70WVM85LFRGo59cv0xwmPOmW0GBA3C0bZQqiscazkeGrCCixey+58/lM
1U1mDH6tiB1GWd88bXCXwI8nPFWkOnuJY/mXvo92gWO6RQzmiY1bwWCGlzjiIePhP66t5HvlynqL
uTBwcaYkFakoarV8VfqaD8ySIMRyoDlJZkhAzigELTEXJxLKutMc9XslddyfpP0edGuxd3sp8hvs
SbBhjbkYoRN0rH5O5iSzKKXHXqCtJI0tmoeO4RZVNywfPFJlHs2JZaLjj6NXRoH4jU7mFsh+zcv2
ZEaYeCZWp1a3ycVW+qX2kXbeLNdf5AaDO6jcv3zqlYkXiuUZkLSZssELRisa9mcSwDyaFfs2+yZp
qnDGK/xL3p+i/RQ8mscpXEk/Q9dI97JrwEGAYC7H+jjNxMHDywEDz0Bwhorhdqa1eSaPZ7eDfc3A
IYiUruBG0Ddzx8OlMLEmsIFUe9cumb+KMv4OW4Z+pwLogMpJ49oqCS+ZJ93BBYk/N1yyhJXZNW++
4l1GfdAgrkZFGHdjNgxkvmm2lAbwOztPMZT8uDtD7iGsn4u5uDXlRmrCZjmW4sGYmt2N9Y+SaMMR
DUUGEwafWNRCJo9avfmwond6tlX0GYQMFTbmf0mnQcsvJ7g/iMWd8aEd6JFsavVvccG53Xrolb3t
pDTrc9TSh/yqgHcc7zM60mge+6YufU+pRrEleMzkjXYeXx0kIJ0WIRtOe0iRVFVPnpKW34Gt+TXV
IQmfNvd94hFJ3vGic9dAmkhruApXlusprILxROTTzSJBPlpIP1WUJyTvbCfKeDy/0FOXZ4BcC6W0
5dYizG10giw5+0uL69eVijYyMQ1dcCMpl14VkQcEjqDoIDOzllUyDofTlywoW5CCY8pvvGrSJMDu
qxhmvGGvdW+N+pGV/d7BMNTpPpbsi60XyKbQG2RizgLBhk/uiKi9FJpTUA+RycEILEQMOVrb7cga
Dp8rBavyw6RJoHKb+usX4tDoKaDc4tqKYAma2FStY8NFzzoNPCPgv6i/+S3ZQ3yxmu9f8j1tHk7c
QY6QrzulXlRvShRSQTB4+YLQQwbEC885YpSRsi5mtfcFjco+mt59rGK/oRs1AZ6asMUGTdke/88b
nzidh7cLaXByOtRxqyGf7f41kVN2BtUFKdHbGBEIgPbdi8rm1Etcmg19qZkAy0y9DLex1+q5XTbz
nZyX4/RDl1HhU2X3HJK/MBZ937lCt//Hq0CrGGUrKe6hCHer+zMsZ1Gzzk6Wg8vGmf9bSk9KE2jf
VmrtaQLV2gPAi35pwy5yheoQmziePPmsC7KAcnhteuMDftSiDCNWsPuKU507cUukDPXMNhnDZ2o6
EvDfBzQb4YgB1iElnS47j+Gg8Fo0zi7qjlI0uSStmk8KNOX2oZC13Tn/O34s6KVgc0lL5b30cDlZ
C7m/EuGXF+VoAg5Mul98goyZ3BCoCd6m2OPphNukfIde4Ojudu+SegUvL3ayQ+tZOvqhRLM/JXuw
MNVH7wfXfgiryiZW0yyQzy3O/XMRwKeeGpyeqSVMRD1ZKK/jpSuq/kF5sE1Z3lOp+X4uki2u89kp
gSwWYiFzkMqvIn7Kc2yL1i0274gNrgikDIj1xCO7Ao3nqNo52H5w4mRj+qHTbt7jMYJZ16g8wEce
a+7AvSHJ94qwXTwNOaS+czLq4vtQWwRBke3XbFpadQOPhzfFIETtmDIr8ibAU2tcIF34S2RDy7qF
KOwpaDb6MVADefKi2tpz07s8YwaFplg7WHhJun4oo53kb4wctT5vt9CBbQtQ++rCgO/0b/x9D9c9
GK/TR3aOJiGnll2PaFSMuIq3vbgNTCCO/jWC/Ch//Z5JBa4bUQXKaK8ZZL2xj5sZ/BuL7uaGVh9J
KJcPa8idmjMB54/CvdB/DlWcH8EcafcNRHOm3EqqIlDoT4HZGrwuA0d+CZ83J+5taIYjg5l36N0Q
DKI0fFJSEgl/sZEXS43fQpK3paVS60x1rS3OLT4pVXgoJn5GZqSK3AnhlKzAiIi1vlwPBJhrqLA0
ebS7UFmvlCny97xBS0Ax3W5SlW5/2pzgE554d34e5Db0czjFpPYrov65AzwCscq9jGkPBpUngWTm
ElnbNO8qoLplGNUbFPtogVIeHvtzYNacx2/+25azbuUQyna9E/AgaUKD4M0BsMcYY/YMjlSKKMzK
1tXaonDlsyFv6R+xgfYLEgvY/vMFFqPulpAEVLhlLGczpAgwjuogxGFqP12CwfTEwMN9lWZbmmFq
/IWyUnlKuQcUZi3hK5+nMp2oshzXWOLm2nAZ7WP00Jnitdj5aC30nDCn1hdEvMTe+B/oU3viQpXw
zsnhV4EzUSTBhHrEWqwHSQLPDnXQR7P1S2tZKYTOoSPVTfVInb+n4ow90TH6EPqry/dUlY/ytSoX
TNVFJZeFQ+Yls8eIjsry2vACmXJQvH4bJxmNReiZXwMNz/s8RJGZ3I8YKDfwFfB4qzzFGBnDCtfr
KJjmCUZ1tXHBOl9z/rR3ouqRqWHXfZyuwfoWYewtfTuE98bHi5mV4Kb8zLGEsmgAvGzehNYWlRoc
EF8b4mruzyry3uVSdom88in+lRXMdEpNNb2ehAoCgQ7/qWz9tcqVrd02YQfxX1poSh+vgFSdlaga
l6DB07sZbg2x40EjPeLuqoin6wWjCbXPNQAZ4YQCz4wWgElamtWvCg5Zmf5u4Tczg7c9VBPqQRwZ
Rg7dj8BOZwj88C2usQPM1+bQ/2pIN1LPHKqee9qYipIKFYV86yzbFVAguvjgc9j6ymuinkvPvUpI
jaYeZk7UiiI2w6Sak5XMatF6jKkBmgHx893EabEQh/gQxra0PxaNN4GVi+ioYtpZ1BS8J1BwNii5
SWy5MaZeIduVNuPhLGO3Dcv3bepPjSzG+wT4Q2vSvjEbEvL/2McL/0RNf4JOZGfl6nCnZSxNjCpO
rAEL3tzvLAO6S20fkv4SI94ago4cEfUvqip7hmm90Pce1bxT0yMOhdRWzM3ofjctGpNbpMhmLKIO
lSjm5PmoxK3ze+Tkf4rUCIjXt4M+ZSKcDaBtsLSsrOE1Ihx9QX1e4jVtEpSaIJfg4e/4L2Vlan78
416cJnAi8ByxYdCV0nEpFx7AewSrbc7APs6ZrsdbDwD4prxDXuQCxzwJqxBFrdKf5lsc03TU2Tmk
y06rF3MrCwOEO5qpBR9HexaeaxC8eqgmJ+xDCUJMlOa1vV60qBh5f1WD+8wTRO9G9O5y6M/g1ct2
HqR8Lz/w1l4wpv4xrvOcNm4Lawtqw5sy54PnHrwgxvUDv+sqThWLHpMnOVlrwJO4PAwrawGmrDca
THNvke0QASRQ90iODcl+l0s+8UFK/ho7SKMQGciTfsxazK+k3cYl5hz4PgMXqignOGhfsHFQLSPT
F6y5vWt8nRHZeITT5vcgJnOhQRYMP/T8Nwt2EHB5X03+15S457TrX2WxIO3EmJIwtopUrehiOmSa
bP/pXaqbzRMszfJBWUD414+reJ/I5hUOamyPuF2H2FNkrAbGnaFIWYC/Ou5TsZL+JEqCVKAOrNJH
8wJH+aveNg5zLQcYGbQVhfR7ZJtG6zKg1vEt0upQw2qxWDiFr3RLn/jvkYDb/J3wVXhzN+5OxilH
xw6CX28hNmY+n2M6+Mar4u1p830xCpYXKzN+plZjgUzQ4ahqHpKOxKT6em1anL2T/K2mRFj1B+qf
bbA7HIuh9U8sdWNLQJ3ry7kw4k5RMZGDxqEY7dkVaHIKpNlT2djIlfEU9iYNDInISqJd8hoA8Y0Q
XUR+8VsIaeSzavu3cYWi931f/iLkBYGBurzxS2tzt70p2pNlrHV4hS5ZS59hR9H8wSBMPAH3ipGV
rS6mL/ox23a4VdoPei1oDMOFKp0btWhi1Df4oeRqCBDuoG1hWwTuhZqWnrPsBmCejeiL6AuFWxN8
+KAiA7BPVnajOf7kNSOpoyQPwN7DESSH2K1qASokhzKiOFjKQC93MHDGBRTwRSNCleciFEkzd1nj
jYu9R82ELdviSzTCLVX4kFYODBGRSbtyg4jo2L4aUjeQP1XgT6qRSQo3eZ0AEOH2RUIJDLxLU9Qn
8TuKdkJFibUlUVZA+yQPyxXEv+/J4osdpsWKzl2SXjGIJCVwoI+qTI+KjyfnvpC86DEWYWx4igNJ
dTlEi+d7SB0eWPJCPasEWcPjmoe4Ulokd73rtNwvn22rXBad7tmfXBq3SCTenAoRSGVvlv9lPPWg
5n0Dj068pTvnoFiXnnPE8i5Zy/7HVcJTYWirdB3nEhTzGLZ6J/8YMRc4YMG08dcAAK7j0D24ljxh
na772u9xpior3D74lEIdhIg9OB+140iOX2qTKqi9jBqCwdyV9dyO2+DNd81TP04K9FmXrMTTFYyN
41nkuEf/8gDNzcs57j8G4fViyloPmS/0GfiCayUCgzSbYUxaF4esemoELGQy0oCpdrglL3oeZHjp
/0vaqp58pR8vRU6IURbTKnymtHg+MuRKfYPv0xKBkoLyZvmFwbjgYd2n92wU1JGMzEUDQTC8M8Gu
4O/oKtAL/M6rA+xDkS+RtK+ERf4wy2rKIllkLdmkJ6z71ueKw+R0SweR4pWZ/UQksubGe/xdTasz
ucs/5oeKVYdbL6G1WW0EAA+NRALc9Z/PbQ0s9W2mPyk/szGUMEBJeckysNfjDWV9iXikl/Zryqg0
fSpNi33ELZw7JhA5YZ9J99Mg3hvIrzCV2qRnMumVMsgXtZz9PaRdtng2uPhpf4WeiQRBCI7i7hSJ
QKgZWMBj9BOnwEPT6ltsX3SkRvv3r+6P5WBi5wFAfMv2cm+oMceFZ5iSebd4NPeMMORFjIy6dYuQ
Ma3D/8Esokv75nEY8hDyOPlEsvreStQ5KvvC+omQh/42tdXI18coNE8OX+Fajk6G3F7bwybj+rlN
GUskljN6v4GMllIs02sQbh6m8ZpFMA+adCOtYEP2niWl3yyjfyL/93Fxty0MQyIspGyhL0dIYTPs
s1VVE9cAP6ujvB29IGUU+KY0UpPUsVmhnyVP2lK9Ay+9PmnX4biMANqthUlXfWWnem0zy9a/l3nj
bQxmU7ggvQ9CeFffLX6a/u1vwNlWsZ6EuUrX5jdOBVUc1mlovyWmfRnZOKchgfjdWlh3XlfKuiwe
KSPVzP/VEDiNy/MXW6BJ+HQh2UabyYcq7hUuYmOibZT+j5ylBRtJPYbA6/tET28RALSN+IlH35Ie
ZWigKd5MmC/TgTPrqC9SkK2m+JdcnPK27UKUe4Yl+H9kUakhjGUASVhgYZFdJWs2WxPlbb1j1JoD
mB8k/8E1uAo/uqjeBHZKbkUqXXXScYmPm7zSnKuxLnGHOtsBlhMBJsGb/5hhczL6cgP94FbW2c4h
oGuiIOL4vWBuzwE383Stsr3jOSoMsKqnH8eGE3KPFNbxCDcwiVKxxs49vGgcFwarqcJd5atnM2KD
RUfH6uN0RnwzOhMs9uoE+A/UED4q8IOU9xtcYN6rUQtnL84dW6x6QFGT69ikHaY+MPE8MnrmjRX3
jFnxXjXor76vndtDcq33SKDve2etx3Z3vScaf6fUxUidr1QyHsEjUmr/pMEHhF29CBEEUxHw9ggc
n3erV7NLCfdlJTNNsbbiCqY7BtMELN1Ix7jaDupcXXSZ05JDIJOtTsVO0Gn8DCDNXqI/hq12Bkfk
xe1XKYfe9RthKVy+A7LB+lsLwnzIHeFMyEjbHQ738MjyXDhlW3nl4rgS82UtVOgnx1p1W/IHVJ6x
7h3YXGq/UZvNDFcZFRxAPTsKV/bNIIRz+J76ppQZxB5HT3QMnxJHXqwpuWmZB4VxPEyYzNywPV8a
MSc3d+OfQ3fEiGvxfT002HfNoMhGjEyq+QSVHTVOef++U34Tx86fXbYdanrNbPp6u2ozUgO5wkUz
miGdxUT0aRfKC3JUvUODJrbffV1pFo4zHa2Zr60A9Tw7bDSPODXpM7LHHNkTdD8ZHcFvc59wLP3G
F+dSyM9uC0LM6jzALsUET8oEMqOUIUDNqclAd2+pHWrKQ6giM5gtd6weodBpzpDXgtu7z6YR6H2R
Uucs05GN7PFA6nxkbZyz7XIrwwz8pXQai8KNbJNye1slYkirAWd9GxDHM6QtvpxHP3mQc3ushsVF
ZzvvxQD32UtZ0oJ1bKWdLVfGu6muKu1x2fdh7+8AnYVojE9GWSx+cuklesuNbBn6nqws7zYGdomj
8Ay0JeA1k4Ukk9uLY3eEWf6zQTEIJO+cfy6unY4El9E0Q2Cfu5Ld3ihQN1+eB/Pc2xkamfAwnGQ+
hqFvgT2Q4PByKEK6L7cZAhO6XVp7duEuDbE/sDwQV2KxgeKTYLSiai85ZMF30y0QO1sh8juQh02W
dCjH6RBzMmyQJodFRXjscjTBYWwebMZNShoVlqQm/0/wJsMQfJqQM4QhqtU25Y5H8k+iOwzB549W
03jjcCVV2BK6JP1sX5f/J/lebH4NKcjx58SDboytAxwNO/1iOGTJ1dihk/NKH77j+bO+OARTHIC5
ywNQzguBJkk+ZH8VqIC1GA9Ev0chmuZk7HyMDbr26ZDJMnRpE9xx3qridFxDWd08dF9a3Nq1vr5A
Kx5WvzU5mOqt9ManKxqu2VfNUjIwsnwEXE3YCvsl3L5RW111CjJ+0KDBxIGt0oF7rx8bMuHg3M9z
5jyp5jgB8GqEAdVrGk3MGENlY3WIKBIFKlx8kqupGAAnJSACFde8KQeaTs/xW1lZGSDjaJgKSpT0
O6k0XkCg0ewLkaCcKLbxYa2UfZVVHnhMy9t+Wtc5JT/TpV350iGiFTy6ep5HRhIV4aTg2nKsJf1l
QCaKRvWIE+CZcj/8QBCt2kVUPMjb4tlLXH76if/7A1lEwDhL9cif0RhEilyFtMvHrOSdZCxWPkPV
fBXcCNgf5U2/Y6jUCeXnK/0O7/gZtNKtuhdjfQa2sVEyZHO7vB7atXZp1y4R1ar/YfUdYQdeHb5x
OCs8Nnnpu+TOPfcg8tQqaPRR3HzmZnK25FiHpUX88jEmN6TKU3O8H1vEEVflch+toluHLo1l/Lwa
TTWx2dkrSdQHKHWSTuG68Ry13v5gPKkoh62XWEhewi6zNnU7y/6ow2qoq4vuI1RsbMrYi40SwwR1
aTH2jL2N7npA1UCE/iVKVBhXrV6n8rspjkyY9jBpAZDW60Wok5e2UzfLcnbA9/DiXXps2wP2E3rn
rEbOGSHlNdV8E/xsWnUk+tdKjV7Ygm02v2UmB3Hq7e7l5OWs57AszkR+Xdy8Rv7IcrKxCuS7GHaG
TUkaAH4V9upghPB8RmVmFHa3UK9zpw9lir1uT7vOgk/kOwZP/zJPJa/FBJTGw1ZTBnJdvJMOJIOY
3SovaKWtqs0Yk79rmITpiDpGRrH4qBkH+9k+tNHw0yhqTc357R3uWwbiEy3cwB1bX+75zqnHnzEG
MuXODjZbB/3F//pb9fY25X599sXauxp6GDHMyYmkpFdtx5U+LFpTnLAfoa+uDNjVDLzk3IF+M0ne
SyIUVMSWbMz6X7c/dYnFmTuiOrPno8GqANKm5Mzijjzbs6tqUaCJl/Y+sMEjcl3cEnYR0mETCIZS
v7AKh0N5VJMTNb0NTF93N45J/5LaCuux7+aE5Ox7Od9FXS2T7/nY/FjVhmkA1T4WNwpYduqhtYpg
iiwXkdKWb6xO5pOk3j2KFrZwe3dnJtuxeRXI6McaMWMALqapa5UA7/Rarjojj9Y/e3FwWQuMLHdd
a39OY5ArbHqo07U3MYWlANJWqtCVZgX89prvQiE7Z2hyFayfTQqzUUNTizI9J/2x2qWOKSA8TRqm
8lhUbhAVnLO7jZ+PiF6NfMzrNEzK3AB6JFSIT2zcy07U3OiKOqQXLpSuMYe2k8QpHmQDR+3OcG1y
+AxFmUN6ix2gb2IP+MF1zvM1keqNMpE1D7aUJgSUlIehEtcSd88cROESVw9/BbT/MzLr12kORQ2m
Bh7a/thSEAYr9cTe+oPU4+6EyKCjXqDdCCMh2K7lDg5HAZFMajwM7IrgbxIOisqwWUvgiKb4G4I0
t+wI3fULTqnc0WmBLA0u49OBbDpupR8Q2TmBm3NRj6ELGo23bakLD+VslkdNqORFGxju6FLSCs9N
QNX86GoS4BUwrsLEWyX2YOgz9zDyuIsbbvWhkEM5JBYpoor8zHs1hApSUftKC9THXN2vbpa71aNI
ZVG6y6vpz91yZaMILf2Tizg00H+S6xtrfuxfL0JEH7NH+zHH9ABD4vALcEz/6Tc6v7raoEeYe61/
GXb5prGcCSHdKnrDEPHLA40AEnlPbeENKufTvOvfhKc4clJGP13ai8n9pnMxgSCP0HYWX6+EQiYv
QOkGqa/8r36/eXjVYENZ1uKN6P8eoIY0PbjBG33gNRYvOdQyFEpIvyABIiimfZJwnf8a9x6keHst
84ZrVSGF81fnLbv2rdA3BaIjs5hUqyLY1RRvtrRfvd6avgUVeXR7qB7vWyfw260kJqsLz++Tl0Bu
ndrIPexLZiOz7xJ7o7EKROyDPIDGxh8tewgv8mSgW2SCqW0At7jH+Rh/2qL6bkeFa42rW6NUeJVz
xxurQDLTd0B38k05UyiltlayDYG/IeIkBPLwv4TVoE08KXbG99zNJIDaCLxJd1c6uyeqd2HnbO+Y
ZpKFwC7zkJLqRH5gC0sIEbUDBzghmLONZNOVmoLgkioR3k7ZpcNr++0iZ41036UIBOOG9zu10kkZ
wrD6AKbsLskWHzOE50Ycc+SXr/ERtW4/7q4s7hxG5K2oDY90zdrwLqpvRSC/KNATD7z1w9UTzCBn
CXfz0JmImWXejFY+4T7mFACi+r9eECUyG79eLde6x3J1E4zWjAwiW3qX1bmLR/QgRVh2OybC8AGD
xfybOgQ+Nd7j1uQGpdv77RkQnvHBE52Xi/mv+dyY7MDjVOPUYmcxZyqDmiZ2UA2Zxe8EJXmo57Wr
odDajUUc/2wJwD7I9xzJhRkI1CyCn19UK3khj8/hfJA86RnCt+JpfGvaGY9EO8fYemUuHsM4qVrP
kov/Y5IUNFFDqFMwQ86fkPHYEjV1tfe4k97pRxKCWcvKYPZnRO/89ptV81/YTUhCzKQD1Ht2Dm1L
xFWtaJIP+66HEnYyBIFQAF1XT8G1axLvMZeK71eX1HuAUZoKOs5PChC4TmW7R6+4zNdMMju/iLVV
VtiMpfrMTSU9zyUbs/1S/QVDXIvP3UJqGObA6LIZH5rYTXIio+FhzKlnbR+gjNtQ5pxelMYww9/U
DSdEuInj+SB96m3hUDRKEtcHjFNseCssU9oxIwn0o56GMzgtbTyKBjsyi3lMM73jY+S15DoB0xa/
WNG3ntzW1Z6TRYpGtXtyoJ6x5NVT8WFEn2RpypcRVSokQaRa/vL/k9inyspPJrIecBSawbgTJR5/
vv2sxj7zRGPg8LcxJnj/KbNbyTuWySHkdh+vyPlQiI65N1uKg0jWtgdILD5l1Ewpn7IUKQqNGzyB
6ElDUuFZ8DPlEAmCN7/dODrfeg7jCxzqkqJnjdKjC1eHhcAJO4gFVKpBhpUBUWygOg0BvgepCZ2A
T4qZvgmcLdmr7m1uWyfZwMATlziFiHYftWsrobbF1lyC/sakOEnSIzkH7nSO9XS25/z4XvfcYNUF
TNO6zmbMbV/EdZZ6EGkI6NK1UMxBIOY7dVki0r57o5jj/CbvTHS6Mn1XjVor2RwklGi6D/kcCz6S
HyGAinmkriTzN26d4DwwcTwNePwAkh9rAOCC+ygNd2sh2hV2JdYym0rWUx+U/F0Su9Xx5B2LnHzt
647svCs1Pp9rNUhpfEX0AY3GcpqgjUtAXhkW7IrNpciLhudWyFUBgjR82Nu8LhhbMgHndpF8fi5m
y3eO5Yjn4uukqrJbOwipscxFWdlmOxTt+rjKn+WZlX3ISiC94e2lhnLWFan7b5g0svK/QdKYK0ps
PJOzeead+mTHTqNj85LKP0BhDLs3j5X2wKucSKaCa5ojDc7piCPdssjpK8yKIPh3kGXoswhHCNLz
IUtldfU+ukjV3/PV+pjUxxOOGOphapGSTopKulew0YTM1xrMlWKd8zn+C2aKGcshXggr9UQlKctJ
urQ996OSfBKHEq+siHLqIsCc/qwV6aIE9mmJuiWhP2WPDLOKQO7hItiSQHpxj66srLJTjZY67FfT
yQHQ9PHOJumX/s6X97AwNMw19A5praSNM4J8LhSdwFGLmYFyrQA3KqJlh9vMH/6eU7uedEn5nVdx
WPK7GzyNtRzUaVJiueTbRL8emXYnzChglMDVDfV7xS9fsr+/iKElqTehCdmH2uScTSVEf8JMktkD
NBFaHwvYxESMOPqCVUW2Nl0wvqcE6exJWejiwgfhQyQ7AYmnVec3WMBZ0OHDpHa+J+2XQf9itEpP
nFHYVDDlw9wCHKd6BxGeJ6xZBhiCCpHZzzEbcmU5c0LftfNN50TbBpnMF1rO8iGTSWxVjMwMi5Xc
ulF20WliuVHmN07M2YJq0xz0bjeBEtciqtXcB9LgnDSNAmAYhOt59D1cyxmibCCZ4Mgj799Vgc2I
jVIzkvjAc4gjjqvpLgThpMIcpU+SdyWJXRGHRrjoEknSyfPq93Fb3R6LlCOUmqPPMWZeoh/Ppz4I
PuyQqfT/FFSxNsw66gWwtdd3At0IL0J1OR86bSSGlgvwXSTYFYR1aa8u2bU0kWTgG35xylMT8sm4
5kmyuWBgG74tRZ9hpVvSABkKCuU4hNQ1ABOX5F/A+FE/G1ki96ATdgTIrcSUiUCcierj0VYNcAgt
07r+4nkyM9WgLCXLhzAew/nA6O9tAYDZ/uC+UeOU+6NsAHc2hR3xLiDE1WuwWlPIwQQVXoBIkDNj
+Lq0juPgqIvXnStLc/3J4Oof+38f6Z98NwicPZdfChwUnKyPxf/nvNzo1tb6mJzz9qQxWt1XwLfh
rDivqMDFhvYkbIlaj253Jwv3yG9kgF6nwJ02YCyq+yOBqttXSaZtxHoyt9XUk6qSeHmwohVju0Ae
vZd3fKKgGYMmAIpnV4/D28eGqdrlFmlGYBayYQePBl2EDetFZKxlEmQy2bFDxS8P8xkEtv+nKjtO
00RaKdPk0GuC195BMaJvqgTBu2OwdpbPvYUZY5nIkno/LIIcfgarJ/9/2sOYdZkqtYwxxfc3YVAs
OD5OSBEPPbh8pDG8sT9OsqUDNQQxhtKqtAIJP/b1KuIpK1ufsZWAvBKW6bVGIcwGB2TLbmHOmEvx
gspgleMvuz6A94QcWelZgcPEypGiVQ3VeoY2LEzK+xDsp5rx5I3idIXFeG3k/qyiarTyLcfcUwpW
6cBH1wJb2sMdfMAtsaAUAgUZabLBtl6aynO27lJxQU9BAHSikd8gZ7efNc60hjfVcanXBnGVW/Nz
jvDDwZnfp6iSvtcEWXyDl1bJEUvxSLXjsKbRYAkK6Lgs6LuEdRiHlraMK5xMSvfiK1wyq2fL/oIS
XHEArMOmtfS78xcPcUFvwWBCQXwZOSPKq1PuP5BgWa0NC14IpnQMalIKS7GTZmCviMHHGy5Mkz0e
tNuQYavxe6Dk6saZdHRNAJ8yrtz1wzPVLpaERb5VMu+O7s/K5ktvVyk6O2SL0VAsbpJ18joABCW3
uFv+g3jO7wzTaTSgEmiSbjGKlCUi9ZZEuD2JA6X1RTzFFE2KZ5E7MoxSq+SRrmae65J+q+6AVJYI
zxE1QoEYZUv1Ss14mIg9rH7Hd0URVRqRrJ65n7eGvLMVO9+GO0qk/K09tvdXOb+9gRHLu+70hcZ5
W7pacvyl+VA+UMwWOu3mtfKvxDPmj4enp8ydR+z1mbpIYYfamfS7YafmFuATlWclt3cxA/Pq5vrC
pyPPDDRDcRkzuPMvm87FpyPyPX1hFxwtJgHMKuYhdFCXHWq3lBmD3dvxaoCKXkKx1f5+UjdEiAhj
HhHJVN1jb+SroC9yUZqUUtlHdpgwU7mqwkHIUg3ylB67oH1ZJq5geHsy+lwpQwuUzZqhXtC+UM53
o2mW7ugjshaRDCPowI+zzlRL2/FAFtZ35finjZ5BIX+EKVqVghVG6LebZBld7quZ95ne/4moAVws
mDckRs9SAIAlVeH/D1Nxf2OB7QAj0EjRCJECYYpehOXAHav00PC0dj5QNKXKDfAaHcmz0jGjNz/C
Gs+dDS6WPjzEwUNxpehxO8sE2QU6ceKfmMdi6Mt6+3tota6IgfoNjk+7Kg28ARPYYNyQHMRUHbMl
D3FcEKX1qA7I+Lp7Ek2wVV48d/zVrzihrAab3Pt3AXuKjGzIdpYhZvJLdjculpNBH8obaN8FBJ66
cmfxm5LzaZDJ0e4qIwLXsPqu0S5KHWu8BPQE6gVjqrtfX7c4jFr9AEhDRWzlAn8/lIpfJcRRd0UH
ENIrtWjQirpMr1j9KKf8fCbnpeNNGBy1WKfDcvdoldSbJLgG6l4gyQ04e7mGjj/HUcRQ8hDE2ZJR
er5GNhTnlYsixfVwp86iUON4v2Y9vciutQhTcYK2zdae7K7nGoFQhno6hM0VnOnlj20IhQuEvT29
+E0d76iWEhK0QbXZI6TNb7BQ8UWKf4v4g/mIiFCYOO7QrXWRkabzaOrVJKIoXaLKy66DMvmXcgMP
ibw4m1hwgY8qWw8y8iG2gc6t7CBspP3LJJPGlsYRnhktvTTOytP4uAVi6ovs2Aj9DDetzWriLTjP
+5VAhzQPsfsL/XN2xMVsQdKSt+h28skTlVs+ivL3DPmnYyxBJOo+eYklR1vL+oy4gpqRu9vkymIu
cPo0sxS9i5Ls8+cTxVSMdCWfeMK4hobiHHZstdxBNdTire0Ti6sLwA12In5QYi1l0zgDindA4i3C
5ZMr3oLsu1PChtaJO/UULmPbWiDN4i/IG/620bI4LNrdyZ2diImd7HLR2+CwDOvrs2K+AwlsUzjh
x71Cd5bpd30AEfkhL0qu0LDhpUnaNA9CmBsCZdMBSIPrj1xglJ2+h/JrHSTpVu3hoRToFMae4oPn
ODlEVKMZG2h2hJTiLghpdO5V3cxBjMhj4lcfb5xRrYFgtaFXgbSn6xq0oZriVcu7jwv7v8lMmknG
VUjr6Pp+x0qX1aZhOSVBK9GNR7XPKaOBLAx6IV3zQzAhVSLmmA5GPxbvc4wRNEs/YU26SYZ3rvHE
AbrSWy8yBqekzY3vwOxG2ynK+/eD8Jr4zqPB+ZDZTk5JKVEmSO6GFm3wDnIFBKlhU7TChzku25Hz
ivUnlLwkafw5OgWBqHvwUsS4v7LYi5YXBkNCf6NkOHazBHyphen/gZsXncoeh1CCKPEWSzL38HCy
Hz5nxPaeBmvk4YR0olgJDLvOSVATu7zmSZQW2Pu/wx7CQKbUO1OtjD42W5dP/A4+f68273J5VMZ0
Xt6OCYFwVN0RojhqGaJ0WqfMREV0aTpHPVQGZCFn3Lrw9ZnL4kZ0K9zl5N0nts1su6xHEE5Gib/n
yYABej4+Y4mdcWbivpSmJ6DxuQuMN3hoH3a9FYtYYBBzZcrk6yXK43KuwFxiq4rQrJdrzcUgvjJG
i5yQA6EnemCq69t1P3w/z7y96xZZVIYkxRTEtot8OP5Cz0LDVC1rkB75Pl3fPEC4s2Ugcp85PMVU
kDNjqBLLp2oDvfEiH1c35im6IXAm7xKILT/PaA4Ya2UX+wzGaV9292/nbq4XFvzNbKSaxP01BG4t
4gvxhF3Vh55yvhypyH75JFMAp9y2tntZxp/HvLwAqHLr3OsoDzZq2nD4wo4fnONySDl0aNpIUzhg
8zY0Nzsk5baOGlRTMZ0AMhaGA0K8/d8YPt3BisX4I3J1z080jOzti95WPdlNuziDUlLhAXzAPMBH
jJaQjr38s3S1m/So1H3A6AZx6d5YizZNNyaMzr0+mYkDV6k+Y2klOkKrfMdxyfJ2UYVqupbf5jZP
AbwiJJ+k75RkhAoVLf+3XTO3Ls/UtM3LJNHm4h9e9XtCQfxzRCEx9IF4qaM43FfSlwKkzUMWQRLa
EH1n/23s6uzE9rZoOx3veK7VrVJ+lgZgUVmao2Ri0495asjxL4g4GlEbh+rNpSAeY8MCfVqQZwpc
gGvoVHkXLlJGGbetiixeOv40BIxWO3VJlSh7rQh5o8ce/8RzuhboPOr+Me/XBbG0XPvCvi0jWDxk
zPU3Fm70F5b/q9GsMsptSBYxzy7nZplHBBiY72aIdtn31cmcnR0Sq4wW75+46Z8AWJ8eaGlMA2/R
Gi6eu52ihEDuKo8vQh//K2M8dZ3IDn4N9GgzVMQqtW6sxF8yVpWZbnYl+BBlG9kZG1hMMejIU6Y6
dAZi/TIonCrXcMkQn3XXxikn1tisiYCBsW3FX8Vka518N6egRQY2NCuPhHf4RpbC09SF9kIKJkyD
5FD1DLWLsqgLWIcgAUavJ3rDQI+4M4Lc5Tl9vE04QX3MLVANz7/m8+liRywlvWg/ljIzwEzg0yIn
DgRp+OrZWVtKUsBpzc2I8jUz+EKz6GhNzPaU72ZRH2czf5L5f2pYoz6oM28wg2dbuHHFMHq7xe/n
pklmjN+0UkTSIUlwWT1ZUyReFpiuv/KgWQCSgobyjQiyQvzuBcCUnnQ4w13sQnRoSAmY8WUzuexB
wtIrY/E2e81+PyZFkW9rAQIZYPgfpKGmzopXePCSyEQF4xvA0puXTVDjh1N7XmKx2ZYQyw4pRmEj
Zi0FZZBx0+BR9iT+cbW0OSBUQeplW2ytkTtSbhpQ6OzHLDVKlr51BXPn3j/9qpL5sfMaMXheS/nF
rIFtfTNQTK8OaL0ehsYEgN0PqHwYG/ItyO6L1Ib9W8g8jLuAXnApzxTKeco/ZLPrPJsszmNMkOgF
a6vLoSOWMKf/Q+xY6qP4SDoPYtWltPW5SnlzZ6GeKKVeL4bsFDKEtOeHj/yBYqpwTF1sfos2Khp/
VPCLSoGLuMvbnMlr3hTbEAuM0WjULDwB/Adv1EEqSKGP8+o8GNHuVgFS4odojFp66PCda2dnJAOU
6inCemBox3F6jOlqlDpbHxx+wA8MXNb65IXYBygxXlZKC9KCw87Zd3qTR5N4u+nLX+TdYQFkgVPp
W48lzf/IxQyTugCgbG7/5fgc+oMk/9lAulemrrn2j3DnDAOtqDTrTBQreFXWyuW8rfu/ZU0smJtm
i00EB0GVg0XMDdeX995X+9XAxdB4Up1S6Iebr9e+fNRtruBv9cbtm3ljixcfbqivlC3zZ/GzAXmT
VbYFBDvkbq69NkpOLwmyVzFbayZBdmSnXeMCnG5fJfNo054WWXg11bb+uaVhvCwv5dV45SDMbOW/
CYNYtvyPhX3shLr7Z6FcqIT646QI18ALzsh9aam55T9ZC7x755Z8xQce9BivvmPCDyrBjO01FJ91
zOK8mD9wYuDsjp14bk4jdeQ9wVy4mbLdxgPNJJiUKraJZmxC7D0w4CY/V1PEUWGkRAZ44N1SS+To
XvAALJ3g/QExashsWm2jGYcoHBMfDpZwFKC1I+UViIudVVxKVhvWFaMEsdkTGAHm0M3TuUsfoIHB
dIVGwNMll2FrochIHBWAu8JYG/mpVDzGtDmFKXidY4UdeoaJw0ueOmQroWGHRy4j5FDV2fiouCWE
64wxOGTxvCeVoen5UgxieTojQPFEmzhV/YUzeJS6G3LyO09mtk2XF2F/Gkm8ZXIIWV7MOSbMuQLb
QshOkJR1m+qR0oD+bkNLjqWsNBkQs9uV929wxfgZ0tHAwtIg/ggiEhHTwq/Av1wqKowuRDGtxDjV
uav0JiCN+29eL4jRkPQSvCir9BBtahB4WCJQEtAPZKpQ0RpLr+QdM8feL1myY9KzGyiGqCW6hJ8k
LSfS+gn5AXT7yIehWL0idMvI7mcSt8rb8zEs2Z5URRzeq3rLQpNoGjBIZr2sfScPL3EVJzv7JZge
j/2/H5lkUVXIBStZ5UOzk7keSLgRk0z3xmky+vSJdSe2sL82h+jtKMIPn0OV07PMK20ADSWW0tLo
CXmiNmW+aiKxpFBcxcYm144zEj2mtIn11Qv7swRrWtmZPgSa+yMv8QsmgiZhRrm04OL00S10I2kl
ue9TeXkGBbG2Gw/t4GbjkY7vUJ9m+IOphI5r+mzEk1dL4FVyZ7x01P9ECmRSB2qOkzDJDJsIrDwP
YZDVouNcvEA/+pCHfdj5RUMHUhWfkf4cUrLbqdlo3eMelhuQr7h2TNdGZTk93WCvPkbG43Lk076L
j4ntVQWiJLxRdHiIUJmfDKTpdILT2qS/CBXnQzjE5cWPgxIK5J/x6DNrKQSq6rgoL2bLp6RNek5j
QNhhSHMNNYBbyf2PKZURx6Njd8WLASd47kqvvBMN+2hsf3XXIE1Sz2/d9XnRtJr1YFZyYUZC1ljm
+NKrxChcU5MPcoHh4NhLnujZa49yJhla5XjHZgkQHaf+vKsnJpPpSc0/ZZkEWPPh6aqrpMNFAqme
N9NjR+6O4X0PiTtweTi/JaDxwQwItV9b7DPD0MIASE2Ka3p9mslZvLdkRb/+pWT+urnqmUTrkHaY
6OEc478dTyorG7k+fk9VWl8AgQsVDmBmFP5a9WqjA0/snox5RO8B7onttnfG0Q+4mm29oEx0rODn
tBDZKXrwcxcwNeewiGPVkkvans4+ofg9MZWLLDNtTm9oF+51yosD534RXM8enVzBti+lxxXJbw/6
XK47gXmCSw3Znt1V19HvJ0bVO9yjatplWcCc92UPgClHOn7UdEskiZAgYfvSkzzIEAuTbP738yJn
NmfdbaKtW+5GuP42I+K/J7I1hXscwe7uO7YAKjUdUkXE87l25vatxM0MTv+zSiHHTC6VMsKc3UUk
TbNrBNtj9GoMSpyxxJTDl0ikq3CUcyca8zb8bcYhOFSEltbm5FpsP78mUMUiVvVEmhjOibbQYT9Z
wqaYtfjasOeQijlg5tV9LTnfyL3ft7ad0TQRhz6Kqq2H5o4KjyY7P2UeLkVePFFrm8R3oprdrTYw
5QHiaR5crx2gxLp/wFtFG6Bv6MRmz/L78sGq9jFV/I3/R5sCnbH4ErDmTt+mtYQEfQi2bDEq+oWA
RsI5sKWeDsBVoaTqoxpo0fy8gjcWfzNhKtMUNBC1psu6OkdvH1fg7lgLSm6I+Zjqj63+t6tgXRto
MbA22WZzCdJdBYclRRltZGzdHpfoSn+sMTpG05J37EATW5J7jYkOy7q0VU/YQsoEWM/pLvvZPp9L
CBxpuXFhfZ6sZ93u2FlDjeYf8D3o+zUL2aQBIvxs+CJEuCAIcFhEEvh9rY/UR+1VexJeLh+1YAFn
V6Xm47I9qLrmSCLtbKWn3ZRwnzTHCwKrWrFKwCtad6LCgN3ISaNZVJNvab0vOeF7CdWzLgDNyD8o
MJ5/VI7hcj41m58oNSULOn+UVmBgS2IF+IzIK7j5Q3gBn26FVxEemTdRTvt9s9RE1NTvDWq2GxOW
w24GQHKNzFZBjrv1dZGP1MVuwksaCG97cKuh3CkFKkKMaTlekPzpLqK9jgTksqYEhwVlvbk4p1BF
/tif5dHB3M9x9DfT5PCrNRBJnvTz2hvWToBcwcuoiKMR/uKM+FJO/m93rxrMp7CxyYAe2WP4RkKb
sq2mebWw9SWMb+CLNvrn9S7u3mJLJZTQV0OfqANTgy51zlPhYZpIyg60o2gYhI6UQKjhmVMOYgMj
UGE3D4WNxCznPvLn1pM6zr2XGQYujYS5t8SAHaqoiaPM3Ixtlp4naEH7iEWlqNTYvI4J79OAUd/2
K7KZStQUzTfJ1M1b3VDWUZ7wb/TG415AgJxwHVM+GchnNNTByWqdKkfN34yOOKK20XpdYDflxoqr
GaGTKM7Rahbfn1+y0dPrEpv10nqKwvuBp5j+ECFPFviXl4/bCkRVH4IpRFVN45rn3p8AaIiRqhFa
4Ne5da7C4QWw1Zohe3IWc6TRC2sRtDqztsa1krYlgHO/IpH1vELCqGgYgl15jaf+R+rSuSvlm9Ux
Bu00CNvCvZJQa8eV4DH9hKIYW+1F8JasIm6tuR8LzqlsRnZqY0yKNB+wnr13pFZ+siZcQwXh67Pi
wjgNfpLZf19rZ64dHnGj6+Mh73L9/COK7hBh8M8zrqCeynftej9dkvmIeua93E81zqIhRDsuUjeD
vipk3f+meF0emZnhaUwFUFwWfE+EiZCRRJiMBTs9ruw7C9zIQ7VnWbaJ4l9H70wdrBbN3l/PDiZw
g3IWw0Vy6ByUNdu78L0RxA/xNkPE7vaIzSYlDVfnvvPT1mfmAq+P4txCHNKDCdKPNeP/Jz07mmGu
Jn/gKvpp9i0dIUxQYb8jqR7HObWLPsXB4BUfrov3ZHVHTIq4VArdd7S0gbcW9mpyE4fa0hv9d66U
WgLGuBMR0a1kDoWUoyjqhGu5ehWmTxfeHTL6pVX5049VvmbdIEmvj6j6azbfUu9a7+dOs8melshy
/Ph2YrbxR3Hr52aC9+rN+vCeOfMMFvfo43zAQGFA9WLJdYswXQsTpTSQVOm1jMtygE39TcGSSyIM
wR80xuCEUzDgCQC2sQE5t2Hadgr6nEvGjg51/RnMSl/GnULXM4F753t5BLRrrpvrmpCKeJaOYjCo
2x2ha/ybfMoyU6t17xHUnl5noiSq7y1x2cRVrIBFkxsaQ1UIEr3Yyz62/kVQQ7u+yi7uC2yi8Uk0
XsiuPBTvLKmJ0ZSeIbSu5guhxDulJULNtksRE1vkKhUEUqEaAyStftOCzrXpTKC/gfA2q8UAvY2G
PKF7ZxPkEC4xDPOEKpJl8fYVZhUCdoebwWU7+aocNogyXoUsm5qKTpxaMsalaW0VZv2Xgrr67g0u
IeCPlTYyrFyicv/E/jQ6EYGmQzEhIFZVSJZZOWus4sR8tb+JBGAYn/d6P90YTBVyeodv+NmxagD5
yGeUVMFrdWUbTeIbb8fKfWjtGtabWbkfeJ9QbkXFVNYv7bPFClo3+Q1JiHGtgMBCNtq46WuGbDt0
S18SSP76mUWHcmmiJ57vQP2/Xqyv4bsi5mvWJLdu9imRbVJbGLuJz1pjYF/tdQ8k1qwgMmdPP3bz
M7Qo76Ldou9LvEn2ydEI2C+Ff/llxXoeLF9A8TXXfd0CajJQva6cCIrH9EBL6jLqcHvxYMVrsIvj
YVPFT1xwK+zGmRf2gF+gE6TuCdmTZzr5u0Ur2JsX006HUDqV8mZDi5dJgCdxxsxArA4yzHF8oobh
68yKrGL8VsH/xDHoKD+kjFUb6YWNbva/0LJPBOD7NFlhLxSByGZoJYatwVWpgMNTm3WkbhC7TB5f
4rwJK9pEfiB4tYOzZ2h4xfiIXSkAIk6+Xz5eHxB2Lnrn0CFGeQtUTTG9sGcmObCKTYJy9pWUayVB
rUHPKgkG9BRSRExtD0fA4VqbaofUvMh20QRk4wYhPHF29eBZAH/dTWNSvSWplQ8mab9b0hKzy70V
Ew5lPrBDQaACtKSfhgOUZBGzM2qzgytmsRwhMDWbsdcvXh/40mVYuQB9mLmGRHkDnJZn+l1sW/t3
QAZvru5mv1Kp6VguYrQFIhxzLZicZ7a2TRYrwL2aI7/wb22VWgSDAh6kUThKRPeLLruejJI0BTKu
vKX/RmfvHFkEC4V+CCcUabjJg6wHfls4p92WA7BVpvp+fVTlICIdnaBWRub/61od+cmK184BTORz
3LU3K97mlvb4y9zwc9Ili6jh2ZuC6o1P7Z52DzgIictKImqw5A9ByPv2AEILdIePNjQ21yNo/gfy
EpU0tJsDW0ufcOflP8qbCS4ye4lC2Qmm/O2D2s83AC2uns2V5Tl+wQfB7cp34rKV57HYpH4QOasB
Sizd/fqFcFdaTVkRYUuDl6f9dKSCYvlXPegqMGv8kWBJ4QvPR587+c2NogUeB7BV3wDElp2Ew4PY
jflXS7F+LTQJVuxchXDodkbqf4CGvZohyIQs7p7zpakvlyP5A3vgYIIbHi0zZ5ONdqYJnce4vRR7
pc65Wve8B+n5c7UixqP5ZcAprKwkAADosxfMOhuclL9ddyUVDYSxEADZUuFgyZ7d6ueLOtdDzJsV
0ETnvInelJu9vsX9SiQM4xtGT3+QDbJd5Lb6LiB/PuM3t6EDrEUCFww01dfrzN8WIRKUenTc5Ige
zeBlYB/UvuBGSvnNiIw5Zj6A/4rg3BuZnK41eK4Q08bbywwQcHxDI+kW0bwMLvNvBNQhaLiA9EaG
2+ugE0fxbxt4W/zGL0shEePpa057D1fBIIzPZ36VdSs9/fs9ixOXouyvvrEGYFhIhNwjQuRV1lEY
rln/EBmYIiTctHYg2QOZJevYz/6CUWmYSqrD3OhM7YVoaaUx1TsVsUyGKtb4cq6IFNHDhPMf5HbE
S2ubDZ1W+PWHw+r3gVoFHRw7+X17gpunSnURIi13VWjQsXimQsPt1xnt75T1M7K53rZfsxZhHJSh
GCIXIEwmc62jJ3UhGjdK0hxNAP6Ky9+XznOuwbNRaXodrv8NYqTvKhAEZqbUZ4njkI+rp1GKWHIS
rdtt6252qoCfzW85ExlEmEWukLRXaZsq1GyaEgOIRwnLoa+aSGhbwwqLPXA9jK1eu1yk4rQi4jP2
LnKdHNpf8EXOFBoCTIcb07gsh9+EhxLhxKjFcG56uc3J5PHjVRgDdAwvnZO2Q4KBBd62KhWsKVH4
uA7n7Q04PQFm9eckwEX93KJvCvSvkAS1d7H+jJlBh0mx6N1qJmd9DLUzzNE+/Dk2PuX1QbvEmYJ9
gUxlJgnl2ZVUnmZPMaRosE9y6g6T7e8fY+4CzV+HwZOwVq5p/Br5+3nkz0aW6RWCR9pimOU1lprS
oyiPD3IjACgS3/ZXLy3qCZUjTnxHoNv4zzGcMT7Jq65GTvBbFcVvf6cbRratkYQHrwMTz+pYJSkB
hO3DL+qjqhM2galj0kvvsgIMQogeFLT/MypEbYvFecIfXjjhoG3ZuCI396g0ubEUjfS8Lzo+JBgk
M4Va5HkZiFQKhJBIk7CrUAbIk0MLdRCuds5rVPkK8svqbwPJiQ/sCNExXLacdkNsCiPsURFZkIXK
IQXMWAaK9kNsX51e7MDOPWHXNe2AlPNvoVUTVo69DtjcLY0jdvvvmFLGZactIQjR8Nqm6lXcNfew
K1T7KT4I4z8jpT0z1pS5BddMSKlhCwJkfpe77Fa6lBWVXD2eNhC05Ki8Km0xVg3AtAgYlPEjeKeV
jq0hCg9EpXG3nzg9BU5tcSLw6LxA82udtjI5bqXogcP8LRzKWljwMr//HhGBx3mpsfjUFgWvICGw
T5R/IuJFCA05fEO0lzlsUA+4dGo44lKKb84pzthQU5ETIwo0PmRVX9+FscgJwrnHk+BCA5O8R/Yy
aUAXAHrwTHHeEgJVsQAvwQHjtO3wvOLWE32zsl1YuXZpUEuOjGib+LNCCf4rlUxl/bdheXBsTF5V
cnNRrCQUNTT7yPGA3bdJX1K6SqCMz9qpHFxl7nxQG9R+6MJmeEOumasU/3Ys/6zEDKPnGUwIumUV
NTL4rW4cv1J0fr1VAzgxe3p/zon0fWijUk0+vpVx7NPxMPR7mup+2W9cwWj4dAHPd4bLc/kR98ZZ
OKLZ13cgQRLCZdYrtB1ZSNzRchvApsuIyScvBh43+vBTW1fg+PALcIjtX+Wmsy5B7CXjvzIAKyuv
JX7Z3E/WKFB9bQPGwl03n4C0HsADMiDOIAkDS1MxFavOJh0Lycjs+tFRnEoisGmO5q8XAw8ZQcve
o/+BFoYIzYzmX49LfxK9QL4+i9Z5Dnen23ah35tEVyDkz4DZwibZ1Qy6Izmj4rJqEet7TB0dMVO+
1p82mzbD+AsKB1bwu4K/yqsyPtAB6DwVe86mzRjOCqSFkI+e3bV2mCceMpMMTUw7oVbcgzGRME1N
EQmyVjQTFmEE+hPxT4VxU27auSY9b7WGhvBYREIT5z2LHlySVMV1b0QsZ/XUEZJwwulWrDrll3xT
2GbI3I8/mpJbm5Ez6XeHmQEq9gnob3aneawJLKMuZUI5i35smuTWGyR8jA41/EvMvHZOSX3i+1rN
9QWPSpTGuWZ6DvyE6aRSJwgEokDNASU97U0dPTxevm82lrjTxjgojtTU6dirmT5pvzpUVWftuixH
fJLH/+5HAbII0GWveq3FGH7X+Sa9oHr58waUKYoen2tEJGWO9dhFNKxKMsg1bFS2lJX4HS02jIUE
q9o9Wwb558Kw1uqqo1kVg0cYrDN40hH2bJCwHC40scoVkc9YO+cLDqgHFk9PJeSjt+Gi7FqZKnJZ
FFF5/IAk4AnHdnzdTgrKP80qcPTb1B/VR8FoRhSppdQAFwywTC8vqPSZGBNxfQM4HZSioy+IdUud
cenuu797vO22u/iYIoqCLr0oPvHIX7m5qu6iXmTAmWQpLczfwxfDbnm+mnPMqFFvz4Ni1skyYoXC
iQvECARBMJfIMy0nnr4YFFExxx6U98Wklx18AOgDcB1wCy/9VJ07t4WHBRPFjwiitvd40fv9zLzQ
NRh45bf0ya+sCGlbvCIE+s47/cGVcGvcFTAd91/hYVQavsGA91USBDkUH3mWCj3U3kp0eXmP8lEV
YK6Qd1ycrKxnGWATYrwGFk7w3cWroS41NUCdWzGtGco9Sh2t9RCnSgt9E9u1C5XQUmbBohvhNg4V
tNZ8DLHoLwjJooAWH1ojECzDqAmLx/LBVDWcwkEs5HBc085jUeGbyK3KqtotEc9Y6ZIbkc9iSoKg
Bhy0/6dpgwi5UtySM7ttCpgvWntMmURdKJ8IdCRBudqyHGp7dAvNQaQbZenpDIWaJLb73GF18cph
WCOBxgWxxC8IVuMvRk2BU9/+jqJgPpnG2eME1E2CSD+5NZwakPh9h78fm/kKY/F7ALzc/WgngTo8
CXPtvHNWQ5saO2ti6DkY6FSQi69QK7W0tuZfJTRe8vPm4QT1LdWEK5tJBT4SVXiIn2YdzZYlq/cH
BdHfT82VZU8relth1JzpIT4wt+at0gBAoipQ0l6NSL7Yct6gc6WQGhzpu6U4rOWxfULt0lAU/RqO
wKwWIvRmmxl5T7TEBkEcDjNq7tRsU0ANKzdi5siwFe29a3/TUKcT2Z0V74wJkiIBAcWtpuohY4fV
VFEBEUaYygrV0ayXc51LRECN6oCLe+hfZKCuSoA7r6skwwMFGty88rifD+a4B/0dqsGXgcfodxvl
a2thO+uBAQVK+c3HtfbuXVs0cwaSwkhS4foQ8dsBVSg21sgyygRD5C7ypxLiVEw9ixn17dizhzsU
W930hJuwSMlmuZMAjxpXXZ9FIyu7sQawyuAwlOWQJV7cnJYKIDnqHnO17+iUs8/AvHxiZRBXH9td
4BWiq5taLlPX8ID2opbPSqAn8LuFaHMCeGG/E5BDg+zH3nXyCy3a0R8sJSNCWimabs8ve9Hz3QZb
XO5EgbsbYlqd2RVGTg6KbBffNjhnCMyVEmERHWRFQfRzv2x89aqNtYzHi/U9QMre9pRz8NGfYP9j
MHZ0aBId9tpcRfsEOv54QfRMNl1KkSlcwmpFIMtO7pYSFGlnfh7duDFUSAEioNE7LN5p9gnwNCvB
WFiWLQa+1iYnwiy4bY38DbnGR3k/xcS2XBb7h6ARFyJgDk8jqg+mpBw5AhB87cAlC+DFhkohaIFJ
+/G1mJdHRYI9sCXS5tJJ8ycf5b6LUNFR0Chh0kjMUy4AzFSevxwJCdUP5XQ34ZKxcUfyPOnF979u
hDPeIeod22vwBtwwN58yZafBFG2YxwS5ZX/A8Zpal6u7gbvxtJa+P5dZyXTF8+kqEjS3Y5ZgAWlx
CMG26nLy5JyNA5LJ1XWP2BSKgrt8RxR4mn3z7Q99R+i02MzN0j7si1gthBOeQOkfYNgcm0FzmuWv
jngb8upVf43EIDB469NMavPs+WddL+lmRyc5lcQaHfwG8ifm1gv0mNAtnxXT1RDSuWT3WZKglc+d
j9KhcezE2lFLhhQ+WWYauppvx/klMsVV7BE+Mur6i7V/7gay6e3xUQ5pCIKMYlKCBjW5H49N2RaL
upkGmkl5LIwgTUuS8AymnkViIdokyj9G6IJRgsf8p7+mJ+fSOI+WkpAvuSKmqQMFyUdbw7k0U2dr
6UkpHNmSXkcFGan1RP6zOlKiWC0kv6PrHm7cwXBQloEY7bKVCcaZ4Af+W9l3YEv6Lfg8oh519vIZ
Cw0Am3OC+7LC78jE4E3w+98O6LHLyIOdXDeAr2aZ9gZffFylQVSwu+jS8hYM1cGiJxCRMUi2UBwT
qyqhyRUjuVTAcIy5oS5OrPTv7w4XBma0igL/bKAiw3sZrozZJeBDJCUgMnpQ4k0MCiAY1XkYunsx
nLdYMMNZoGrfhHvxuMu4ItEwgLtFoLkt7+E65Za3aBanUaVbXogDlplV5qDgUMPWQKCuQEMpLxyE
ihzYiX+r+g5FDTRnDsdjMW5w7uXcx+amSJh13Gq8HrYmIlhyDq9YGiM2Kx5sowi8tXluOh3sURkL
Vhju/MHpSBhwF3nRJl0CIWihNjdELlcXrtPnAgMJLiRfMg0vzQF3Da5c14GKydDRNXMZvlDekask
77OLINIZjBZRblVY9tdoJ5zt2N4HygddUEMhePsdx6HPGLENk3M+wbbjQbtFiTizBXJGXhYhcwd3
tTC71SatMilHwXK2vRdwwGKW8eNOyX7Pn6sKScAy5IdWQy0oBVg46I09zZ1lGCMBGSG+SYS2ipQc
O3tAQmaYjn9t6CQzXxKXVtU4Slh/6WaWzshDj6faNmLx8uVxLKe3aHFVuaLa6iesM2k775Yh4NHJ
wN6n2nInTq2Od6cN4tWU1kihyIamdsYxat8wW16lE5TwUXX/Nmayh0dZdWssR+c/ZnuqL8DAd5eP
/s3ZfoFsWiSdvXAvvobwRBfzIZx+sZbF6FBMHCBN+RvAzEplY6yeohr5ZaHQf7Exm250U7poCyse
w6VPEcr9+FZ6ER2x5YTIytOFd15wZ3Y8qfMUf/A3ffy8UK54YJIM3xKm95wnF1BE0moDJhJt72G2
Mhus6n3s74Wh81oZ5HscJ0v2HoEkvI0WLUI+FSaaY11QvflZWXwA2hAUubJ9l2C5wfWmF8h5mZob
9SbD3SV2nMTzXR+XbeiIExYmEXdukJZW2UXybCGpnnRlxp8uhDGoSZkV1IPyMVMgzmjUqk/mjR5n
2VErUgYkOmcQIqkahbnC9FbuFMMEwEKJh0ir5pvaApQNSwp6rh5jdknQXGLBciP+l/HkvGdIfo6e
/iWMpgzBAlRQ/s44P303OrkJTZELubbZ9dxJ9ocHftvXwM7kStZ9FK4pIGMcMcavxa06oxnPbBnr
+GeHjwenIKnwgU0QSdg77u55OdfF4PYyLAXnPlwxhpGdX1hBls0nhZdvd1eS5AHiv+e8/h3/dgKl
ZqJ1YB13zuh/gXv4isD3P1+BdR/fXNfNFsGUH2dCtTcfT005PlWzMm3r7G/10JJt/Y+JpCRQQxMW
bEiXVqRu5COHHKOtbstkMCNAHMs7mtdAVlrUm9E24irXMWJVbbYDRUHu1KIl+jhVLriMJiYRDdZf
5CxfxynPRYBRkAAIEKwe8gvi9IufRqqWGeYrP/Z6lJ+5E08ObJdsSYiYHmHfnkjrDqBcJjozPk/l
k14HNzC75YmWPSJ3C+IRd9V+uKKCi50H5ApxPEOIttOgCcMYMuybdjftYsRVpCWRWIGifIx6V8UO
EYmGgOjHAfQxKzSgGNqiLe3UxhS++yXq7wvjRG0odibFTpxwvmw8kUjbKbM/dISUSD+oDFutVW4h
zn9JA/2T4q9gMb4R6RBTyC8uRxFbH1AS4PqF8K9+qu2Lr1zRCULZ/RZAvsE3UwiK/Wodyk+I521M
2SQmbv1+sZIXuQN+Mj8kuuwJNIht8fl1TMnwVHkbJZV4ipQzC3HfABuDDW8B9bUtZhHxrp3cFNhP
q2z+3P7BsMEgz1JskLbXIb0rpHcUVOPoCkLCYD4jqqA2qcRhENOYJEJFzc5dUw3xFXIS8d50eqeD
UrObRrx013zjUK0FvtbPFcJOJCm5oo6CtpJoFSkdBWIk/wdKKwogfZ7DT2gQkCX7gHpNBRaGmxQA
iQtY77Wa38a2TjA6AWsGpKXdNE0syHsY9qZZdIbGIblo0DMvc9mviTEQvSDJH9nUge/bzyBL2Rxj
U9Ap8307FXtgduSaz1TvXqpmnH4tmb8eREZHL7QLfac/lnCPDP+0bLrS1j8hbVa3sgbtpCvjH4Au
+J1foP+x3pOXb/eAwR3AX2c4rGA9Wh+QKn1nT7EJfD4hFu2PCYQYyM2Yiv17XNaPn7sswEy/o7bR
O2HtF9DnFOfHTyd2h/XozqoMDcaltuxBpBSDlM4X+G/y4yXa6r5tCtBoVCEpR2s+T4tOmZpPCogd
lpt1j2saG9WZaXPxz5OpzS+SGHHaMu370bxMnAi/uZxYajyqLbNyXy8cA6uZsn7ovnd/3/v6bY8I
INCZPM3hdxctBXCSDWOOsfgNzHsIEQTgajgwG8snZiLSgEhU/+ViCp3XLbnPiPJYunivz4Am0QLd
mwO0iOGFahxP7MYp7Ck/Q905XTSorRtDaN1pAPoEGGWeftgkwOfJuzBHWdL9P4RPvQE0nKtXAdb0
FfC1taf4qUld6gnHN9g/ueWjZ1oGy+x9VK0p39IyjwlxENlqpOEAdTyl+BcNGW/5cIYMOPW8TqyA
VHA32vL/IlMg1e6FCkEdMR1VXRwCfPyhNxV5BuntR7PG4TJD3Xe3cxD3io9s3xe1uLfT5wYK2XN4
NVjL9sh69KTw+rsvHhTVpcsqGtElHUe3NGGpdOIDuzJzsdvwjPfW8zSqJk3s8NjgzGd0y56OBcdw
99cU9pgITkfId88hDQJUDYsl9WPhrzzMbTPhq437REwLB7SwvcD+NFjOfvZOD/itKPLA5PR7N9mL
N+PRR5QQP0Com+kIULQ1gQ1sjiXgA0y1+1bxSu7dfRZmAp5zeu8ue6DYoPt0WvTaB7kCJSJ61XbQ
EK+zJMzcySJEEuGqxrg1hdDELprBiikrzxTrDUdaB8xBRj9MGQrN/HjfGm7ota9v+gW8y+KjblfS
+DfaZ8ApEOspxVvs2NSaUqsLML2yYZ16P9A/FmBJe0ibHXNiR7mTfJzDZ7Du8Np3C5P6rSX9i5uC
/8e1+lTtjUeEzqJgVVnM3DEVXJyeGvOXLWWPKM99TPqXu6lWWAWIrYUe9+FdCeGVkPrCJaQd8dN8
DHRNaZIPnSEyViuuhi9IHV4/ZnRJUq774whbxaEHFseCV7eJM7qbvnOWvxtHInsppWVxU3KFA+ST
nnFOM5vxTXIzzwZs9JCVuBhkzkQCXIhG2wbnitzljvbTzFc7y/45Mh9b+ZRNi0/aqhX70N5lWbMZ
yyN0wTcb0r/M7owwcQwBOWFNJWzfHWRJrjTOUIZkchMkmFT6n108C6OZdNhp8GeOisNNyQcziN5R
lrsJpw6QX3VBG6sDRlUKbLgOhu8gkxi4/S2w0tFAyOGH9onCc8y5dgpbII2ODL+3bUdGA3VNAzfO
1IKjF7Y5p+RXUdneiI1puEZmA9UfFW/thbSNkleJfNdVyJvJiq8o5nj2P/o8g8kRKsc6awPxTh+3
qdVSgM2nfgphqw530bF7ORkk9Cj8SAxFrBTqg/7I95Kg1OsfJwVWOzV8M9uZCDSaWGsT2SlYHmpZ
kYskoLHI4MVSBggBCkHJvoWexDgntHse8xcme2BDy/rHRwwCG/ROdCYAnmj6vZjVnW/CkS5N/T4r
pBYZcqWIZJCPTzqRvZp9qyZBGAEJsLfnrohryfZudvr+dRtMOsomvJSoE0CZlW+5iKQaTDehRSdj
rptydwAM+vKYBS2b/4Dnl2foZNlK+gfEQYUFv1V1pJ6fPz0XCO/gWQ34EhhGSfi1Ulxah1f7S29f
VluV2R1bocM2wfJsTBKRBQP/KKk5tlgBNJz4rhsYSO03SeB15VGHMaZPLF92ai1oz0Mfut3yxKGw
AhVZl36FiZduFJOXak9eqkeJDOzceqIvFLN8ub6JW74YkY7SY08c/UmvXey2dbq3XpPcuKu3NnAr
p8E66OTJHwmAfXBXgPGH1pGheAiHVEK+VJ2zAGiMCEFRVf/Wm+/Qf79ETlykhSUgMLb/764D1GEO
kLk/UdA7c/DjQd8zU8/er7V2j/CjouWIL0DUl8AyuG2bpL/9NuoTYiLZyG7pJmzm+5QKyTUsxFw1
mbLq4pMJGr7LxLvhMivasEvc8S7vbVnEi6/VdwFyogIUWuTgmtBajKDlzZcDqyU37AKxUbjOPMPq
DkJfyCaQS1jnbckg9dCP8Dz2h7BZnKOghd7+DQg89a8mJdZiFr1ei4B9O2KCURdV6ZlYSt3dnONu
trWIZ7y5fnBfgXS2amcYnQyCmYf8F38ygW1sNW220pLNHptPBuYx1fs5LaT1F+rMU3KFryvJCQBY
FIkw+Y7gMUPgiAXXAFcGKcbDi4+Z0gWmVPErORnulvE9x+G5eq7MIC5EF0mZBGGDac03HRsCJecE
i87ciwdIgndJNRDf4sX1FGAotEaWFUs4aiEWPL3KUpERThDWg/TkJI5Q9XWDtATOKqjX6zHOZJKp
IQaKH3Mi4U0/o0e70H00ORfEUKCl3/+ohcmzqcEm8yvfaWvrz1MGYCbE56FFpW1RamBTSfBttNl6
IqlBpImXqDskHqeUiAn13ijD49ZKWasKZqFzYUHNYcCgfUeWlYToK0y4LzoBzB5gaobDYAX926oe
lV6tQQxW40fWshkHrMfpvKVSYTF7kaXkkEj/JnAO6yRGjxDVeAeqsZy0gBqCE0HYddfVJpE0a/U+
mowUZKAe76JZeoeHLIhjZvDdk1vuxgUcxpionCwvWo0rMCt0EFolPRtQxe61kOVAQmHPHm/LqfVy
oK5uqtQF76HcOUJxpkYHT6ePALRagovhGVwj2Xc4uo5gLiok8vr7ZjhreHrP4Rm8YoiM4HU1Zvmt
v/r6e91sAhTc1VLLsTxYrAHCqMmugL3L81bU9BTjQlLeUYVURGe0l8kw8Q9/TdFBVbKC9yA0b2rc
PFrRzbG9OmH800uYQimRxZ89gfFxDEniGzwTC9Z2xkmOZSpRImwF0QYQ4Kb6fq1sAr5TD6yJIhDT
lb13fHhDikDywzK6+qnY6//ForrJt8qabtfhzSgRQGkiotZ8RqpTIaEYK17rieesIuzy001Nap4Q
M4J0m33Of4Y9nV7GdhRFHvc/REBXIVPLP4utXb2fv2gZ4Kttwua1NiHzKtMNQaOqzRqXtkyW8A/X
kjjTk6Ucd860lzDHoJTEOv/eiepTEwYmcL1EgChZKGtVWjznlP9TJPjmexg4G6FiE+O8LtIMTyx5
XIZ5MrvVnDVVlkOetF9ZN3HSwggge20e8Dn+WMYwIMwU4JqP4manVwBz+F2b0LwLzpgYuyy6whc9
QVYdvq/jem/XSCtOlTYwsGTwiO9G/DSPsfx0F56gdsnh/4p1uofeu5oVNsEtpc7GpKkUCRkDoZcc
NiIhMyNyGZi4COCv3pD3nG4FQlUeqGdup4FqapDkOHFpLQMZeyoUpo5ppKwaxv9yfdXj1YhDCoVL
ph0QnzsSYRc+NPYfvcB6SYtJOsRD4sbkt8YGNqGHLjp8t8EVrSzUFPwOWm6yoMVZblubuMe8Y1Px
rqY/y+Px2IikBwWyuqqe1DcYhAoPblXYBY1PBDESbr5RrJzJzy2R9DaMCO+2olZHEGva0pcrZ/it
ALGBQK3l8MrC5YiqGlEwI9LtvIIyqKEmFZuENxZ8+GD8UxpfZWgr562Uv10hljxLm3rT78rzNCNy
ceauUm60oF6AJMbgXpdHZ1y9ORANNgSv2GxJ4TtWhTND7pxgHqdK7A72v5t8pwjK3LJpNmC1XVpR
FJnG5pfz9BJKQgFgSKVHgE7uV23W/O55Ai1hxGYP92yITeN3SdXTgq1t1GCaQcLbDNEHWDd1lCQC
WkmCpjcvTkPzlDSG4jKfESYUk4G+8mORm6Cbc44UWxN6X7k/T174FsMlaBaz93dPqN1Qi6NO16Fu
6K3ONipmmoLEzgzWrPRBBQfh+W0pPuJcMTEpXsgjYuCn4fVRHBqJQhgRWF+ut7Wqk7VW4fuHUPhC
dnFgcRDq1L93Fw7jGsoriSrzqg16oj4xKA8yx2wH++TLpr6Axj/rHTdZdrgL7xFVKpuSNaugGTvx
7LDrDr6iqARYtJKuaRiHZVqK1nHmSqjUE3VkuK7CSqCFEd1KyC4eXjdlncbdiW4MRiLOagl112kv
hVxER/nkfOMTalySfpoIuHttb4QPrKBl4ZV03fg1PkXvshUQq7SKTnG4eej7hEW2bR8eWuK2O/2H
6A9qmANy1JaBbQ3U0DtjcYSKHJoy02KPYGh1Q+PB6lp3Jrmar6AjIApb3V3IHfgOPEfxhcDKrJ4W
aQFLgW71rr0ezPd8wrh5M1lb4WHa6OTs0SEQ543Fow9f64Uj9M4KEiNyLDSGBIOQFzlxMDdrBVJi
3rRiUHdDVC7oIgzDE4uarAWCJgdk8D7b2eLb0UmX58gIi4AiCkn0uk7zbJKV+s3fSuoyJAWgiP3G
0XDoeMBt/scDIkpo/d8U52A+qiRTEh2WpPzGuSekcJpLH0Dp9u1PpVBtgVIIi1AYROfjunkLt3qR
YmENro+TfJHcUXsSUNjmiE0j5dXl3xnR+eHB3mhwXoAJJ97tatDZw9lmSoZBKdUateaAWtfoqH25
yuZBxzlANgltaRLgj2+or5qR1Pg6Nn5qz1KIeU8z+4ep4SrJoY9oBIG7UnYPkq+m0Q08zGT+/7Y5
9TceRRQ7nukjC8wfYmISZkTXdZs6VmxN0i5KrrYtYYXyNwe+BdqjeQNxKHeqvehqysvVKYq2oqNk
9AhvknIDTuttI4X13cDiJroRW+5kVfDPdaO/GbtdMB/TpjQwwcgWGEQONmrNMFjVev3kZlpm0vfo
eXqsca2p3/gk2goN8v4x0nfCfJrMM7dFqm30lWhXuLV7cB/1QQYIaJf70b5iKCFHynz4cpCW76uy
9sujs9pSXVN1BFlvVpqaeC6YZfYqqqKhs2Y0d+2YArlT97gilSMVFF4XxS1sLVZXH8jTwdC5zg80
v8LBhOXuDc1lsQFjOd963FdZsgRaH2s7djotEkK2zftlj07BqWZV+5zqsspzDkqxgacmTdjfUgZ/
CjS19gY2YOEzR6SbmhaWRsbbrS8bqtEv8F5kKmRPHigCJDO427YtUgYe7dd+6nM1LUtfx+q1mSjw
6KQc5VqvKdI4bln6vXcNQZKWeGxuiSErw+6RAuzkgkYItK9GOAXeo2i/kZaWjLP9dbGIc8orDkxo
7pniYY8VvXVgPebyrM2I79jg6N0m41vvDtc1mOEtke7df+91Olml0TsGc62QKSaHVCC30pu1GLUX
UIFGoFGAXjB14QCtfRwzcgo+k9ykUavam/BTR3nbzF9ZDqbPMsdKc+aHU9WxDpjMCU169wGt79xS
ku4QLVE3Ceh2eQx2VNh2UHJu8SDs8asp86eHqgzGO52EdPYE1M+ePLJKfk4xzrgUAhqu+26f0Zou
SITkJR9ezDJ7KlbIbDlIMksPSY1vg3KVKmIuB0cysE7cs3nZWJ1U0Iv2aLQMowOnKeJf5KT8v2zs
yiBne7rNH/5GuWp0Ciru/dJEe/GCYABWlI/Wox/vz+Pr/3eyOlSztVFa6R7TNB7Ln2sW+dB/fQKa
9y4WmeyAlIjDOwSyFq8Vz7r1YkdjnA/ZOEV/wpd4C+8fcgVMLH4CVJ3Sc3fEcDwKR4oqT31njyPX
IvDIZ6uUqXJ+EtADrzsYv9NV9kEK3//I/I8E5zISMhDMcSgJEpWnJmD5DFt50Sgjf8qf/JfQPIY3
4JhunGVFnjqIITZzRGjfIY/Jodd0LQVfWR7qq7Lg9ymPiGkJ7bKDXnrDmoRu4SKg8oMk/0ehRRyl
of1XSZkz3WGGLGRsE/f16gjSu1y+fnV0xFTY9PW94oVz+6lbaSphZzxpyvEEDdqnaFKAoR5b3Kgd
/xEX3RcvkAGUqJIc2d/5vPnaU38lYEM2eIrPyFVaY6z6caku5IG78HvUHaoAQnbLRcYZhU3N8UDY
YUuV+8hFF77I9si3tIwOylBjFzi9r7oKnimVgq8HJF2I5RExlQEhUPRMMyvIJlDyvqEYnOV4aAMO
R/pfuavIFa80PigIUie67U4xs8lVbv4md5FnJMnp9bTCbEXvHGX2Yx+gi6GBkbFeIOxqtXSBx+4O
U/HSmo6jPklvuXjmbd6zvQb7BOWuPWFgJaaINGThHfs7Q/RIIXkmimn0W4akEvmT9EHdK5SGEymX
wRRYYlJsLLlePG8HXtAD0fJlyNaS/N7h5SPbqfIw09IXp/gSRYgPdUsZoNK7vq2jluR4zm/U6hQ7
DEa1NQnRivsLILrZtS75abSMms4QZXzZOFlFItJy2u6S2LFxJ23z7df9LpaCV7e7L/9d3xq+ZqnA
CKFfxfAuVgDN/kUFji8iwavDniixeF8vvasNc4sKZnLzkES/uDV55f8VJneUC2g4ylDVlMem0G8h
qaI/pLkHliwbyly6S/7dVriMhJMR+NC5snQFCkp4DiQR4t48FFUlAJaIuQDZC0vsJv4NgoYQZ7Nm
zhD4rOaB3QTNL6yt79FY+UKGwh0WskLh/O0bO3fSOm6Y405QpG06aLiDbd4u01um0WdzUc0lWpkF
3GaoO5J1RwxdT1ZcYmTtcdY373YRmpiL5fk5UkRzqUCMS8BHWllrJVC3WkmExMVy8UbO5/EaAGi3
TDMVZqUzYTdNeS/uSvW5R15zREJAPjuonTt4oEtzmGq7ein9Ag3xaJ/v1HnxO07ewqCR3Zap22tF
Der6UcPwAS4x1aTG1+NJk6Sm5C/UGCGeOPsRfjOadnguPUDYprupp/+5hSTcRoYv1ylWsYk/ZkH1
U8yaEzik04uoUbhIS45ndTQysc1y/RiF0Tnfka0Y0AuMrA0sEcoGG4HnFmSdQfEEbTOL7bkC58QL
TgZKgqXM3Gg2H8siLqwX4whYKLjSnavla3oydQHEA5Xyc7MUcBOCotvu/kicJtDruMzHBf6cXQ8k
dVx9QzbIq8cdKXNEXy0H2Qb2CsQQ3f3tRfR8dQ0HNPw6IYYEHwa3wHNwVSYLKawd3TTsPLZxdbMb
1DbQ6GYyjlpJ7g3fLKblfcQQEH51w9P4lYBlx0Cb1BrGQS6ZDgaxhao7BxWFkjJXWfj/PvcDtCN8
imA5nEqWQVEhgrmKnSmCo2aM6EtVhKHRwOtlFxcoXHGoU8Kh7kS19x+DA9l5Y9AdIeIZYNEiESzo
v89Z4F02eKrcgLdYDk6P+kqRhxrxhF4s2n81WLp1DMMhAOmoO+0pRl11f90ELbCiS1NBiX1lZeWa
vhpVX+0R7cvDcRtmpm0PwzTj6EEZqJW/23WhLIXGBuKN4oc/zjBpj39iSvEfhkIYu2lGgB02bTIG
3+vianzMPmA2L3Ol89ycvExbobQPwn8undT6WDLGO6kmG5USiwnHSLRe6MdTORPnEZzdr0qvW5Cg
mHWTK0h1iLEUw1Q5PNX5EXrYIAHJQ8vvxDV5F8gxwdpr+bTbChFNPReqi/qx8FHtWX1sigV9RMUb
/LFoMhQ5UzHxtqxSXun9VEmmTbFh5QD4DNdWpESn2nBkxwppZkHFAyzcYbJcmY9QYwX/MCwhvxPS
3+kxMokdO8HaGd7j+Dq7XTaQgzyg5tMwky6iSaALhMWpmrSKi8jOr/ZptlQFWtm9vm7414n2D+oa
24Kh/+Hk814+rUJ3jkJ6eDslOJCFO+Rsm/N79j1AxhQ07WC6dxSbYu3L9HhnP7QTI9ffR3V25tOj
dtOFL84jCZVGqcPymCe05azfCxvP5pTqc9P2Xtvo/xlSEGqoiEly2eIgzk+THnr0OBaxb2BnqjPN
OrkNvt6nbVfmeS5WpX9B411QP+zejxvM24PQqX0d8L8npY/5cSvLJgxz0qRG97bLcq3GDXom7pfe
dB4xvfaz9F9P33j4BjhG6WlyHSPl3P80/iPRLXa6bukbJHsRKf9lDxM16YOMUhLHVzWM3Lg5KDZ4
X5ikwdny83XjDjTW6Pa2AcfMJVTTRYWtuJ6/x0nIwVqSEgsYRn5iYyD0UxgUDOQnbaFjdolVvQdc
KjGkE26EzGATw7OtUPUeNtbfcGSvmanroEjaBOGuj9x6iAKyYjdvCgzItBb1YOXD89/ZYuZJWFCF
jMgqN+4t2aMU3n+6/bdutDv1XV4Ld+IGOK/mx9mC5PP5E847Sm7bbW7gLYUIPT4bxi54Qk3CGUCv
2N+t1/YHCD/cdtE1JnDaQnFlii9utDhiJZSxloNuShxT8svXRUg1xlSHfZydhzAg9WnNokkjOjdu
fCbo80+c2+TmV2l3CIGK7E0Qb+SUWh2zbuM3qBAt6c8MT2MxxFUaS98Ht+Y+p8NcB1NR9OuGsvce
WxuT9554TGJ9N00hAF25uJqAq9HXcmVt3GwHEWKok2BLNr4q7FH51FNG2elVzzKY+GfDp/nnnw3w
dD8q0g4e9mA/JV44fR6JRqdWsMQ6vvdeL0FLAgP23QMx8ZWNQewd4L2GY2FyAlS8tP8g0wXhHlv7
xtGF1kvKCwSy/q3nQucWhq6C8VIKK5bu5s4A9b3ld95EBHsZC4Ljxm1EGzHtd5L+md7/BDMzh8dB
+dSW92C9NeylPqrsyDIBIKkuAq2i8w6tAFfjoXc+n+cngkZpEFtbjHQzn3I3K07F4XdqikCBjq9Y
tcMY7A3AMs0PtLgayRo8aOZ5ixgPckVm+xFFDEEhybrGbso3fAx97MCn/CdNVqwqfGXh+AHW5KH6
AngQHRoVeT0AtjEePJ83gmRfqzItejetmeRz8kwqjNSsIlOPwAv9HHkVqQNqDOOu1iKBPXRyP3QI
wRVMmV564Eb0fddCDfsie+zMvyNUfCnv1oc1RlHNu/Ep2QaDXFOIracSHs9YQ0Vj38rCkSfh7I4G
TZeMbdHGJfAYWx+ITav31NIMSCU9c/ZilC5KYdNk0RJ2B8/4u/I1w8lOy86Eg7SHsgrAW9OZnzrG
8QRHr03idu52Th+jHKLA7JzTdDgT+NsirNCBBSrXP4XDiuaL9RHx4enmBUDZISdj3qn2IBYgXdSc
D4Gsaqty4Uxvmis7gzN9/aGknH9/xt+AW9jiHFIPV5nDtYwSF3R+Ox5xzTvwyI9BdQs3pmpmEbwD
GzZl9XdOIzTx9q6NxRsrf2F8KRP6MaLCCAju4BSbt58SgCQjyftZZTREzgbKyQBAU45SDvV6QP0Y
drhcfIFcNhJtsxb8h4tUtD6sj6kV6k2vjpJY/ad2fT4QqlH6dFGNRcsQFuEk1pdgxO51++bj8rK6
mFYSxnl5aCxy+iF1o0V+c3PDIptIWSoDz8dZAA7pwxtZ+yPw+ZPCnTYcQYcq+aEW+xJ+5S0wmEV2
PlFULWgExA5fiyo8z9pUqO+cpB/XcXumupK3SLnufliO3JxpZN+L97xwxPfZVHIxx8Jwr3pehZ4K
WB82TJkiPexdVynNH7MlyxjGkqPm7DT5bC3hA1Aik4sUKtzu5zlihEUHD2ObQ3B85tiv7eNBTHp4
FLwdsW/gMol41uirGuHJIyR3zQp9PWe8nbgw7xjtsRJKpCGnhxWe5kwHkK2ZTUhyvcm/C/6SyeLc
5v5HAVASiLexPvgD80dPVaqk7xdS2YzGvo5MhHnzESWF/VtOTYyftu1Ht0GNc8816/TPuh4hNFnS
xJrW3c1xk2WoC/9z2Mv6YMm60wQ+DASuWzltTtjGVz77xyrV0am0h5qd87edwLYgZUXM0HXRVc7G
RzbwVc1O5V25CKTRLt0YvDveV53AP6QepBAxP4urbsfefzNT3ssfwVOlc1iAM01FO7lZUcgrHWyp
y51ioe/f62NUa3IO+1oa5SFAkxgDLP1EAVcZ7h0MpG5hk0nklhV6zt4xKvH4fHaRHYvLRlXebzhy
NSeejvzzFZlWF27pDQ+w42ffbcOGOYBjMFdigJ4DuxKDFOHpJHtJGYKgZLKakdQsE/lZIs6bbC01
SBNRXJXyjY0y9AVTPwv8RQl4+b4KyvT8HcvPdTRcdMsIQ422KXINc2cr879GSYZceZ1Phz60uvDJ
qw+MeAfUUDh5GYXP/fZyUELWdAbEhoLmk0h28lB+czTp8bFck88UVEDNK8s9aN6fLl82cjzjKwQU
a8xUPfHYN3euSTwMBoKiq3xX0Mlj/TOt41gdXEBvYQRD2cjdJlI1kGFz9UYOr669WVf9J55whJBp
rHsYDE2VoCPILIn1vUs3UPrhL6FXNSLdVt9Z2TPwE4Qf1/eAWGbbY/waL3dKA+HVN5hEmqaeZNop
FYKV7SFUpWJWUs1BI7xaIEq+neQpk0tFFSMR01vJiIGPQC0mpaZ328SxfW/ah/ow5BGwgzjEL7od
ks+YPBhAZSEd6U7NylBV/gmcWYVm++SYbw7O039qI3kfL6sagz2cKlFA88UimoxLp3qPkhfMwr/D
KkUghfdFJLsTvoA6yENOwjIKDi8Qsj7kVvDmNEstMQXtvoYL9SNl4bLfmqMMvo5V6JHDPh/i/W4D
ByVgA+T9O/IMkze41nUlRKpdhniLcKiMQQkRAWyagyZ8j0O/MJJ5Wsj+UAWy7fi9MHRjSUl9YwzS
gB609sK5E0cSZAmrTqxH8f5whvouxEDJo+ToFm82Kc9MU32rJkR3Y6qdjlJrx5l4Qn/Z2jEjFbxV
8iXSOaT5s9mKKBA6QUEU5gMrc7TazxMHLfdOgeWxMQM4N1Dr1t+dPyynyBR9+O1futf78KRJWr3c
rG8s6QcmyNMoKJo2wxZdyFWd+ubbXYwDTuwDJEY/wkTxpTvGPlpIDAXlDadn0pcV+O1XW4H1B4X5
7axVmmBlvmxk3iZQ59icXx2h8pv9z9JMidBlRdnUOQ/EKlU3Foy5mk+wH3yF+Upk7xCnKlv4q8Li
1Kd3KEsFRleWXIUI1YIfhePoEFjQwW+ccRfHtNcMicJwpwyGUNV5eoeBS7dINUmCvgHohZngmqTI
vM0hATCrD+fOu2qbDboHgmk2AmcIOt7tsfaBMtSfg+09xLsQ5Fgfmlg7wxhW1vWSALaIZ399uWe5
RxruJ89JibH/3zy5vZjiY9hewNcTOqPDmM8n0knM4SSxH7IxucEETHLNKT/29f2yray4iFlCWb6C
Sb226zy6tvW7cssbiNx0WgUFywKOShGlXtnCOEqg+M2IqLIIc/jHW1D15fFAAt0OvpcrHjDr51HD
V+X9EfiGyYYKdSq92ijwf15JJ0+RsEe3j5+jSc+u5Ofd8Ky2LO+sLoTMbGvE0sz1wrYtrbDH0qzK
U6p1YUt+XSIy3tBL5JGvI+HXbgtp502vCm2gpeay3aURcSU3gaEmBJx5CZY1WEkqDwU75J8Jx/wk
RZKT57UyihZEDWNC/1uvIy/q3NvkNBKdR+87BnHselx7iyOUXy8PBJ/+W8zNwCHuGPLw17c5ZBnG
kdtoOtvQuNJkM4MeT2NMu+avo+AFynCugod2x0N3YhcZy8/7nKySyI//OVlFL2sRD7H1YMri+1Nn
NUsbN6Q44xLqNw6JXFqsoI8/91XH9UzAlVJQ+QSIGYg3xUQMEMxRB7MSzPicPU8ICbZ1zD2get2c
ayU35/CWHEnfrBtrXUgww+IDHlZ/lKw+XhsYL1VAaJCIk4oO0m5gKRkDVcm938ec2K07NVnzJ2qY
FyGWWA6qWLx4NlFQ2AhPzN5c5O6aUjd3pAoqRsYCWd4eJKw8VgKh2+grroU/hu3FDGT8lQYEGjNk
IxC/ca9v+1DNy+m6rw86jSnJ+4jg0B/JJhsfPnkrW4WMLJkgqOTYVGGM81wqgHc27krMEsmbNiSI
uekQyZ17sAazc+bxKZkp6GAyIjJ3gLJ8SvHyDknpTN9VzNFol+j7+jw8QuuMUh/R9UM1x0xpREwb
cxp+RWogEFTezPRzZzXgoWS532voNwBWxfTfVl9eB8QOY2gGBWCf70ytylbSVWL3s5QeK+GwykAL
RkSB/Agi+NwkuG1MI7XzAcUH1i2apBh06J7apfldJDt5vsYQp2RSNFbEO2MUtSwaZy1AaPU+exA7
wG/9Ifj8frAvkBpZrAVeuIubXT+qrJBnHZ4M93y52URP+8W6Cn36UtJNBWs+LbeYvQpvu3amEIhe
br2O/51sC3EcFFO16K/yPFPgARfgGFmNAzGjYfIQVW6Wi5IzaTnE14B70U9qnF2NA3F0cArCe9ud
wyo3RuiirNiIPkN/BvW7/LXQudvXkVpz0IDKbQrJKbv5TLBNCWxAHjgYSnx9LkR6KzKwKVDMHAse
/TijUr93CCOxKsUMoTz+A0pQu+IHozptHQUjl+CaQ+Cn4uOCm9Zal3UwgseXwCzI50O9HJsDBCzM
0duQb2SD4oibCxh87ufyBPHLw6pB1rHKDWjRvawNxDRyMZsOaK0L37Ak29PIkQe1hbkR+Rp9QZY8
HqBdTahETE7LNxM1BC8ZgeARYeezWLJGoMq4DFZxY6swR14TPk60R4g04DLbEprfpwlQeDyPYZJz
0VVIAyfSYEZ7Fd01AP3ofxPXnyeQMVaQfPWnKbXeybY2W5aTObm0LdnH5tyMRw0tuZA+O8a89qRg
zLz9nizYZxeHw94lowSocJl+Jb9Zb8WKoeS5qBX3VhKG0jD/gzdflmN82nE2TJIHTBghhoUuYl9e
wgD7LAK/IglGwPa1IGMI3IVqsJao4ujC4V3gnBbPadpdu/eMjKY91N/LDBdYypzhx3DdzyTcOsQ8
GjPhBsj8+SsMh3W0GBIuOnqSi+tnkgaFXtUy8WKNf0PHMtntsbL/WXVu7lIeBqC/nbMnuZp8+/P8
UxaX3czUiEvUCVp4SCo26u597DbjmTcJVfBrI7mrwkybbcsPYa4ITik097h5xVDibilmBHnJN00L
X2K5kNTzDCnhKkZvqNHvLJTMILcDtoRLsJQjItBS9E9YObql2GJ3D8OSlaFW2MPl3nJY7tokOrjJ
T+gbZqFWUlSNleUwSwKrsdUHQn1VnB+w42xl+aaFwOzCVxVSMCbG76NQ4j3LRXuG4AAT2go1+L4i
J/AoPxTic1UtFr2UERY8xwJ8uglz4lpYU+BQzvdEd2BXBeNkr+BnHA00qmonKDv/UAU+9lNF1E3u
5mdLCCYIXtioyEJjhWBMUudAvWtdtzCZG7krsSCJexli6yYIl77te43P7xk2Baj+WFXsJzxKs5/Q
OkPPfmPBa9Rvx88OcXd8rKY+/fZE1ePNMl75h1VxDPsRtnVrjVgdjYv7ws/wAb/dD5bOiz4m1E82
vpge1kHeMyjzNFaumo68O8FjBOYbJ9u++EVgW9XLgAoAp68o5FFKNiMRFMIg/7iCyk1x/ekZmYsI
BeYip5LUyvAaujFvwWzCFbvfBaDr1jJTALSOWoGOILkXihOuoBt1RArhCB1Y9OT96IAbj//UPC4h
qRa+SGb/uH/TvLlKfDWxDDhDgitxagh/crL0zru4LHChEKXdYVlYXmCRqVjBWCWwJ8mPRwqwT5P2
/Kv7cSTwxQxdeNa4CqhZFewpa+REUywwD9l2vIRzU31KMvDoSCLgnYBIgeKm7TFgqfE1g2h5mCv9
4ukHEsrmzBtgDJKVR3SktlQvlOtUtSg975b32t8mqtMTgkuxWLV5kq2xX/MheujfXssWCgHYu1su
1JBH605YLNAAB43/3ATRJPLnF149ZZblyFwr5+0TY0DHAKt4O0fWifhFnJeSFBpZmSMNcvmpPPZu
Mu68nxmvT6QyqTotW8Sdv/08x++Svpc2GdJaZ4smteRdBBL3nXEFewhdwbumf3Mkta9J79D49ISZ
ZIBFwzwPggCRv481LWlPkoJdKZ/ngs569XHqOGkg0ArnxgYMYchXfaqomdQyp6LgYLAKM0Wtxn1m
imEp7dFQx2uYBaRbICjX2EUe3qeAN69P3olkJ1iN1LViI7uEtIeQ1rpqAwzBdQvhvVUI3bAMmWCJ
Prrt9V/c+McmmZQZM+G0hB3IucYU1G3T0yfLOu+jAP9mYABYb+cTtTNBVbg86u9ch9LfCyfNiHd2
m7zxiA/8FW003ZzY0teErThDf2JUavtwB3gS9tjW7xncPf3Qz8IMCmmtCa9Qn97imsaF9gK56aB5
6HzpQDoxBsnC5hyOIOwwUlxUllXwM0k/bsPM6PBfM4kg8Zn+9gl6H7bciJ04az2wpxSphKAyoCEJ
zgcjFXizJUKX13DxaJ74uXf3pNm3343gwYT23lLBl2bMV6RUF/FGhRYRzg90hL4Q5DauoaQB8oLj
mrrOhfmzzpAoKKX5VuBB1esQWjdHfxZ7em5+vteSo4fIa3eq5KCd8JDY+hu+8Z7Rivk7Q244LKuP
NIJo0fbF5dGwU6O5e9uVl5UKl8qp1dmS0V0KQDNVRQ1oInn+RSBp71U2X9y9t3rqSYrU2YBTuThR
HKI7otO7W2YdyG9p1QrjEmH02TWfIVzUSgG1JyRTXmzC8psce5bzTl3hyXB0rk/GctxPvZ0pgwq9
QCbrxnP881a8P34Sy6M6sYhPDyfmb8aWQH/SGZ7k1zX8D56ztX1yoXmwNsizbqC12nk/hTMV6nbu
IDTrPhcgI2pws3/sLlNms4kqo5zHN9L+fKk8JnQYWBOZ9XtzWcDxcPYI0+t/zJRdw/Ljga9T9O/J
+gOd5vPI8eNWbB9MDOYOLJI5doJeWg3SYGqTqrmFaKPXRodiPI22U4I+QMHVD3GpzwZAz2Vd+kio
Wwl+LCir9SyuqrWTYHeIUEv//V5YI+9gseADU/wBZ/jqbAhnIQsyGZA6xVJNW3WFttoY5pG7a4LN
VW1pHObGF9EVJ4f3cHSw1SWVMXk6h/uJsRzYsMJGUPqk7+HOJvuCD4GuxiYBV5SjUT2yX3fCvYeX
InX4gfoHx3V2JmR/RP3Ep8hd0C7tuYfmq92l0huDHt18/Egv7AtXsjVTAJpBcLVstqRuXQ+8Z6JF
4HeDxoGiZHUzR8K+S1g+kXbxp3qWcRoRaldUQOfIq6nAQrRt5IkC+78MOu8pq/Q8YSis/eUlkg5O
HL97tsufJqPd6QCsEm+99ghafu8ZB4sJW2aieJ/lCnOpM2R2Z8a5I4U+//yv1A2A4BJ5uC5MRRIg
w8IC1YQOjN726FJqqXlfmKIxleUmeCuD9EbnIxGsSGJhUwmfmICYDZ4xCl1/SMrRDyH70AfkeOJF
GW/rYCTfeKEu3U00tTH9bYWmUgY3WnCh7zxrcilkOkrQbiJkxBTQlC7tc7rIMRnu2s8DNoSZpH8O
42fY3UY0eZNASSuIcvz6WZSe5gu0mV5atbHgcw3kvAhALLtSPLayX2A7Q8WYNlLRDRcHDd/k7hPq
LcmEEMqL/hF+nt/KOaubum4SbHsxWnUikJ6gIXJph5cDd5Dmhaks5m40ubo2XaDOmpc5Gqnw6fmv
IYUcctA9sIurL+lazz0wn3QRRTS4PLXjmMWV0tkCVnBFck9VzR5xbHT4UxReysYvJGdO2xXGKZhN
JlJGT35aImWldCd1Uw4OcsCMetw43b8UBrfOfqG/8GLoL/4aGc26yImZ5KCSSh6YmoQVXHJvKPZL
PhxCmKxSV8a7vwKWuwQjce84RK9rWyrvlfFSdcIaTm0GnSm1l7ILB4ZGSmj7B8vdxORD+UuckNK6
ygHt5W1xADzwOzXa16rqFFxHr7f2hKkGwlGVGtuF4aZ3qNZXg1Gdfc7j0Lgmi4o/KLPv+EozH4GY
3XLvglHmxiXkbiU29JWHpRBNdWk7Hq4bZ24gV/hmttg1kkCyTNE9SHLIAZiuyk9WCMvuPwbWwG4c
1R5EZWaKQXMqvYDJKkcaOS2/LiYXJOl2PXK0+8Eqa4ESyR0bSSaWCMUm7SJ8dRHBtPtPIC5sjNcI
UmeS7JsK3JdSp8jk1K46o2r+5+yBCy0ppWHkC6smFKDCvwNVTFWmvJQQBFgXxvE8UXNj5KiU+VoT
Oprb7OjZ/6+cJApixwp+TMwd9mIbdjMDpOGlAVHjeUiFvV92EPOie9KIcDMBk4hxXlsa5JvvEQDE
HOJ2sJh4mlcRuuj9GB27+YxoDRdcTIvYeZKhrr9M8Ov47oLHG6Mz5hRYVWl/egqVke6ZdwDNEbJu
3g5N+aetZw4DLRqKKf/AigVMmVgg8RKhKsknrj3xLzHjadY6uMnIrg41u0LKh9zf7222WaItILQj
fnuMnG6IcSVH59EHGNZxo5WpJKHeFwD8HsODSIx8r/nrRIOxZn2cRgpxGpjyttQRJ7m9s+n32To7
Nas91wmEMI2xW9w1r6goI/etgUNRP5xkAiIimDZqlOPvKMJJ/tyZ4gFrlBa/RBtUInWOSiE/AMKj
m5ffl+OF/9GsNeVWmGK9IUN1jB3F6dYRwbHP8+/R1WaAsOusM4JIcyJ13d3B6yjWR3zovqu9lpog
O57EehWNw2J/1t+dzncdqlMwNoxjPdTDlIKsxX2wjAN0j5foIkyXKZBU/M7VypbQDwrG9Wat4HRn
Fn1NTOFcHxVcTHXImBaHYYU/lImVXDG7W0mYxKZcMr/KdBf2KX2PstQvaZ7FchhA50fIaxRsqUG9
a+LoACaJvtuNniqKR38UKerYwXzcU8fTKabFCCgh+7DwYiVeYsG0C9e8q3zt43V5pHb5Skfsa+Mv
YMsMNBc3gyJWaW6oe7QaSRzPuuoXLeVxpJlweNordDd8nc9nVYINL3L80JZVfbOh5gjdZTLMOgLS
4zjqWr5FQWI6f42HdpTja18lx9uPCu9SZ7rUzGgvtULgbolNXKZby3YX3w5co4mkBG43uDj15jTk
SipHJHu852awgoxOrr5a/0QVPfUnf8NmD4s9uhQPLte2BsGuP/KPD173fU5ShlonVKM6Y5Q1K4gb
TETrSY4EZghrMRbjb3vSZ903UmledEOm1fIMnDDy+yr0QAzfUjohlDBqlrzND9OoWMNF8iuE8YhM
Dea7W+9c8iJWbGbkNjEMdzgE3pQxRuTXGGanaxi6JifwVwFeodva+xL0hp4uRfaMjJg2Ja85S1g1
RoD3+ZzdI8/C+aNcN3/idIuCvAszo0Udl0R4R2fgt02ROK7oMTg++tildPVEhKllCPFIKNA21pKI
WT8M/89j5/6dBA6xUnWvaRJQtAulmqiRHHu8678Y5bxlyGuqXfLDDaNhJHFOBISSY/tKj+FkLar3
UDcwh0QDGjLQOfogBipd8IXQGt3+eTB3nn6EpZHMVo9lT18BrXw7pMK+JQGaeFei7s3t+pz9bsqt
HzDe7ILhc21NFgQvjHm9qMid2J7fv2u0mCrJcJy9E16JQgXwLzrTP3TWU4+iqgLB+YyXnvfzzxOV
GgZTSXZFeIgtF07XjiV747vDt6eEuhGp0jWgEwdLVYiLyOAm/E62qDX/7nPws0/0Ie7Md3gcUaYA
d7LR5lVvgWR8uesjbumiY5dRqzT6XcTHPLqP7TFFtUfmdK5z0S43eLZJWMmwtcbxF21BFvMbRZZQ
Y+91nYMxJl7MQGUEC/X2z5QadGQzmsuWmmLWX1GErNlNosn85W3bVVFuO7ptoCokjn2uYZb+WoUu
wxNkuRAzLanKgljRWU3Lv5Nl5GD/wU6fhFsWWdHVK0FbOCOfP3RBUG9kPzfDWNmD1WFnMGGDDd1h
KNKdY6sj+rwTWY6mVdxGOgJnEQsyIR+bCr8S4dKVzPcaULyAbOdF0tHo56iFbrqku9YQe6JpFrL/
an7vo5B8h1BNYra/G9L/1R6gbzu5AzwUrZ/6JMnPrJJhKj4bA9te4hVh8AU1Hc/RC3W9lOowuk5M
J2G172t4O7mBIhxvUa+hYO6fN0KW4p51FneDejteT0cVATicIyayYyxQnf6F1Lh08qasO7hzA+Sw
eHWCoORj2eoGdYuLdUod7J8+3sxEPjIOxBYLLF86IdngG4DzfohtVB+w+ZUvxrehLV1QgKvwFXLZ
NWcYf3zPpWfeHIYb2/LmwV6BuSQUDHVZDLGu+PWxg2aWw4EgPINVgGKReou64/qzm3DzMEBa7Qs9
74dGZle8L7zEIFvuQWQdcYQvunRpVWPPMN1dmSBbj/RtW+DRfAZG66872dCG1D3aPPIurJ6l9CoX
bAkXHRbfunJ0gCH8xhlWfzXmKwT3ds27YYYC90MQ6/nafqOGZsCwt18sYxMnML6jLNOGYEZQT27v
jdqcnlZa26+pPbdt6HtzSznha2SMOnYT00S5E164fMrv7Br3eq3GNo5HFKb2FlrW9eA9WkIwDoS3
L8u6DHfH3zwpp8Gar6PHINipIRvCqx/4gIfWQwLCt05Me3nwAVougKW9c/lLv1Vr9rZPeOmK9ftB
9Q4RsQLcmAO+bHnZbmmPrN8FOTr2KI19H2NEe7sG7S9jNMpVPMEEOIcMcL5ayEB+qHZ+0FW5RBa+
83jLXE6Lkpv/owNuWC1GlzXOjqnS88sSBg0QNMnQc6U6oUXHH/W0sVdDX0244YVVCRfIOhj2OV+o
hV8Qh+Jgu/Ba0/IlqqEhydnlCCPKmu6fihbvnGll29GBJDy7QVRN0i5+FDC0NhxuZgTmJFyvWw4I
NnRFRhfTPOYeytW9l/G74LmN86qJR6y/yLm5YbuJoiS6+uw+qVaN8oJXo+Q3HqoBwTKQ/p/9oHuF
5BRayUe2uN3q0a0EZudgfGK6OChuDNs7fs+IQUkSKZIX5OJcdOmwUQMjx6YwDRStIeTsxW6rkxmD
adzUkBYg1KscGgniVGtpZb4PMFidmkruzLPDSkcnAUuQ2sTvH4+45ozc4wyCjTUsdKlntEJumic2
lXH4NXAHBe/PhqvHFSniiJWOn8i1Ffoo/HQp623AQHNSLiSP6q5ulg4y2eb1D6YbA8xn7hRw+0Z2
nv2If7P6ItTZKi/pBMFQUQufRtW8mTG7wm/G9ijh/8UiGuEcXmzw4ybin3JaBREgh3ODiyPeFDMq
J+7Gp79V/2jrAquTn5yPF53xRX0gDC/SN8xdWTU5bbWVD4nr070+srLubQrbfUf2I7GUYKct0HsR
+hLtbUATau/2W4gZXB5BgCeQUIf/Mp7mRT1Dm+UhD+TNz4dqh0kn7pgxkkmDKpoLbDFtvlAk0r9+
lBXR3p8v1Xk4MwY+y3UuUPu2FmR61B9r18J/R+TZ+VnKq5CLwT8JW4jUrNJIK8wtZ8P8l6crHjzB
ZPFjY6Pvv1EJ1AEItNy3ziA5FiDnEy7KZaPEJXsWKirCwTFl9bWDEMHIqElVmqMfFbfy++cQwKpu
chzGZhi32d0B3y9sI+ouejM9F4EJkxOx+d930I01l/VipxlNU1zLTIFUF2XbFFYP7ILzCUzFufta
p7nmzuypGumqdot7H8G86UKBO3jFRZ3jRZf/eLjSA3orWKIlddXXesmEnZ6vRDEgakdy47ZEuvdK
6trD5Y0YP6nSf8OzbApAAaBbV8rJWcWlrOTHnTvL5RyOUX3luagcLFSayfuMQk8VgSGf1nWokBPd
lk+Oob1wOm3G++mwEalUXEG3AmgewSi1NcBp1lDbjO+llePD7tbj47PhG9iysLu/9fyo8t8VI3Zv
2qzH+NHZejj2jpJA5gRHwzXNN3mzV93gmGmxHprc36+d7iZSOFzcMKBZ6MYtAFOj7jxx/evWXlRp
uGah13otkKUI62duVpaLxvHfK0gW3PBPdHuPNmhwyXQhjCEQTJfokFpK02OTLlZJ1JYAo45LV1jc
MXBFN0hnR2htkWpHLWKsd0qM8xKbfxHxVAofZX8ikOD9tb/g2drkQQAD3quK7OFVeNsrC6TP2eLD
RD30CU17thMcb7QcrV3vmdDuZqVZjNfjnCLhmhMkv1lDNgJ5vSCoQasJiT2l5xpu1DSPd65TQm2B
4L90+5f9TQkeIqfkpQ7v0Xe7JJAQ3gjGfN/Vc8vgp6+U2m2JpFp7rNfyIscvWNRGFEvQwxoMx5yh
lI8v+pZHBAVDUxYg54EbFcxvaed4ELiAMnfRY/FnSazEwx2sSSacooSml86Fu87dvBJSjy1EfuNS
LqAPOpQIfrmmg4ctxovSfRrhXoXswLMUoj+rZOeBu69KzpcUYXREcHuZarU9NjOKx/H3nYPECFLl
ygEMZ0o7t/wJKTQ9XdFl3HGe3cxWYKWyz4wwwb0FHiFzkeR4nXdkriQH7iE80H/wH4N7c97VtxQ+
KxhN71sunVwYAMvkBpAVGTs9Ac2ZIuhhVd6KAn5shu1VYfRWxDP4NxmXF/gpzcdo5y0T2N4w/5RE
eOWCmzKdQuHBVdq252Zpz6a2QAk7ZjMn4T2e02cD7xssbF4eCKw5Sw2qVWsPZePMTU1f3cJBz90M
zWBGRQ2a3xp4aRD6aK4cIbD7Csqw80rN8QJIYu3rxjRgUriwbeS/lPOqO0cEkJoEQQojneOOx/6Z
+GISWTlDuAelUxbT7lQUe8oVuGmgx0gw+yXG7Hxx9i9nD4tb1UzjWsCrTBMltM4mqxs5V9t2Ice8
+TVLml8bOcTK3VDuxnGWbKYNT7OgBGsZpUeTomXbvB5k0T5xwuCCpfQ3I1qzpTsUKTjYD/hvgrkY
Weye/h+H9jylYbi8McE40wGR6qbU71xeGFr9s1Gtsubf9HeltSz4qhcfoPibYvz/pMabyP0CsJW0
JqOGeZP1ZEKce+O9rQMNl8cS767A1GYNl+AiyPMk0d3ekSxSAYaXBPvqQf4VU9q4VDG6o3FdrAoZ
DU0L4X4jr2zbzBWW+ABUgG53qAsvYA0vmn7Zmr1qFzMz0dK5Sl7Oh+rP9VSF2OadT8EfAjUSGqTi
qdT/mFHbsXmsLPnsgZ2llypCjuzaHmFcXoFGvDxWaGiob0HfB69DTLHcmHjRO+nC8Wp8QgeDYhyy
KY43xOG613HI4jBW8D4T/wQQCMF9ly11V7GSUg7XQROojv6mkIZtB3BODzgXD8n90JKN99YsMtks
uBQ4RM5AGN1KSya7S7ei1IO9mRLzveweNP+cq5iddYuh9oKEl2D81AGGp7ttYgoxkaeV6TQX4VQl
qakcCqrAUSFPAPqeEU03rYhZcTbJE9YrRuiXGxrgH5dukPNPivg4jJLjpMZ7cO1+ezlMMuLzAxgs
bThHC4DIjqTbpgfejZ9rJu2mD2z+aVcfufoDqoilFqYQ7eTJBGggn/NgsTh3BMW1YUd3KNdjkBSi
f+A+ebTRbsLpyNjqfTzJckilUa7iQkixrJJ2kxHWL0+j8SGMJflCdjg+hmeND+MFSjk/wpQy86TP
uDdAAWZbuNggtdhCjxfmy6gtS0a/34dIgTMy0EObNZGZRJqg7CckUQAKvmje0meMdioqgPX8A9xM
B2Ro451bxVtYkcxyGa2Fou7gC2i8zrYO3r4aqRbqwhlZPdvOqJoAvhAZLbzH7nrHeHWmLVYhyhOy
DzG0uhzHl/WYPXdGGII90wSzzXoBW/sFz7CKRUClErI90g4mm5HeWT8IzNmQNWRAFXTisNawGIy9
sC1ZiQMg6bNsujktVMTpfztjiR8sR0yt8s6kF6UnKhg3tomfKaaAgsDRTkGcD04YYbfZ/oXzzwkx
MnVlk/OlBg0O8c4NcigPp6hpZw45wJIS5gVDFTy7Yrtykk/yf7mAPJkJkmspyH6z2EWKD3yfdYvw
jlZj1dDbaA/OGWyHwNhXkqGXfZqSm7gFgfnoM6y5rbIye0QdjHkXPWb+l9IiPcJa80nE/1/f0W7M
sEzD9ousblGBplx6pZDM12ceoMKy8XbefY4vWmD+i2KbCHxdmtEcp3v9lEy0knyOJcCn0xATW+YY
kwFlvt27B6lL6j9s9Y9oOrumx2X3h4igWsq/Di0vZt9nGVhs0vlHJrZPCg50dAuvsWjBnjSglKnS
gRrnqKKYwh8EFyAeMu0JmLh0YlHe9A6MQ3F1I4Dzt3COWRyDTHFk8Ocf4Bw2xkZfkMvj4EPZT01X
Gf7KnnPxBPgv5ft+hZUvQlR+ld6vL+BO7t7L824VJBxcXW4CgEMEvaCHfH1QC8q7d5a2ErIi2ORa
A5TutilZdrkVujPMCt+qJnFIefpx5y1W7a0gfgGNdSK0wclLnWpzxUcthZRzTV5O4j4i1X3WzCVW
vhfLwZmdtzFjYILTkTk5milvW/YY5dpoEP+OWl3P3r+aGHq2mYrlXS1ERPZN+Nv7DRKvt+/EjUhB
R/2kfTRVA0hpXOgAtxlMqgpiV4H90mjqZf8+zKCuV8E5fmWAp4piKHk5+jDNsIjMLs08ms1T2ld9
gFOMYdXQhJcZwHTBenJCNLAgvpW1G+5Q2vw7Ks+WeKJLWPu8ujUhHgxLSgrIY4ypj/5TVceHkbP8
TED9UNcwI/WZ0hRivalgRmp7UWL3ZvHPqHLOXPnFHs9Ik3eHNllNdK1VoI04bsM6ILQdmYRte0rz
52sN/gMVDGKzG9Z5pWjGN3uutph+fYqtrzZMbCdsYUaaQU/zPXlJojmSmkplM6nVRSoFtnRtFalr
om/yL1KZ+pS+edD5AuioLfVj7hUpw09THUdCSfgDIX5Jm59RqLTEnwFqdBYAT6rRyq1fI/ncTMGU
zvtX2yMhQSsz+SaS20OIPFhpr5caw6FCH8vE2WlCYIOhxgtFEarcjqtG7cqsvXGJVnCBC4ADLY4d
atRXYUTAr4DpicdJCiWLEVkiUt6MH/rclczgFA4Qpl33TDu3kjZd3BmImndy1xPj/bNmWzbrYR1R
ZKoTGQ0aXCaq7k0UVnQVPAT1a7oBX2ZipjulUSQ1FFXktja8n3uhaKa5diJE5KyQUq+kJ7w/SzKA
WfEUP0KqNsd38GQqz1S4oEo3fGsyxoFOxMsCNMvlL/3TkzQPf5EYHUwL63agI/M6qNreIJ3rV3QA
Ve4G1zp6LiEC0bs0qC1NmhBX3jyyis/YGu1DiyTWiBCguanAcXGRnujYVBvUvQPrNGInig/0LEYA
t1keXJCUHuUoDk10tZ2Y1yLbxpYiREet45SkBlzCCf2U+KqX0FCe2Ef23fpD8tz+pfvgNoNjQAjj
NXPCb/2PAchgLi8ZGAH+IzL12g5rt6Rva4L6tybfYoanIbSSZliUZU1/nEL67wmPSe7wB+iNxKL7
MdwHFFHBrDOsfisZc8n1srMqbNC2ts1qxGQnsAx9umlNlTEJ1LhmVJCFFBWG44TDl2CYfg8e42jO
PaeN2pCsWwszVWk7Gtle2lDHp/Sx7TIiYbPaJEYOBSZtyA5l/yj8vgWHLs1libuU6MVrR7r7k8E+
ovdTDn16k+LKclzxRM/JLfv6sL6XmtfOi/UqLYmi/o9X4qZNojLcrgPHCsDelRxJMluPRs6ajmZs
+eSQ3PppjVupKLhBiDIPe+SFwpJWA8lmPApxO/FmsQgDu/aNfPANQFiNS2Z69YoP/K6gwXkpdEyG
7VF5Y7GGI2DLy4T9DYnWJikxO23u8QpBYdWrIDIhPHNozOewLX/DW59/iv7ZC6xn1K4Xn3A8Fcue
1jVKoeef7vP4CfSOoLYifVQWMKqgENi0ItvckrbNQqfwEsom2RIMQEDaDvju/FtN/9UjO7CM/qj8
JJTXjfxUe9P9SCg4K+o1+wLZnjizCgZ+E5POc6Brpx3vfQmnCLxHZedSdU9CNqzBGvdUS03tQdRc
HG87c/rDq2T1bSldaNXlgiIVQSPHCnUo8ct72+as02xacyj2hv+BdfdJAfZm6e+Yf1OwZ70bQ1MH
6MY7Hzu9v4wtTelst3f5STGgDVGelSXGx15SYSYp2jqOrUxOa0QsHtGOFhOKeduC1Vs1OCFv21ad
moEIPlEzBQwWWMr9NyCjzOjoVo4MiCThtQd9ToS3RUJU5CU11sOHWexdSjzdVzoxeaKmb/oeDTtk
dODHGSB6EQl+7spq/00NBB+0ZSoZU9/cSUPgOqcwk7CKan++iJ3OjLJkEhsIyZCRqz+vYtlyr5Ai
qGaHlX8W1R0+bxqH/Ghie/L0K4eLzxU/s+VyIXQBDqKgFTJHlpZ/AeW5LW+91mSHCvwuuB8xm4oY
LCj75ToKM76FtbVhWcuFX+e5I0Ro0arpDlrWvTyRvIazZnwyFXxssgz+Q0J85uN/Hoahnzcj0PoL
aKJ6Mug36vlNy/BgyTA7UNJJ5H/dyVovR0Mwf3wz/xnyI8s5dgBnISq6+QnokgA1onifvqubO5Ch
oUU+Dc4Orndm7IioO5pl3KQ6HNq18OzuQSAUS/Px8qStg8xs0NnRUZZ8+1t6Zg4eoO9uGfKnEqzF
unkgBRbLl5ynHochcD3Gvij3MBI89xZaaXwEg9HQTkyP8jnObTtCTX/gdMasRBWJhUYLvvxRyM+H
ZeOmV19LvdJGj3gdpP3A5bnsMGDW0s3Zdyf4KM30vCh6IdXYVc3X5S7iTqIRQltiRNsbuiGOisd9
YW4MrCFgHVcgKxE7ecZOhxxhEXf4n8sIPnufBhtl29XvAfKlskiWiJ0dgi7ALFRaClxsSK9XAsXL
SQQu6Ek9CIHp6dYFXil3LRJmQwpInIyfbbMFGf5fSIcBEyzL9RntteTku7Aw0CBTIp+rlVchAbgS
7SVsBswrRduWRYctTv+3nh2t6zz2c/Io4/3blrOMM4SWkK8Gdk1QhV33Lm17CTQf2x9RamSDhs66
HRiW5OlrXCIJ68FYgkKC8QV3K+2vPxQlKXs5tKmISkRqGMeXQ+Uf6aMPN7zgCFlkrQZYB/QFdpby
W6wgxy97UnXn3nm7lzTIRfHPyl4CN9otN4eUMpCygbeYieGlmi3ZOx49+rzGp4TD/wwT9ngeV29j
lkDsVK2bbwa9gPc+XMXAFVXgTzWR4VZxnGYpDigZviqXaHfFOerWYs+uEKc/pJyypDl4YMIMJZp9
KboYWmIU9kePTaleRDADvvtqIK0/1nk3bt1+qZhy+mxRoyt9nGFwoBsWDVqL/n1u3giA2rdTHc0F
Lq48WBuQNR9O/XQnGLI8w5JukxmvjxCwVd2SP4Vbmk9nMTAYOTXWveaz5RjRb4gOUSNLhNtW7wQV
bmQpZ6wXk5C/c8N99LfuD0ptjwRw7BHeWTLTS53imtA2tEp/tDHpem022WNS3cQ57dBvBelu9WTS
CgEZjjUHxYtCitQY6OXYg5uWVGrrTkbU/w32ahm4hPJPKNvCw3UzTF1Gtxwsq58bL8SmUUIT4tsN
lY8Ip1YfRsYclBKuYTpOBZRn9rkoFKQ+4xuAMqiBzBR+S2EG0zFhW5cGrYrAhE7SQy15KA1UGnRq
ltvh+S3Elk5d/pCJ8ZZMHOQAmHVka9MrlDlEWdrMTP1+GhJYn1ZM6L+RwFsmv1+JWVDopkvFEagB
LvX6QNHXdsXct/RsBVyYlgsWAGACh43O03ZUapo7sI+Zdz/floanOo5tNgFJKAGEb8gvhWMmwPd0
Yx7bOtdjhrKFMLHnqehPEVSweXgYbdTrRclVBvxwx4pLW0LyTAT2OFAtkSSUtT4wRSHUsD9zhTkU
QZzNIKI7jx9tFh/7D9Uq+iqfTKWlB1+89D8NUbbK/ax31pY7U14QajfvhBp9dV3nDsdWGXO4eE/Y
TKAjPdYYOxx9zCauxE2U5uHrgl2uQwHR4QEW6DYKUtNGYr6Hg0EMOqj0cYYPB6ifrME0bihOIaxL
4g0yu68GkG6RA4SGqg8wi1Bp60u+2JPuMz66SSYJdAnKIcI3LzikHwCYKtuX1nYzg977gbbz8ZkF
Go2ULkDXEjWPlvU4d+hvvoYuNkobPkdv8Rce4bxYNyCto82PeJx99sNXeKaJ/315gVpS4EM0qexA
3ltGFSf8wh1D60Izkh9yF8CK1FVRr+3x3xG4zOFvIAHNX+IfRu2i2wim1flHWBhck4BYfXtYMt4b
VGOOLZl1ilYRAGrN6ScJXVAQbr4fWhFKEoCfoYPme5d8aTTBKHhYRGpEnYA7oePUioR8/IoS17UG
ci68+TFxzEuvtYTvtB2fnzCqpD66AN7KZDgrdyHhDTp6FQEhI1jDf5LoJPX9DaaratHJp1FT/efS
f+Buecry+9WSiDWNdamN5SOiSWKA6hkny2lW+Ww7xLYmsMcJsSMARbxcLo6Uj0THKNfJBzzcMWzH
hUFBb3z7ih89pSnlmeDbjR+OiQuzMVcXx6bh3tIYTtF360Re6K841h6dI0Tinb8TaxlYkpjRE5Nl
riFnT1iFWsfLrL7S4oL0fvIRTNOOKjMEf3KXtqMOYiCQu9mIMB8WC3ZMtwZAVWGMY/on7oIWL23J
iKRpYcQDRrcRPo/1kwA5TKGLlwFl9cjqzHyeQNqgxIIK0Cx1H80ZCgIq3Ay7o/ouqHyXTwSavjKd
f6734TwrClCxS/4oNav5cGGam0jx9kBTtIVqvst6BEGAqOHGwy/WV+72vAKFWyWQ6ADN7+HWCzo4
4GPmK7kPGriHnpn0IUx2ai0iyRph18hrSbN73ULU7lPicX4zW4yMQ5DJhZqJZhwaJVY9BCWaMQ+7
o2gKwuLF+nLoJbtt0oRWG5QVHhMMrIMO1ynnIajZzDsstqCg8ZExZGCQnX/EtnpB7ba5Rq+D4xo0
EL/A9r14GJGPjJhF+75PX4aWSdwHH9YrBhtvIG+xnMdzaUTsJ/Xv1xwAHvYZiTnYyfCA4CsrF9XV
6uOiWFhBcRor3Gd0YgjYiRdcypm1V+LGaUJPycailXWNt8jyp3bjTPp0b35yciBlIe7+4oVtkJe/
B9RPiwcdLxk2Enxyi1+Wx32i6ho2Sm4O5PbemzvAJUzB3ul8ss4ouNgkdZgLoFz2rtWtwXGlVPXA
nNsIHu2KVwE7EzRQ4a65nakAFbs/kJyhqhwI8cq3SfLx/Ym9yi9tozplZzvfK6nVNxs1Ni4dAxAN
k1VtAGSgO+HUlwJJoVVTqjVBgNd/uxtxXNuEmtV1gmXgLRPbbgrUcq2y4YHqHXttDf3CPLtKFB4r
+trHk3iqUuO0vweou5hh+asWwSIy/jC159XfzCfPeh2ketlULcyfEFqA+PYXUDZOkVYuYMIfY+xZ
UlXGuy6gS4+8aNbu81Bq20Wn3rppnkRcEU/N2T8/Bm/MzpZ0tvpIY95u1DadQc2JpU1QvMFE2zpa
/qShc1YjYH3LhOIIDCej/y7TBi2MbL8mS+oEpKZpBQAbc9+ncQl6BS2aTYzBBvk9b4SWQMxvrJzP
KuhuAoVz3vAh3gzTKFWNTylrYBkO0QPg5Tc1zSfDbbpoHiIxHBd7d03B8uz6c5OKjAna9e9uwkOH
wBnCTc5PMWlIX7hdQb+YOi/SCrNYDElOgViregSindto2pP1jVwPxf/r5drvqYV2LkhMV+Vc7WX1
hKZWDo/8PeE/miChE1wwmuFMYuGfwR5iz6PzNX+hBN888+EOAwVMtj/F2z4Eiw1vbFYTIMIHsfSe
oVbF2rLJCwh22aE0APDHFRFqOAgV9sinnvxPCTaBojOgHyCDrSBFTxr/LK6QFEQp3l5iEeg/9rg4
WGBMLvbJhDPmOTyLPz7MKAGCsFqbZnY4bAB70rD89OgNZDdTmSqZ0s4LyxDOCt74ITSfHyOUSp0G
cRSvzzZ/ttk5+ktIFOqMEfKz/yFr8sVzw8+NMO/46r69EusU3zdS1jAfM/RDPehH4nTAI/5Ga81b
4ARmeDqvc5bI9+jfOPmnbc/+OKVZruo3oSByuSZrOf0He8KZYPwtbMtfe4UOESldsJCCGWrAJJkC
EEd/IhEySbhj0+GQDOMIvZ7rqB4c7pzfWI+WaMpdOxvrcyalhLmvj/pZSTSozpbJJjFli1LnLVV/
Y2CeISr8EHYtQCv837TtJ1ovOQUJx6NBF3G+riWCpFyIArLUyMKJTYcEP8/mXW8SY/CSAMXuH27R
maQ2t6A4ktamsBDC5Xttk9MyX8zH2TAaCfp8Tt48cLNuXqWdlhRkNFgS7gegk0DlaXSUSt79aHFS
kOZqMoA6q5c1XUO0tNjNUuLWiTnA9gHRkXUSJHlPIK1uFuZ8h6GTHAVwL0gvak4ie8O2opq0ZMPF
kM8RCMsvEvvB95SXTeOqgcKCUwqFJGn32lxe9owSdAV0F4r21t7pnMyYULpjAO5VHL7KVMAKNnlI
e0HTcIkbMhUgTHtSJEzqsBapVJmJzGYCmwq4siWflSQcx8jwG0fXHr6pxrQvYmyzYUN/AzbR6SmG
WAtVxDzXXXP9Ex/IahLk1xoqtzJ2Zi83JgTALhFX9QDzcL5vD5SSxwBdQM8t6L7tdw/VWAd2vKHb
cotYVcSIdKpkbBzNz+MM4GeSMRH8eX3ZCzYQD3/6QTdWcrSmKJIZNuxmksrRJncBALYOTGIm/f/j
3MHJQgpUvvIsruQcB/Vvs33VnxiU7YFRYvcFdygxFim6iUeUqrEDU8Xx/yF4QEvAat8axfpY4vXF
5jCyc6OLOgqrJmt29M4qui1TFO3PfTnrmltDZm5WPSAi+CGx15krZLzNX9JWy817WkojtbLVv4Py
nSNyh2pbTVg7F5+Tem54F2M982e50kTC5TRe1lsCunW7RaY0r8r85zbMMyJi+y2zGZpAOyud64Em
32sUeXgvM01SHk2Ompxv9oAaRZPN2cINL3gyAP4LH0wMcAapHsmlr6/CaTh7RM2yt7e0duH6E3YE
VguarU5+DFE9SXBWHoFiCdJ8cHUR8esBeP8V7QdRWrmjl/FXm6MhY3nuMFwqPaLhvk96XHdH/7Oi
M8SSJ/Zonh+02cJ4BibIl3T6dX2GkN1lxcQ3rYN1fORAwrzqyDAuvNqReDY7NGXsp5UVrQ3Sjp5F
Mg0Z0wRmQiFdpdCGt2jB535zyRDZEwCG6TLgES2TyKFzcKaKcINuNLFPYwLMQ2zXopXICTxfLUnr
4XBrwryXPr0DChnxrTHmnC4sc/V76uGp2eu/qLh8xjW9U+fdFM+ce2nMghlMVIFFfJ47hempF/Fv
+yXQWA1WS4vAlYjOR1NnzAKmTfKH15EWMKYxoFtPf4AsqPIWRVGISrTfingaCDopJDTkzdy4NKkr
u3dpPeL+tsZs3EBj24ZUKYWIijQgnBUX/FgKwRetEsmAjccBa8/CBWbNLOShMy9VsdWXccIXitn4
kHQ74huaDAUy42oInBSb/mDnjS/4/gpfEhRMg220Y3twkcrS/qsxm1a0jv/h6ctXnOZOp2wG5u6q
euNc1eYklmtAHdrkykdVkHS2OyL3RlAdrCEAT6M6l3clQo0uL/CYoQh8hZpQrIJhhwYc6GJ5PYMK
cs/VGMIwM2YAQKiCD1BbyPypn/uYHXYHa0yuIS0eHuKo+Mk9YfOaSN40wLxnMrFiGChW2gifnAwT
13URUyTIxeeP0aFUs6emK4uGxCkNHqpLwq7RBvJtW4kJCjiTNi9+FzyW1xUH0UY4/uojp1RnM1QN
7rajc+Q9WXG2xDHdhDzRNGVU4crTcHr6PF92kyiJ7gm/OO6iK1hTb84aTGIColVPyk33HEa4LqNv
gxtHzpihk+AUICnSEUC2fIFnqnq4S8+Jq/4OWV5S+sqpzuFPPGtLtbetLtjYNhppZzxvzrWUELRu
NvpuNtNfTM62Ne5qiaDLezgloKOvgjn3+1jlPR2mXb2sfJjTF4AlbMfkcDWqaFi2f6bFn4Al/VQB
rHITYnQJY3Yk8P7dzNz8VgWrz+WKIHziRDqzbp+mFTo3+TOaMkGvov59O5SZ6/KjV4auh3P4p46D
BF3x/v1rf4iG7br6B+x69e3jFcnoP4PHHsoR4CGwXwnX3ueJXhn8Ek2dlr5kWIW7AZmsmGP4X4ra
8QpUxBZYKK7OptcjvIoAbo0a5EyXMpwEDPZ5bxBjP9VdZ59WYpDSCUrlGOzyZlzQI9wuHRPuVe1i
7N8ZHUQLBgOu0kC1SJo7pqKxx7vgSa3/6/3A2WCK1/0IHqkAQQ8as05xUqt5KGs8i4ZJJZiZtDCk
MI0kemRcC6fUuH1/chIx43NQuUFMJ7a85y5qxr0bOnbm7iW68wNwHwDtbQ+A7qYXVJnuMYmU7WgB
NscMlnoP9xPqMPzgFoBUX51/80c4OSfp2hCMTSeN342F//ItM/dE41Jy1DFMuv4MsVy3yjmzt5bp
Bab5pqnDn4lnNSEIHYC66Xmb6IgNXyAvCV5cRy0K4jJ8QBUVRhTX1jMCzx64/3SxHnDVB7lqCWu5
/XSbBcxEb2RXbq560f2spZgmRXkm1tGP3Jz4l2d95fJ2q7tDGiEAqz7j2giADpx//L54eCPwRC10
bcHmK4leBum7Z6owNZrt1M5/cgt3o6vig31qyA6dCkJyWlxhDsWLjwW1KN4ZBY2byfpawqNv1bgN
Bd3uc2NXR7YHvbb6gECvXi9lumdvVZ6DVF5hWd3KjAxIhif3FZ8ieu1OWTNoZy8LIbVb28LUu4rh
jci/moe47rpcrH56Wao2R2xc8xHP1MrYRKhTPByNJBTCjXHlMqAZohPhcpIi8rtqL5DEoQ92TRig
43/Saxi5VnXbj7/hprJEQg4v1SZiEvF8vsbl6gNABB70WBa187ERDTsOyi4e9i0mTPZCdHFUHQ6Z
O4Vzoe9ZLLXtK/UvZveYr7j37QOi1kKpiA0TqRt5TllqGou2JUm1RzKXiEy8tSYf4cb319BLwjJv
n62uDlpckCGNATx0w1udk6Bxxcy7mAvSfmGv5U8lMquQKPsCH2EMjb/AWhdJbZpJrQX/5gYmki7Y
FE0Ba4uTzYZdiw8CnB+rM0fskk9rI0Y+3b9XppN0jba3+61B/aCcAfz371t7ehmMbwhthw5KTxJg
zEpmOt7lqhk0mVumCntHTtUji/qIaKR7yb1mB5UxFj0pfG7HubjSvZutbE3h3e1Z7UfsPf9SrMe9
N8h9zw78nRLTC0e9Dmuo776AJy8DuY/x2hztaLkYVXv10E+H4DliekK7CLEmB5NIOVXm1NrllAIb
E8VyfJ8KbvToHnn3Y6gFOakuWn7N7aEGp10FBSC8jFt8gnuftNQseXocZj9HYIjp80yvxKzcnx8L
KsvTW8jniHuqaBaCrsj7PL/+11JiFdo/+DVSvByEp+BBVWFRpVoRzSYXm/TRgGqjNmuyeDltFvck
ddCE8+3ffnwYxPu8JuDE34aHRnf7tLq104qCAmQ5TbRxBK1Uap1wI8Nk5h2un+rdf5ci5RTf/LYl
IKZSyCKa7yNM2aveTBPUr5eqCniEZPnKrsZBpdWLM2yG1mhu+61wOGgy4iInHP8NcU1mKENApH28
wZv303QVj+Dr21XFmdrOuhq315b+VKobBLIKeSDPU+VEckIZmfV/nQVTb9AssW7ztkFc3P9KoYul
kvDGTmhy/SZXC44pslJ8DoG8yjqVz2rWAlUKPIwF/9LDZUUrPrktLxX+k6DNWRHYt2+At4Nne3Ur
R3KFbR32sadZUcg1cyF9GUMD+EAkeg5yYovWgYQBm8lJ5Mmw8aZcKRpKzn90mGtA1mey5JxPyFJ7
3Ge3CLnYevDUQDcdWB1j6xFmojPUQghxc+iEj8q26j8GNpbMSyNChrCz5R+NUwWzG61meiLSTLa7
wqe75K7AhSWfl6mVgBRdnopHW+vj4vo/IwdLZ8MfDPe2MnZ9wjgiK8nXeB7Z7miQatjFTQjFvoIo
tOWSTzysKHXCdb6zMVTT05JsIydbUjSEm2Q52DkF+pe9Splhd9uV4lOIkth5nssLxVa6x9vrnwto
LpjQmqB+8cYuCdiYV9+aJlyacrrylHvSQgsPKYYWVZmJMBYgctcZVvHbSqjjX17wM9HopCvCkRox
oMXaDBNw+yf9U1878uJEvOJGbMV31/5/nN8+K0lb+LpYlXxXbDQLZaYqeJQ6Derb5yaOfyUC05iQ
LD2cmTCxLRJ94GzWp8TgKXynDCslZAFGfDHh9B1MlOuKRC3nQRZX1enIymaQRf/UeSQjFjMQhtqs
FUi3dT61u2GT06060yiTIto4N1k136X9VMTVilqjZD9ePnvSRffmNKo7DpDKZXVSjQ66sLsI/+1P
e0PNEuDdq+qv3Puwrnj5LKQdvZILFYnHiNmpt8UWlP4R7shULEWvfDUdaMXangMUdyeZsEOmiHXv
PONP2uxLMbjwxN18cjoROZU97xyzSsuWRzeUJmGwVgi++4AIVNQyqWZaB6JOpvSBcnd1dh16Etov
0Z+6hrzM315THHRKMpIoVPtA4fTuniRNp1dPgKQqdTHWxg8g/mQmDtzEdvIJsShm5jz1EfvCdpw9
8CVx/bbdUsAU88lkMaCud8F6bhusoIIov1ejUxnl8nRttwgddpYnJXerPng3Dr3bAxPwor0pucAM
5nQIYXyLiFcInnytmF3inrHhuFZhCEP09v4CrMOgQ16CzmQVJuVFflmxltkQUmj0fvIQbexMFw3r
PsAdizGbRjfHLzuNYiNa4xOEWy8hPyTP6DUneDdtUG4S7+Jf2W4I9cGvwyGQr5nEDSypUpJv1Z8B
e3YlRZlve0C0uGZhtx/jHp9G8/fLBenouCZhqYoxRIqLb8AaLI19sZLZf7erKXExjEBvxXf7SULn
gpBlUnE4K+zgnISUhFe04wOCv1wUlca5BKXAR2iEsH2OlkyaXJjR6Um8Ynh0elCkm0pLWSvntx/L
5JWQt9yVOU0RziSAWwKI6BqtgPDaLFe5h02tI8CMXmSyYSVm2C6iI5UGxKsfa5i5LYJH69lzVrdx
X3qrUNNdv+mvgXsf4ly68gd7tncPASxp/WFeC2ARwGp9ziUQekm5Aeb7mc8sk4dXbIz9pVviI2PM
F5eOSQc813lYfgNhQu9ByWU60sC5kXIc5onPVOtyassVxuOakxt4zIIWN2zmEo3AOJKcN3kfLJL5
1IBLr74XNyUzz2AKNeOqNbcPGl6ch1/wghJQYabPw/etYt8e1hOSoqM3Hj6Fy1jtjHbHfrkJP0nI
H3nQght88dcK18lxjRTGk1FqcYTVGB35RSZsvlQMwE7mKhcGgklVFyRrPjz3kCVPxuSJiNwl6Eld
TINrOK3opTmFjeFeh7OjyoGlpZurkVzYn9t0gTR40wsmo1+vAfeBAXCTjSMCu2UfwsH21NFreFc2
hgXhy+n9+GNJTVBkF+iZtXiMu5EFBb4IYVU/jXaWclb3VAl0bvZJG5O3/GsJzzd0SZ4s+HJjAuS9
DfKaK2JDH8+mV7L/CmzHsz94J6kb+bEWsxseO+aJk/bEZC2pohi7r5HnFSsZg8WKiOyXjcAKUkEf
31OO+9T1Cj0lhCQjf6GKN3wU++0wI3PqH3U5LqykCKgslCNRoeqRTit+Zxffq1C3V8mOfKtfBNgL
zjh2Qu8bjzd/IZNwDa6xcSXJGc1Z3KvVNIRvjOCMpUGKoxM1yxoJrbsvtkTCZKWnwYshM3GHhQ9h
ZmnsZOL0SXvZ/cU2DwzVeL9rR9iHMLlsU2Uuj4xPd7nDsweNfww5SqwKE7ydSTWZxMSfpUWaW6pd
+nz6bPRcDoZ6IragOqIitzjYY38xXA3czMEF0K8p3qqdoMGTpBhaHA8Gb55FxjrVn51wkhvy0IfD
gc8J/HL3YkYwCfbLN7LwA6JYL1UHmqDCikjpVPIswx6UuwVI027YYKpSAkqjCtfHRfNZ+ySfIOjP
Z991ucxExBntWpFjaFSn/I4AD/7BUN+OEn4AZZLhIAaWN9CqDNzvyY6/IUE8L118lCqGvLDPuCtL
Nb+HZ00TLByiCzmHpvFU+8pcBApyDgrAXUA/b7ucEMpM66xg79Njjq98uCZNkScbZ/9h7Nix9vfb
HgKA0FwzREHgCvdx3PNIpoahxpVSd3Le1m1Y9o5jbnm+ERJDc3OmBrvNetbnegxoNbg+8dgiMdlW
S9k7OHzyVk6xu6sm8zIQMJcnZxb0JLmYjw8ASmGIICMWmirv2vTOracFMnu6DD+HJTs8beWLe7wo
6I1JeyStLirGBrbIqeAiVHKntqaENvM7/VV/e8WylJ27sfhgsvBS8ffc+1eYcsSjSuCupmmhEG75
CO6aIrz/7UzR/D1vasaAgiWNTZL/V+VI4tXUv/55Yum0HCbRmh4CNJG85v3FBJ7GL2V9KtdByBbm
Z4cKYmMsG8oNBu8ta9i8T6uybgA29xbVmCV639tCVN0NMTVBNFooTO5jMybhedkOKLth9PplVefc
QyL65JMDy5VGMztkOpmOqkLNeiAuUTt3HQtDV2Par9YVGP6pji2xaTJTPWEjJbYyMcoZFGUHnQy7
X4OL4JXmMz9d3YIP0h3XC+9EyqrI1s4l+751xdKgfPmsIZgbiYoekEz57c5Q6XnEjZ61FS2HYogV
jWeY3uF4TaYXZNhhd7p8h8awRxvhVr/YrD/f4goW1d4JM7N3xl4MngRw1ycvjbBTdXoM0zHKnpOp
x9qI66li+7Bl6z8qzI+wtfhPGWwxqf1VTj+jY7Cakz6JUWBjy6u29KuKOTg3v840cn7gFiw2lOf9
sj4TE9U3hHAxJUNYMAV7/XIqB+BfWBwZVvLSjVhlpOBmxr/NNdTn/CXFJMQx8D/Q5AhGU9ny02JI
WqJWHGdkiNdtE5e62V0w+YD3cWNspqWrJ6rv38P2pkY1hTShCKM3pcx4ayE51iZJ8nuFbgzUDqZn
yVwcwQl1mocCHfJw4PDH/w0+1nHBgKpDD825+gjsmMGjC2wJpqyP4KHssWUtd9XPvmj36xLyYDDA
IOkvSfBrMNPDEaUDLYCPHm+ym3bRIHfeYOLruFSNKDY4Q1h12i8WelvnIKjHiKBRoYgO4cW0usMX
lGgHsIwpPMhjjjMd/O6okvnJAdpqKE+HM8MSZjcLmalBV4XNQvgHpA9FHBaWnJso3nLHA6x3+w5T
liRMnmlFR/3FlkAy/Oa5M3EBAL0P18jNSNWieYmX8ejAp3axgiOCSgqci0J/7DEY9JmCcnip8kNa
IjJh2/FTmu4RPbb9/MBmE2zf/gXmL+R8P7Wp6FXyF3RKiDRM0bndZfmz2Ho8zZJTRW0aMJX+fA84
V5L8J4OBZW9k6snIuc5vxmzESO2jDUztoA0W6rPEzADr2/gau6hy9y4OKhCWo/jLHIjLuMNbZbsQ
BVl+QWotouNJtFX2J8byFVVEAJBW5PVnP5Lg7HNecbObWKglv9XCbX3glqTRyvmazH8VhufkvCQW
CLTvV5x+7bGHboyugbAbXB90BH6eoOA6AqJs9yimE7bvJnsVZmc3/XXMYaEhMZ/EdNzGujC0Wf/G
4wwglxwYmHEQUY9gOAne3w2zoPxf7HNU0azY3Zy494SXJN+fVJTQfDJkGGFCijYH8ZRBqlCK/y8h
WBRBKNQnEtHiPfz2RZdngB3tbZhgbmTLhNf5yR0FLZMpOcliR9LouRH5WoKUnwtNFa8PyE/TlK+N
eVrDhRKkzb7HnyxwxogMjNcyQE/UdMrBU65/LhsYWb7w99dEUXlqpmOvxYdYmyfc9+gwJn4gshHS
k69/vnIK+7UZUjybnjhrvpUzIKtBkJQqo2/HW01P4AUiHEPsR1qoBoDM89tsxo1sspTPp9CgE7on
duqKFdSMSIanlcM+S822Ne86jvOmtuoAIx99PQx93412CohV+tsam14ym9vjIyDzIpDZYCvbBaQI
pGCeLUgRYCvLrtEEl3CLlzyTAKWO2HDRVfKxnhb2mUEC1PCwK82OhV4Zjt2Tbq9KPiX7sLQjc0+t
b9X2YHYMkmFkIH4gPdL5XnN1I76X0rjdEgkMq0eZ7r8efOJE+Q1TrO6G5bMbykAdTBgpa6naloNR
X764kqoHqbqRCMAEdgKVQJIBA8rDucdA8GWWWULeofB8R3R6XQlBXvk8WsEK2IqpwouA7gyOUmwM
t3CpWZkelbUjES1AihMWyG4CvQdhSRn+QrT+p/IGXpidG5o439uG7Szvn6wYi/HB6xpY12v1Z5MU
Usr0L4k5ISMm14OWndN0CMOJ4McIc2tUModyyoC8g+VoC7gxhJEye3+0vwQmyQ0arRA0qmkoYQIf
WB/vzxOfopT8Le2x9/DNLPLlA7Bc6Gry1WWHPHSOD4zjXlHB6umGw/zemxo5/HzTbgFqmEWEIayg
6agKJelhPS9eB0QNRJnpquQwB/LVVugDGPRrsO//cjLx7p1KrAsz++lBeR4SM6CYwZL+r2ioiVqA
llZDV1Fj8uUZQfN/fKJ15bEnakyKMCRESLI95ojfWq8VLMPlW3IRBSbod05iVgzTmd7DjpLrrX3W
ZCYYpetFW6pYeMvOZyVhuRkny8/uQLduvAFla499V8icUy6oX1t6ZWt5x9O1JFRWzGvduPLn/SpQ
B8po+hJaZSmZuTCtcUyg3YdjOiOp3JOruUiGLHt1VXj+8m7MZF20p0huBmCbSkSSXQZZjUpueDCV
oA9F7BmnYJ5ucPwqSxXm9cFOwizrygf2kcdRK0nmz/dl25hjIdM5+/KSDUn3R7K9puZ3sr8gSqwU
46WLimbMuN82J31b3YR3SIA57nDWADzK2lRBV5ZxrRJ5SWaSfJ4WIk5/+DXhefkSAXhI4kk4TmPy
KBC7Sw3PJ8EdgUcOpWE1uV475BhPURVOebScummEb6KIfRMlOeiDp1B0Nb2JdRp2Fp4XPpXCNb3M
vUA65cMCNvl0YKuWbccrIEAFUFkJMDSOWK4jdQITcayjRWbTlU0Y38iQEnNa88pnixhx0tX7l/Ob
MSHhNmThNrRfud8AMvFBX1YgoI7bNtt1R9qrdVNsJcfzYt60voG/UWETeXKqsEna9R5ajior4E9d
VGj6tU2ObS/OAVQzaOjjHnSIDSrsb0FkX1MSeqS8cQfbKWujBaUBrKPtsxfRZz4BmfiM3f7C7gCJ
6wAT2TpNwqYByqi1ssjwWmxV2oOl2sUOFvtj+zHf4YCIgysNwJfUE8h/xQNqX4zm6q883Mkfuev4
XXxTF79GfB1sSdKU8Vjik5lTtn2/1SNGjv8eiHWVFRkL25R1OBQy60FoicV15C8Of9FyTLW1YA/Z
Hq5xGee+rtnb1do+4sE0fYkj/dOgLcCR7DcgUk0F4cYanYc3mgU/GkVRh/8F7kLjxLNWnpAnOrDR
jHRX/KeeITtP702d5IfPDcNufZyLL89SbRZBPqVZ8+3Y8U7e5aHDXt0WIWNQo9VG50c7w+NmDzrQ
hMWbr2fasvv5MItM2Hztjbz1koq+t85CUEeGWoEEYy1YEmJLYgx7+PKHn2wEmzB4LlhZyn7DihBw
FgJ92XylcR3JJj5on5bWOBMWlFBEmkyjfwdER3WAl6sm2f08rAW+N1wlV8XsOjDpKfBbVKAM82t+
SqN++Tk4hXJX60Eg2eMVrNxH9vlil8XcHQ45NgM9GWrVmqkmEceSDU/lTg0680Gwk7RBmJJj0fR4
ozen0ZQFYGAaTDgf7X7XIzvfQAZCXIrvsEqNscsuSlpChoo9UQhJG/a2oociAsVz2XRuJ3Fl4m56
LxiIOA02yL7hwQGvg0smIJtEL4CdOVqhsGnvHA85vLyS4RLgT0uXEVva7Ny9jrWHWJjNaF8cLYVg
DfYXztRLUh7z4M/1aKh3kgSgk/cUC69svZRHP8HLku8DumRhRUsGP+pchmjDHlmNLDne4Zsx/qLr
ha7tsmSF/l15XQEc/8wPHPtxzvZChnxnMHV4r6rIUp8yw38ShcHK0oLH+I4P113EngGSZivLhi+n
RUcatJ0D2HICXShIgP+82hJPG/Ns3dR8S66+ybUOZNO8rnOP9oDWe03mahOFPApAw/BuHDPvUmko
3ngU01I2RZyJc9Zcb8uuxv6UtbVc01otzmrb+v28Djz0y/uTEHEniZHmj8WrTCcg2NavcEiN3laD
Abzn/kaIgMxEn8h/BrnLBvi5vcjP6js/Rw7ns/dofCyJ0MF4vVJD2mZHR1DfDNCeCqFICCP0Vcjk
aoRNnOIAAevT8tMxeceR3qtFpKsQbHnukMvkZz2IzAU3pvQzh/dnrOupcGIcjRcneWLLRUF1utV+
gmogKhZwg9ZkAP0NpeJ5cevhjtfJg63cgVzgJlw+/ghTeOept4UcXHQmxpb5Tr6leTzj5Ts/WjTu
0HvRZmOnX6F4370CVq393y5n9Q56B6RqOyaqsiQXO9vSpS5AwcxIx5/TdLmG/wtMlqx7f2qJimrx
nN6zmMDxBqgaIJTqCYu2wh2DGglDGbSM7jyPyxhraNXFIDqH6Ox9RpXWNWsRg8O8dZvHSL9/jFhA
7+lw/XCRnnoE0KIbaPiP+l8E10XGE3zv+J6NaYvgGKIhYG6LOyq9SR52Kn6IiuLoAOls0EA91AP4
93DKFoMdfXGD1CRYeKBNhWacEsoOx4jYihqGwkZWBjHEK1ugHdHNGj8Rpv4tLbp3u3MIwfogcMT0
BepAlDgTepfmhxh8L/ZjwvoTyG6L2wx2diJymU+nGonHozOhqgOCO7Wmc5G5hbiN5kgpViaL68uu
2f/W3YoftCsEIW/5lBqrB/38MXT75CVleUknlQ5/IHGMQf0tIpKoeCM20cA3TqgjFenuSeWmf4eY
8kS4SL18YrP5JcmnEOp70UCkLwbmSo2WFAJ/tr7lpGOLHSH3d9tAldQ9fY+fJqP7O/S6Q+ifQ5YT
6moumHMAEjfV9L29MdiSngBGVA9NLfNWTETInxJrbk5rfMt6kv1gd8DZEg832FH2+fMwy6lAbxQW
QmPoqJIarLW1TU4RYNdq/oIDV/hjTcBLQuO/FWLBdfXLgn9fGLnyflLbr2/u1lxx1M00bIqGna0T
KugTbTExtBhIFMd32RNqv2SHHh+COelAfu08WpFBGH5J57C2/Z8k8EB28Hg7OVZK3nh/hKDKRllc
XpSjkzP8xbJzFoK820FYrE4zZoJgfPPTlWJtBQfl+sg+9qXWqbLb101xHgMtU+ADrhHG5th2KgPT
RaFgY9ZItyHxsf0Ed8LxP/dl7VGiUI4EpaRHO2pa6gvGB/Z60vyVLxrog1p94NqgLLB1aJPoqXi/
92rkpj73b8Yy+Do/RgPbCPlkmbBUdjSEkyY8oO1yaMWKTD87B70CGTLFXnfSYoYfP+5xdmH2wG6a
Q5TMYlHb9VdBRXTMhMB5JIXYZpLLabja2BvoeEH+I1cEB1GaCSU9PJNcLepqOw9oSq0BONJktgsf
GwIsoE+HhO0UhrRt/Igf1CFzExb/iFD1zz8FYq8a7zEVI/sTQ45Yzm+YhVqZrho/uf5jl/6Dk2L+
KG6JGr+mmFoKCnnebn8us4T6T4NsYiPbjeqs6XRhktW+OAcxOmrDcR7G9ehK4bHAbiEZv7TJVcjB
Q8QOWZcDlvihye7jN0fUkzJivvUSPtyt2L3mkT5W7EsYi34k+p8qlratyYwNLe7sBahV2K6BSpzG
sH0cwXhcQ4f1ZMdoC/NVKO0GbKJkq2fuuaZ9omRAMzxTrnGPUB5vxtKgjit0RQYa/L1kYFDtlg2M
GHVBQ4zQmpfqITOfEoPhFYlExUBeacH5cnA33EfN5SAE1lxbxeG8/U+x1X2wgsRYRlJX9DenrBJP
5NobnP+hNHcMYVleusyPLdWeFLS8LG72QwQ9EcptSkPBLtMdYHkLQDb2H94p3tjqBQSqRO3fpXzS
+NjaBOOS+rh9yVCC31mBofvc84sCmuT5Q1T3DL+PwFUIr0YTbLknh9b0n7cm2qybM6MEtSppNySg
tDUHbq6RXa3KAzNxhPJxWRID1+fX6wOJAUo/5qgtBsyoFROp3xHL7EvpfrHGEVTn/456Rf4k+mjP
CDIQVX28P+mDPMOw6qMtPnzhw7kZVVUiZt/E2KUn64zvQaNtpux+lpSKbg9DG9kYBSznt4Od7Klz
twgkRYJJ5F/fy5+6C2JbSgW3GjNzJyZBBatt8J0dWUL67yqSL6anB6+JTeZMp0mdOOirFgCxCMMK
huqCWInTySPHl3/2jQ/pAFt1ma+ogTu/TPctNmuF/pX6TqKK5aXfK7DOegF7NJfl4rWOV1MUGHMO
v1RpfCcQXMVy97rjF+dU9vC8ZRzgAcAaATKo7orLexfMj8YG2rCWm9XI9AiQd9J6GqRoDnmJBarN
VHgQ5u8hHJSndfVkqADan6UAk+VWTs57q9t8Hf24JsfhaCMlXjbVJ5fHlmJTbcYKmC9FuC4AHAEs
A+sNFfz8Xk0C2v4OPC8DJ4rhUfw74/oUkkTkMqkHc3MBLc/FW+DLV4fZUhWwZ+/mMJ2W53y7yac6
6WzGXbcSxDawxEdKUdNq2ZGoJeRM2gyPfpKkf4O3S3QcLW3Jb87NTJpfzyNh+9fNi6UpchcBbuRA
aZcx4pqR8FGt6CboSfFLgZQDbIXynKYjIMWu+HVOZ9juidJ2JLxpONWPf/YJX/+5ElnNIkpfvqxD
vE7aUMUTTZlKhEob5JQDZ4SAlul8mVlKDCR7ltJmGYGuV5E+50goGn8xayLoiLVGHZG534jHcUHY
gr8jj3o1hlMlundT5SQuJlOtARw9HBVar+6dboAp5pKEey3kWzNTIRpZc7KH05B9/tX7TZfGSYBL
JtZZIWdDudQcIizFrAvs5BOyneBJsKeObpOQR5dx88Wu2Sl9JbFgqkhW79LjrL83WGNy3JMI1Ue8
LjgsgxvifkXisN4sjdfDiprG2affT8MTR/nRatNUF7TE+mMwl0O/LBUjYXO+cTMMCr3pE6+C89Ob
r8dsYkuyV6BBdGlBvzAXq8xhA8wx7x7dlvuZiTeqHzImWFeHk6X9Ysmuzci6QTTPsLPSHlAlJMfx
FJoDb3XEs/OKnEjywUfips42X9gouV/AjwP1P0qyWRPa9Y8IEPEbCM5wfWQs85mOd6sG2Nh/2fRI
zrwedFvqM78Ewq62Bp7zyiBemDrLfMvXpoQwp4IYPzvP5tvS8QsaU9p21h1wMCOraOBWiOJP+v5y
PI/z/uFibCXXI1u4KJaE7ImY7xPXYzDKQR0Rq10HIfDQnVScHHoquMZv/yUEZq8kouuOsdlGi5bs
7VZI5sIFjuqs0mcepP2eWzcgU4PTNXajK7NVba++dWQGLzQriR3SxNii9MMYqGVlDFFCEn1VM0yy
eMPDr4wltBwZlvBzNkgfxKEY7S7OmWbjyYF68uNMqHu1az+W4PR/LhWCnxmhNDPU08PccYUuV1DA
znVQEFj3LEFzNzt+5DVNYI+iEc0yiAZN9tmOV18WT29HG/7anJUGHfh9iF/OEdCpNMSqMbyljPI2
mDC1dKH5TR6lhf9D6578DJB7KS4pOHXR8RfXwixqeKjsA2oTWRUpGjSXG2G884Ww6k8F84f+ef1d
56AN4nwnRRH7WpZGhL2Rh80DCj0EHhbZHXQ46eJmPx2OjnLBNUQIrQ9gVLmb8+GIEEdLSMzUuwxM
rinpBOxJ8U7KcAAaNlg1SVBL1nRxIFl793YKT46mOfzvaPjPudSBMHMmupyrZ0kGJGqWXUHWMjHv
FMZKOn+JGgDLgark/n6Js1LcK0XSC9aS3ccad+zjRRmg9YZ4gCHrd/pHZ7v5XyPBhLN1y45u4Lio
YAOPAMQAZ8m5TOk2z9obz4xSOo4fPTYwt7lZhd+Q+Us4B6vM02tm4fKQHC5NFimUTi5dkTGOsuXo
PVZifVz9nYFCUl79MHjV8J96uBksgcC1SxV2MhKtSc8twJ0PB5VhMakMv/Aq5SA4AkFI49G/oLNn
AYegRFgtl+KlAJLzYsELgMwIT32K56YH+7EFItQIgfZUOHFaecbQAGisF2sG9ovx/N0AulBP3nLH
bZ68CVZEyEFT+nPv/5sPkAHgQ26IlcChI8KM4R4HiPmIldGiIN3aCgLB46gWCDrigJIPnrevAgXP
T9fEkC1zYGEil3gHAmhnfoaQclTNOsnSx2xQZ4AdF/ZSf2Tf8zxP9feE1o7jaf0mvBiJ8wYB+a7P
g2Xm5QTj9VsPOdwSYHo8/TPddbEO0itAwA3Nut/lhuF5LAzhaa0wUWqkyqdzUzcTU9Nsowsge+Uf
0zXDfErjqysx9ORHCg1v0Y2wDmlDinJaHDiVTtwY36qCn8vM3bNZL8QQ317YqcRIjrsc+pu/Cqq/
rzkQGw+5FuqSZ9AeW6VdnbYMvHHvvB2kXBYdKIVMq+oFgf4tVWD/FPqJnyeUd5DK8J/rFs3bp+2A
2bfJ8lMDIyUwQ3/XeOCADlB+Mzk1Ecz28Q+uxbdclKYxyllt3k495Z7/pOqd0odw5Zz9pbTdRjV2
H4XxahapnRhFkvFWfFMvPnQNeeLauS1JpdCcoIcwAVLfLKuyhZq3OM+snd8BGwx++u76v3a4MdGD
3U7E8vOHK3l2HeEuOXZ2TqQTQ8CdUbI2fsXxJr0rHKcJ08rxZcniA2EjQwrZFSUAj9UzffF6wTjN
yE0u1/lAqY47EjEUMLI5HBc+1rT/zF4xt8WPnaQtXTDrca0Aa/Ci7v5+lEiEmkVLJ7ZzdtoBrbah
KCT1naYW+JTqwNUdu42FjyTMIySGpYdFh1crWi8NgD37Vd/vkBDVYEN4Ecp5wlp4OXc7nfsWMc73
SqyBPevKhygDBN93Vurpy5FCgaUggcdAIhdgIWLuokR7dfiuUnG7JoGGCLpuwE6KXu2YLScCWVs1
crE1RW6hNYz0vEm16VAISLKxIWF6l3O1jjb8/yoSLlxOPOFhrvTpBNpMD3NgaHxK9mUHAZwto3MN
Do4nWV7p+PArHiBnVNvxyhhMgESSC6AZ3gnymTCew7eTvM/JCAGGLvkDtKLNTCsHdJlJvjZAXnJL
X3r7LomXc+D1dIHnG+A0ArRusMtIiEhEkye6LYRi8eJ5OyOkiV5DfbW6m1cmHAUXa8wy/fn9g/mr
Dm4hNdAO4JUB7kd6lpHMfh6qj1oBfBbWS3GAF/e91d1zdsfg00tzWh1vFuXfpot8PSPq6CFoFBzP
jWvHGdwc/Whx9h15cQ8XADATxz71BrwafCKM6X9AYTSD0ZTVl8BFdPeVCtaXWK6wtRhjVWQsO69D
oqW4uu7bLvojDWfAF+mdIuHWPOdb/X11GLVZxXbQNHD7OoNRcp8J9YgvgWWhJ7wDZRnq7QN69NsP
S+We75uLaHcgzsEnUQEG4cJb1kD7UumQWdLX/MmIKoz1MzAAeJewxlhlyStZl6ta352wzFv1KZL9
qT7jX/gxNTNS1Qmi0x2sSIaMaHYzyKHLxeW0JV/yxsZo4DF41ZA0KkKli3LJdpGGTLrvrBQdeVkg
THQC+hSP0KI0qWkdCFNysbbPj/CN8K4ENBGV7vMYoKy8bEw6KWrLF4cGEKxO9Bn0p+Ktp5StN2DW
+U/GvKbOAsUwSG0z82ofkKHlkmSQX2ZRqVOOnlrITGV8qzZ/5KxlR2wnsT8EhJHZhBQj9H4hReqV
rS41vf1zwhVs5aKM8QizLa5B1jnHbHY8HkPTs1GZ/IpxaeQkqyoGTtvNXYc40UehRKczlBClfNCb
vOROF3BPWIkq0DbfHcYGOVxZa9ph+w8A3phYuT7Wux9aLk5AJf/FenZWM/ldUymsrIqVQyJD3Uou
HEoTcde/iaVFef0MALGXaJya1eQLxQFntBx13Ul3jyCexgzcL4TR6F9WvCdQr0EOEzTm6h50A8gD
Fm5O+8GtOZ18GgENL2Phvbkj0BXk/PfGGgbUoqqeXpW7VTK0dJY2miR+px6U+4Cx1DvY0F1Zo+17
EhawE9nOFuP3sN4SOXpTAt19Z7+P6HjOimr8HBuYELjss5MGhEyNolODLd5r466YADnpeLg/qRTO
LdiAbCrjpbSqOijC77n9V8e4NACDIm84FfIkQhIM5YVvueQtGXrK1vgI8qMp6hdSo5ncx2N9vxXh
Nyf2+Iryby/vDmIhCpb7yZ0iwrmH93VTXL6TikABkhV5T+PUQxSW9JyNzQfv40DHMO1BKpkv8zqQ
pixHVfisxiV2A8STLoeXK/cASS7Zvcvljv4beAGS+JMnz/f4fB1wh/V1RWEoCo9dwm0+je7quG1+
/z7lF2MLTwBID6VNKPI/SKqypqf4eNaxCFoHkic9FBD1vmd9tevFYnvUvGmJFH1tqcaWslwnt/E+
O0y6T7jIEgC4+irb4Ylm4G5HbeIZnKtxEUX2tP+9EPoOwl7FLP/PwDtmpAjP17SmITZKkkZE4/Z+
o88DKidkqwZUAqgKrBhUn2t4NeWKhfgjVAt6EnCkN+1ABch312Fmz4rUJiJxii8YHleF+gYRHaZH
deScUUMUTznPH/+QJBpszE12sokvkv04pkJiuEcu8WZNzscqbnYVoQoiw6FZ+N72RHfW/1UhxNBF
Ez5xZLig2aukKcfMtm20z85q61NYs0BH0hwHkATyQ9Vo4ImRiLG3yrVD6mcs6IZOICqqepabRiAr
+DogeEKPgYE384bGs94iAy07FfnsjECwKXnNQSlJ2jRGWuKFouWb7WXEBbLCRLO0HJDITucntdy3
KFW9XUBRv8R3dyUjUcI1SDMSZbNbDCqBFIZ5Cm+1G8teQBa3thdofBsWUZrYRK6o4EaCMAIqBCGV
A0+5kd3hkIYZcCv4QYC14GfSgb8N2WmNmYmUylTPTX5hgQqrtSCeBbtVmy8CH6nmWNjPRdzy7UZD
QK6o3UjK88jdX45+GrkZkBA4mZw+abFmLSJMu+XeYK6a8CieUBlJR/pWXWJo8/zVp4LJ/j0UEd8c
7QF2vEYs57Kpk/IuE7wSSBZCGQLccxl9MnDSLDZExxJrmLyD0FVD5EVmmuKKENPRl28h0F3JJX2/
UC7of0QoHpC2vFaxQ6NunahXgKieXpWge3ttVl9ODYDWAFFvp1+KnnZafVnfiCHAsqBpzF6qTqb1
9j+UIfjxaMCeY+s8RieqC0BVuFAugDNyc09OxeNqI8joJ9GDFQ1PBO0MdIaAGwRY1Qok/ILTeJhL
pBJBPChaK1IKMweZ79/EBRGzsA6g3YscMX7qWLA/FiB24eebQ0/3yE2W/V2X6Sf4Pz6AaGB0tJAV
ybXtIWvokJeMACPGM9Q7/rfGaf2yVkBEO0LfLyKnQUFyHcgineXkgpuD4GoEbG6v6sMCed3z1TrT
edzxgbPeejtx98O4HJHHJcx1I53v4QXSVmyjqvXmvQPLDXzrkg9MavU+eJqPmgyIXJNpZHWqm+aG
fjIiGUNmfeUBqifvQWNdy8DRxdyskLXCunb1WIhyyOoNqqCDIU/jK/48lwSlve2GTC3bTNm6EdRS
oDkh+qyHbej1nLNWBCM9AUHyN/nMjHnfwQEBjcGpTyGbOxaLyQ62MOFYyUYFLJH+caf4/xFUtW4Z
yeRedkWPdSFfXzToXVMusKFh5RpgcSbrzajNcbCcQUiRAkSSusJW+EMnNUW1q0AipCtAOISzRu1V
IncmoAKuHmebJHBlV8TyujPp5UCxxrCSVlyqI4YadM2I/I6gMnPPHTJP1vqE4SldqWKFirwI6lZK
ZahK5tYgC937m/VbJhMvuniFHizFxOJs6XHb5etpYMDi9LJbZmRsJOtuKp1ofRJo1lEuhf/ROTjG
6czRVvxmcpEuZXk4gJPnCIirM2M1ixZX8g5VJgnaI8VbdW+XMdCE15v6ATOnrmiqw6QWmtEZF9m1
RwaGXCLOBS+Fq6ylPrYT5UUYneQNin8PbaA3tfpHOVLRExy0StDDeRAu8DwdSosAWRPSlctyTWGC
+5E0zuJjxdrmJtgi7/3VNzGYSfkXoJoTl5FpVpNyzsdl2LQmWatZW8bzUduglBJhcoD5+dlgJNY/
pW0jS+9X3w57Q0cXRpFOQO7D0OZRvRSgl824j9uOorNphljqWCn8epgESgXvMTAKoCEgSjyn4N3k
p1yF1NhXp9OqSyvgXVbKYpAEG+BqPLTzr45JlNsg6n57dp7hRHWuYy5iqpUsi0zVDeU6oup+rBvQ
obAU+zHqF/utBLuPVQ+lBB+vNb4YTdJxBdsw6VezMcprV05ylk0dnL/D8ZAbcSzCQA9gVmTEncbB
w5H/TTz1kEu1Y/cRH4HxkJoSDNJf3x9fqIpBsA4hRjVsET0sNZtNad59YecRc6hRDYWfnG8o2/bo
KKnU6iGd84uocWvqVcyCgxTEVhdio4cPY36/N3ogvPiMPhX+r8C30HaUtq5DmJhGOxLXFkjWs+PU
bv6pP1RlWmb2JoBZnJ/F21Ohc/0gobREzUPhxn6dak6zD69d0jtGOlsJOCU3hVw7j6W6ZaPkTecm
3p9NQpOktn67SkPCOGNfbJJAkERQZx3vo39OyXDue0LU0Kl7fEEkD80EtXNK4SZQCAfA5eYZNNnb
I+6Hp7RDamt8ajXk9qlnZWizWCMcDgWkB51dtpunaFmXkBGArtgxXyfZHp6whN/+t+3sD2hxghAq
vMg6bl0AklY6etgkXKiwr1TQHOp1oJ2sIf9vzqLAs1DwD8wE7TA8bm1lBYN+TJQqlQ9eqwz5SP3D
zNVd/Q6HUuvLbiZck/32ItOTnGrynFVhaqtXIofc5tjQtrziPWalYMH/UP0VfviBFLqdLICIVLXr
uusVkyCJPfkQ6/JYspCQHSBq0dW6DCHx2DmsX/1CZuDVwmDgfff46+prCcJO/A6scarGWM06jnnO
a4i7/Pwb2U9eZoGdTuNukdkA7MBgyQK/fF9bH9jYAGaiSlX38Zvlf8JkLIdv0JUCR6wNFSUrLI/n
nm8wrjyCYZuojF37NsioxMqm+GbYg/VcHOBkr/mWESWNpO/UGcRpbRf0ut3Qf2UW3Smv1IiYkQwS
VWjrbxpJCKXNSVTw/GmhcbUMy3MKp38Ow8XwAQPVvzNgnaNGo6dz8E5uakVgwPTQCDjxCTGZjVuS
RxVZl1piJW9LO/exmozCUIHisEU03rHruyfsv3iNQE0TT7KGBWtz0M1HTQQodyM/8ilT7s1JZTMv
m3QyNdVffRV/LJT/AR9MBGO2JT78uU5ksHMpf8m2g5Tj8AD1c5NOjgPkJMbBpXcjAGTbNnaom7fh
p9cDzSd51KHKKcofGGdzQmzb7nR/oLKymsk0mcpis2K4+d+sDVtsdkPJOOu+8B/ir8N6JT5D9phq
EdhFaTbf44C9pzIaNWryN+6Og6WKBfy81PuhoXS0u42DPKUD9jh/AAzA9syKw2CSE/gac7fZlOJZ
zVC60ajSKsS2ALgdDTJxS8/+j34th5oOGQScaVGU5zlDaIqHVhv1H22KQq3kKhQPckDloYCGEAuO
GVwgVT1vWKRFH0ejOwP5gYqu2gpRWmKMYCQGhEOyqLEPP4xVj977HeF/vw/2OhVN2gO+H1NtgCDQ
M7vcbifhVPhoLJz+qPzQGWoM+kNi4lKb/v9CLLrg6uOQvkB5o0ExXqp1Qkp+hsxonY5J/12ZY66Q
80K0r5qE+V2UjohEwKsONKCHl/FYItO2czmdgIZ1wBu6hv11JF56aMO2Ikxzf83NLiOVf3r0Ykz0
+vblFZZoqOJQsVri4pVYBnZRMa+yjuutFAMDMosCPP7QgkTTlG86re0rIjymLiaX4TYfdgnr04IQ
Wl9xAkT/0MqyoTAD/fWu/5fBroZ2BDA08F8IZ8FR3/LKE6rToQz66P0mjG8e4Iifzge0NTXs8gwS
xmKib12u/simIWOq7ZkeYKnr1+iYKc3aN5258Yvqv3HNyHZklHSQhaU6iKqkS+I4C5aU/auyoVW0
SYE3KQOZ+uUjEVTQCSaUZ6LlCvAR4bpToGWFp+e9Lth4bozjmNLR3cBu1jfw7tFVCooLXbv9XHA7
1u9hc/g+2eLxeKeIQq1DpjDnVDuGaW1VVH0iD+U1+gLDhBJizK7Ic0PvCYPzArxNsm8BnDLEyLeq
X1zf7aGXGQfPD5+m2OCIVtGQFV+v9wwrOLirDvcdu55MjyjOVTcGLYjZZVELA1/cxjpxP6ZjEViB
Qe5Temc6lSAARnyUQEcMLTJmzR6iixOPXyzHGTS9LcGSuRt7zgdBlZ5PCbqMFusPX3XiqTaEZS2Q
2ClR9IgpjowWJXbKb44dnc5ZSYlvgY2T7TJY/vv0V47PGtEGmMQjfG10Mv5q4eFeQ9LDQZVbNbDJ
6qt3iBDhlIeujdI+q1kQ6gDvt0ZbwkX43raGH40mu7GaniPX+EMmol5TjF5PFFBDzFWIm3U9qxbI
KmYPXcf7wSfv9zydzNBaaNRmSrZuH0cHIRzaaEyTBn0POe+DREORHcs6I5lQV3UmO+d8nCL1ODG5
PyvNUUvvI1zoPucMczCIWSS9W2jU1nE5rGM3XvHoNGnn5I7h6IEoDE4wCA93ED4nqw+/BHgAbt/Y
2emdUKhiTyEogw38pUqVKKPAk2Rvtwn4FkxoTlncBzaYOuPoP8rpMakgEahVF8iszAnrGEvJ3V+/
kqPIhlEdmOTsPa3uIUlncBMZ/dPyde+TQdQgZDowpboGKJcDnwJzGGN6Y5Gh1q5hJCyfZxmXtJdM
GgOeZqKnQcwBqU/eABrsFcrzugtBeca0O/OSaVsCBBzRrsfSMSltsO4GW707b+VNlBvjWQw+SZce
0NgI9ejjijgjlCpAAoV9StxZG82QKjKw9HhwHia7jEvnk6EqOd+ANbu2MJYmcK+VPDZmHmLztqb6
WFA5bsKzLFLsjoXx41W/mzPcoyFFxwj89jRWysQYfk1LDbpjfA92JnMZfUb16lqi2GpTUmrTxdI3
sfDKcOy1++OT8yrciArkYdKntFXW3eRl33wnodvBl6gwUvfqmwOZqG0+tEBAKmxvRR1L3OoPay9C
XdDXr82+Oi+ykUDncIj4oFugexrCn6fqpLlCiAjh1Rx92vagsjxcOEZ5NeD/jivp29CrqrW8dvgj
WKpqU5KNqz9iLIrbcwspOCAt5g1ynLBinIPJ7Xr7sKSC24KVuQ9ZttUFNYnPMTDKl0QJJgokTtkd
Ki10Tb42Ur1jR9Xw0D0pChQpKUOFbOn4m0bqywcMV44CW/sDJ0vDnvXPKROSrYf10XqCW+vTd9UP
/JENPnpnK5wqJDtJb1JcUkAgGPwBfH37G3woaI61ZQQA/A+XXZaEiAwOyRoCYfpvDkp2GQWZ6Yq8
PLYInL4s4wax+FXQo90fBniIAwYCDeAhZW/2RbWs5yWwh8rZAV0JIHfAfkNWTud4XNGuxOsJ3JhA
zN1FLPDNu1GSuTKojy8SaAT7caD5InDUpgCV7f66ASYGXp/GzHWDi6W82ZZdDYkXVtc3dsHKJzYV
1B/mRERj/MRcL3xOY9LhmMWd0+S+TmRhMzWOGAu8XPk4gpyuZ9gZPmgzWvUe8Qbf+WxFYofg7dUt
XqG75uxW7N24GY7JhahfVolOaDlF8X/+buEs5ZnUaig0vzguWVGup9M5KaNSvrUbCOm5JQTGrzuo
x3xviZsTgsVXEICTVyA/hQI2YqU+9JYgLiaGb3umu/pIwlt9JyC8WBv3voWVE6pfTGZG9+m6k0V4
wBnWUBMiE5m5g3CqKr0hzaK/jhdIqHpmy9FB15AAVax2Lsr+3Cxv1DvkVN9eME9OQf36LeSef0/J
uJ34/46gfTUXVI0WzIi6S7Iu95vTjzR7zGqgvbFLh7Mm8lxx1i0R652vwuS/uaXLqyOqJ/aHW0XY
jzVbVvsx65hHxsXGzKu59MdKrpT5eFLR6m2N18IOVzvvvXdBLgGfQwiBAsQjrOuJg2lVcYWPHIaz
konv7pX7m18+Qn7c9yok4K2ELPFd6/ME5nBKqWd/TWHMfCRord9H8CSsT7QVy9Pe9Fpk65mQOodB
uZNuK8x5HxJUQMv8FdVOVhdgKEGnq+ZKQD4KoTMXgWYva+CL5GhfokkP5pbHtKdhNhG7gT4sHiiq
XaFENZkVooudoAfhfntaz2fqMHi1WdqVZ0iu0i1QrsUaeOd7Bb31mnnCRAyof+U+hAE9ERBJiXP/
zQ1YFb41+cMW4pDOHyhW7fShSEBBKhE8y/DtYpOrNyqmdyNWIQoNs41pe4k6Juz322WD5Cjg6WfF
/n7i6xuJLLj0+ivNbpuf9iqX0cX7Y+39PfFmbSn57osQXdAHwHT6wGyLrsZ1yGk/8Bm74ksceOxj
ngQUJNAYg8ZYjshhxFld7Qve9Nfn2l2SBeXuqtwyo0MiFN/TzHBrJ4/uauM1d7a/JCt5IVnVd0kP
DUdlP5TafIhmJsmZt2uN5vOHsmaccRueew6qyiD3JHScj81b+Y25mk8S+zu849eWSSamFH+zeroj
+UNf5WGZuSazhsceqRmjfXvR+q9JQ32ABuI5RG6/IUKUUPHEvWeK/xZX3mlagoyoC6k9PhTIdkle
eNqGicgBrLGTr/C5q5heQI0lIlpKp5sLtNJWzipHVZkhI85m0PsiKhDMasbi0gomvI1YR6SiSkYd
BK5sB77h88VjyXs5eIVz4Z3R6AjI5viUBDhwDP1SETULtikX9IIMzcoUqTyZQ1kxsRdvCUCNiq6D
G2ODiFtwTPLsOzUkAGa/UNhawrENqJjcJKza/1UqqEC7BU3aE0rN5bJf8Gwj0BciTJoLPQdsW4xE
317jI0oqfUKAHEhewAqIu50cLpanjb9ygAsbRog2304OnB/0VeN6PbOly7vtaRRRnm6vUMjid1SB
iHt6rCIeSmRaPQ7sSna/YadzqRIvCQJ0Jcb8iaZxyOb6e3Dqz2ZkQCPVLI6MgKoxXwIgtIHeyCOL
5DX76vNnD3trfCtohjXxfjZe2h4BDd6vY2OCMTnSSkXvvLSBNN2NlSMVyvxoo7wX4+jVVKWUW625
vBMqvB7TJ2QQJ3iJKLFbwF6R162UffiuBl51Zi9JiScRLb1R6B3HcenqTGLfIbYG5rPeHpRjYLCS
8TwonIESvOvoVUVZQVJ6XsqgRfDQOqv0sIHHYJOCm00+uhjMRFTA6pDXUb6u9NAfwtYX12AaIj2W
bkKyUlgxD0LL10l+vuqopqKHlAE4yPZNqAM2vliVRuvV2l9OMyhIMIOjhn6YdvgFGL3QEG+JU9p3
uhnhJaS9k5k3b0+cioZYIPQtG46CQbVHLIilrU63cs2yLhr8tIr6ZpsBGrwRemNZ9lpcYY0U8oC7
3kSlgve8ZtefwqsbhV/NL4NZW5Vzw7uLulr6tJO2sNc2ALcF0bHjnmsPaMWGxbDsafyzIXOEce3f
gu/tD/nheG9mWwC9/EdFnT12MwSmA7Qs2AhN/OTjK2BrXLOWrwiz8kHb/Zil1QOknNhEHXJU1DTC
uJAuzRd98YlQlJ2AWYJ9oPhe16K1yh2/MO/lN2ZX5sxDdLetI9+5xvgEUZ39kNArih09ajPgtm+4
EddwkMYzFxdYT7zaEIWg1iR90SFbCMMSA0q8YuKGAmOW2MAcnNU1FSnq1UWElNC0yTSvhx9P0/jp
LB+eVK+X5ZPnxThNZuwVGtPv4K8ouq0q5qzg70thBysuQzyYc54BYT+N79+KajDEwC5QjyCmTWa0
ucwcy729LUn3d3HW90gw4wIAUq2o+eCy787pEgmCSNZd1J3CZ2rjc/3TX4hcMA96KrY84owDpfO5
PzgKvZngyAcptQ5RgY8V+SaJB2Q7n527lHTyP9xUv4SRaxLO4FXgSC80Hy6cO+VTKOHH387fp6IJ
2qgPU5LNbVfzOmXlk4hZgfzBYBw65ilO2NNpa7ErV7A2touYmHrAwIqoMWK+7Qm538VmyZVc+ZdF
wNRkEXVzrCEne2X7M7b0Cl8MQKTjdC4gpwfUwZoEmfdUylakIyNmRPLKJAh46j5jViY8UJWHNiCm
YKTLbMW2yAxI4AbkzDTVKxNXGDZYEiiTMcZiYHPWLdSSIBQ0ZL8/UE+1gWm4zSGgFCwRrt3IPOYx
DHvtpKb99g9MGVFZ8qSZTpTsIJxXPXB0Z7oMbxXO/B4bD9cKd/ExAiCAYNuLyXsqET447eH8vuaE
0KjuaPI3+mfU2Ubsc+0xTCoeG5Ijyv3DdMMbXnGq/VglpMjw7NuEL3RQFoRcjN8cQ2fOWwzhetaI
jEll8L7gD1LVJ7BGyRjmiuqi/laSfr8mtsZkBOrF2PRokDmomQSv5HmmnqmRQqZTyx6At347VjAO
c+W62w6RShqIjFk2S9Pknu4Jvd0B5VXozzPUGgVl3yr9RtnfJ5PTSqKrO8QaMZlUcXpWpdxJiZFy
ahRvOeErd9ed6ubwtgTiXNYI7/H3CihQPKDPY/vF01KzKDbxbdQXPGzj7bABme6Ft/OqIOsQLrQ5
Bg/tCEKcBWsPJSYqg0Qe5BN8LpYKKl9FDYNCXWGb0jHM3VlxWpeU+4IO2hcdyK2EE3ToVYNZMYyR
1bUNmnSoKTxXDJUpbMj+tuCPworUQ109I41zm84P65ymnpG1S5DVFGX3cn4td2IAIch2HGInfcH9
WwOmVyYzBGSoRwdtbIYBh9DO2zRXOcApMGHM23zlDSd1r6dtXhZzQEVbVzu7jkjbVSH6lZEdfZIG
lR57fWIq88L+JzQg6oKij8anamb1ozjDr1rMXKc7/5GOktvMqFPd3AX5sNCahNh+FDY43afpY8nq
T8LKOdDKa/dqqIjWzc4kG299jYyc0CiVJSTBhmvlYM1uPBeut/XoehFDqmehaZW83lA47Eg5OfzJ
4EOvVjhBdX/wOdBhomScocy9Gf6+tYrYpYziem+xZnqj758O4KxKIwoC7+cuVydqELeYYkrLDBoW
PDr7Sp1Or8g4imspGRC6zexUbhnH6wihOF186gD0nDzGzLN+tZKj1uKmV6G1/9N2Ln0glX3HTsXC
lzn6+qdqCxKf2a5khhZkSGUC18AfoyFKlZi2EYtEcUh8yJaoPBlVZqUdGau4Cdsh0ogNMTiwXaA+
O4WqQxlFtLOY8UsvGyvuJnrsua3eifALSnFj4Y9sVKUjbvNPmv9T6dHYuXENxBIQjuKTD0zq4sNT
r1/ii+mtS6QY51wv5oXCYuv05WU5TpWe24QYvQLy0YeY5wFfjZ7reSC2uUnFr2GLTYjIUrWYGkLm
ihGaqP63s5QKFrhgarKrO611CnWdtcm9S/DU0NAcvmUOUeti/7TmUeIUAWWptoipD+UnKtH7K8Jq
kqGGxLno+KDQBT80yzouzNC91ZxMnQLHY7jh4DDAcbWThKROENkCc0f1YhmyfEcdmPHOv0x/y9jw
4mPDYTyIzdvNDZbBjeFoXfCI023dbT35vl2Cuj5QRpmrXU//y2DuRyR3z274IM8Skbde/G7EKhxb
OB/M1nBGczjSV9v5EXvNuz/fXCS3T6SjwYwjpvKBDVhr+TJGUfla7vGmszwXwCNub2zbblWXUhhF
HdOO+a/b3QFrmY3vnIrHC2afKyhZPiJ4LNQ1juNRhLDxeQD/rhh5gHH6/adrRJCv//iKBTOS6S16
NTYmigmiYOQPrsAadvocpNlNqelJxYKt8p8qL5oPOeINLBAe2+/TGY8DuzK9hLFU1LtNu5wNbefq
5MwD70FzvCIVwscb3kA+NutN9DLH3jwYKdh81ZFYzMIDRV8x75YUEKXoXvWe4Nlu7xG11Po+SS/l
eW8B9dgiBUuNMoVkjOiizgQ9bRaq8QeYWAUR3FTOBkJ7rlAFl82tFgCPuS0ZKJ3f2FVYPbpP1Gbh
RPs4iM8ZcY7HVCpDaCwe8wk3Vp45nF5Ww8aj44DN0CUdvIOWX4UBtBd4W5mjQRtNQ6MCtKpcfhnf
9I6GwyY7y0clA4WrZiy0ll+zuZfsJ0fM3rRdIKyc6xAVmcvVuc/72jEQ2nxocO2tg92TFjGt6Lrv
sOfbqeBHrKJTTyGiI/q8VoVUGw56VlMkBFAz47ae67hRzok3LhGsJNoSZNvBWoV1J3gK6qkFAdqI
8Zw6D1E1xWw9vAKwx0RG4EgNw6oUokxhP7GotLIhP4UHfT313vwwkDbBMTFloVBrK45kdpBDhpha
neahrMbbbkvVVv1jAlF3SqZsTtHp6mEOZVg0jeWz9mMEWHMCWBjWAzEeT7rJbpv28nRgY9S7zl5f
HFKBpGXJu3WFt0UQC3I1KpOOxRU++OTd/p/TT2+AcPTHx5zwuP6mN+yfAq9gIGjiCC2eO4EOjzte
XT1j7pqAzv9EMd96Hm58nQP/xQpzgj87948KewAUnM1H/fTlEj26yBUdFf0Qzv/gHHI0cOG/CuL4
27bWQxPtBSeGjw/YeYMQFbJ+WL/mUvuTqUUlKKCoVVyqnG2jWRVLDt2cWldPE+kn5Cm0eyx0r3Z6
/kwf4tQ7t/ROMDPaI5ELaFzKy8rekPPIJWpFIXE8+Px0ZQLBfqbwpZiiIZ5V+b3YODvA+yz+LZoe
cniPHVDfI7waeLkTqnv/P4T51S22cbwpvMyiYQmhXyGSyNV8sgXzIWzURWZEjDfMzqTb7WrbkdvC
pJMbYTGgL3rPtn5VFU1g8nQgPt9dG176MNIeRhiD60uAPyX3KxiPfcgZFIXIFomYv/rMCtRZLZWP
+A/5R5AOfFhhgFEA0cEBz+kmxoizYo3I4Cc0/dzFY9csY6GLyRMZ3CResGHnJotgE7uJuAIksTrg
YepVFjcIeHW8pJWRdJfLMrWQA1PXnvWAJ7+1TjfucXqPNs7M6w775Bxu9g8vrtnZKSSelzIUuSHq
T/JoPaT6xvXCUhZXUFVOmG5sV5j0UTCUKSUpJHRzwYfbZ6W8etuR6Wxnjl2bYZvs4zAtmjLvbkMY
IegN7XoeKVmV+MUKwWulzsKdUY2kFCGRQzPnZ6djFxFqqAwvqEojz6fl9UyRDQrMK/ip1WIj/nO4
Jvm8PM2NjUXdhzjPWbOdlecyo0DBJrsVNYUjpvTroZcPU/lJaxlrWV92TgKjl4r0HF9pjmf3QGIW
sFMV01/B4zDzS6rmQQxeyq5yhoTT9JLEmAzciNzsSyYND0+ROgm0WjuCJJXYWwPqNrnrYUV3FYWx
I+Q0bxFEly2pls0N+jBJ++R0tHMwDaMMYULxcIH/n56akkQK3Ibbuc0rPcBlr+WGFeBIWO3WIYPu
7fWW0nmsnN8g+vtvqjx05r2TKttb9/JY8z9JXQvKa5+YtrWBuADlLHZCpUcktlUjlGIAKvIss4B3
Iw1j8BYKlWHpFo/WYfAdUtcW7R4wOQNh9TwDQP3/17eYqQi43jHSagBWwVCxkcGOhn3iT3fpV6Xv
TOKyhtVYhfPaPNB/T8rInEXrc7YVw4SvnDTB1exuS5bq0jGNw+YLCSl4hIdf1aL2KmY+e9SGe9GB
xYH6wWytEqlQ8onThnRB0aB8VNWnszjZw0Sc5iatlUucASVCVvaV9Nd13/XHO/D1bEoe+rrcCNu1
hCEUqwGzrxaM2obnFWBuOjrMj5iKDQXohZmLrpdwZvNPy9rlp+43NKM433k9SgRhRrEgiI6mn2Q0
HQM8fJW8UDNRD08AasZggh0uNEfc2BNK71ELJwA53kgaWZRT6nd1+in4f+m+R3p74+iRdGH8pPX0
rC60F6EMLXgPBRXK+65UqUMo/cqhYbYaqgffRJ66ekztYUS+P2tk0202pRTMQ3pCv0sWIZve+uy3
Wqksja8WG0O3/R4UxkC8A8mF/d9cmfMZNsonk/sELRv/5ycEUXuqzq1VuBKfoforPBBVQ+xRMwbB
wXWMJeaE93yAXvIhKh3J1wPVJ+tKIMoL3OZi+CSYXE3cwb6yMM7QxPI9Yt5qqRC9deFAeubcbsgs
no9IOAL969aiJqRIiBGBeXQrH2HMm8GTYMrAXTwx3oQTml1EchXHUh06zjYiwmKYsFCB/zcEqqZ0
CsSD6fOIWJB3RSHBS9/Yz0Lo3NWgoRcsI7Q0OmtPmtrBiZcZbg1SHnsYOaUWC5XNj8tiV6RI0sEP
LHvbi1widCIhAUbLN1bJezyiIvMSWpbCaKATmSexYyK4n9Dd9X26XyKz9Bo4tE63dHi7vENgjQ8A
tdYo7PjqESwQDWB7PociQB9zaw72fwdl1jNkt1bnUHVXqkRoXP/nT7civBvsytJhOnvJHbdMx5JV
9pjtdXBuBNoq1soIapYIWyygIL5vKsEZeNwVsRA08UTTzMZ/rUX7mltBdAGyurGrjTK12a8dJPT8
ZSx7EByYGqVYf4H0Q8cBe2Y2TwfNeBleDJ6tqC0cd7J/x+71n3gCWwAu243e0eqQ3G2//QK5J65k
4uZ/xXv27gj1zS+BOE66sPiOL2IjzRb8L3F769peObLWwTZowdCl2Ej+IXjOGZn2mOZuIFKLACuL
F9oPTTvVBE1BJOfcNix7ERYoGTLzKzYjLXF1ExJwni6BRjHtrUrxCzhVcid6WZjQ6UJfVvy6XaZ+
JWCfNAaCvR8VhCEYjRq/NTBx2v1sqaidBcnnuXBjNJBCUv4+jPswWASDPeufo6zCJVlS54e/aM2j
GdGNMsfSBsU/TOVG6KxoO53kVtC83XQIEJrb6B1J2AXpnDAnRAapvJ6F3upAygvnElGSePdNW0Rr
sxkPAi8sfVeMGa+SdaUyze75FPFCsxZzL3E6INvztXzdc7KKHC12hLkESMdgtGT+jlrV+A2uVIbg
5t6Rf1Y+e5liflcCWpaGh7yCYp7+NRZn9lHDbdhjS66q4tgveX5qK4Tt9IxVYd2CNmwOhE+yZ6R4
0cLzZNRhQXPFjTCswUmX0XhI4qJXn/VlK4rXbDNlS3mdtjeNhmwQ291h3hh9tF26zCxS9UnSe0pv
yrgzrAOhf4c31BSKYlYuWwNqauY26Z9cj9D1bjgmSwVu7laNg/LkbpWF+AOvYjJ4wp49N8XiWDre
TETOn7rjDkufb7/itRT6gU4NIkL2TtWe3f4Dy+u8ov3CasabvC3U601zdQ3jKDHfVxVqEANsEgFc
e6AdNIEErxfe+ZCJQXnJLKPbV7D9aSjtLgxAJjEa8czdbPqukH3Pq/NTy3O+DVmHfW3GomGcV5R8
HkGieAVeObI7tgGCX9FN1OoX6USrMNSnlCnbkWrnapuV9qEVkdW/qr5pbWntdB4C1wQo4pm+b6h4
+ef45LZy8DIImp/kK5DO8kRXpxHmiVTIcf5mor4Gmu/Gs9TDeSI4js3n0A5u08yZaJNPlQGGN2V7
i8q+Lpm42y36FUCxMbMK7Tw83roFo3810jekauag619SeEE33jHSif8zB1qcM7Z8Y2drd+ohvnto
/2+ofTRFTXNkS2KfQOoMAC82bFsFWezm540I7sFwyxGepu9eg5MRjiEVFGu96LkK5qb3ReLcYEyw
+PuBYbuxWfve+FHvZjiJe7LvYSwEU9V52HrgyWQKqHuz7NO/THhMBiavTamSDu9syin2YqjnqsVp
y6NCJ7FpmQDvIilcw11UTS7D3x8Dw5oG8G+sdU0O8NfXXvy7BOsmuLXmHgFixTbcfhf+0AHOXBj7
biUYHhCE7B453pC6A0bHs9PTuF2lU2RMus9T3ZRBz3X7k/8Zc9dF/ez+aoOQJi7DNvipygyP+JgX
gdzu9Gc1qO7igc9Wn01n5FpWZ2/GSkHSe8S60lTHizwr6RNPIDSvI0MKdlY9gUAa+smfWgWQOfXi
lP5vLm0JiUSBE3vL20irqNfw7jhAeQ0tE8CptSHiCQPJkcYWAHv4nt9JWRAuzy6/E7W02KBSvKLL
hYvgwQntpczrkTe1GNLaZqP1JGbf5Gzm/FxNdXYqFqE53fsTHHBU4mNNtY68HgCWE2+88R3YxKN4
yi+JQVmt5yBGqYULwl4xcPFfdsdHKrQvY5Im4QSYtd5h7IplUfu+9WXaPtVAfwsFGOK5NPpYriH2
aJ8QdC3lZGi2QibW3UjgdaT/YB/q3u1WXrQfBSfIB43/YwUuRmhTgGs+FAx2Y0XI0wglE5muSpIP
uzzrR8lZ0kKjjzeoRhucxKDG3mcCRCg1Ks9CQv5VSzkx8650cj1HBhXx1+vDKUpLsi+I97ba2qhG
VLSYnqxJGhynOMnXlbWV4jUuKKc53zdFuvz/NHWnv+qJYWKR0bK23ZHXh0sM2w19HSD5or63aZHd
T/iaDUUY0b19Rwl0ZKb5VtN5ZYjJWTjDXa0f1aIPN+oaWauIrYmbCfRnaVgPT8/mFLBDL9rsSOMC
V1sJMrPt/zeTwYKj7dxpZrGBqSSz3HEEuADaypOe3eL74VP/g+BCEvtRlUW4EJMs0qQMGY9+AOEJ
Act4bFXIurPJjB0lWL/i0UiqUS14jPoCr9Z1R0hm86fh/nKfdHNhsA20f46D1wPzn8lXFtPedAB4
69ZpDhei52nODbhhEmUqMRquSxFKIf1h8+WSDvWB4orTUrzveXxD7/5MFFMwC44b9IQiV3KgdFnJ
TTjZaQwK04kkeYNaQQKehqxav9XqyXYUOM+XRGcfsnG6vfwGAvL7P5PnpDVnF1FhEF0eSTgLoOZw
75w/E0sDKGNjeAro+nl+uICcvwShEeuK4QdXdPwOUs9pLQcZIiVwQvG+YxRV68tnFbK3LX4g/zXj
Be+seCoX1Abwi3OEZXyiFZLN4XLnZt0n6pFlDsca6OZm/pUHKH01c94PBYSXGascpmWxJpBeECUi
YCuYUy38209WQGPqteLKEr+K+7T19Uk+EsmaLwob/HB4HsaMiH0Sl7B/B6M8O8JbvW9pgObOpCLn
rUpInhq67Y2C7v43o3LBetcme7oO2c0yE4yG+jxHGr4vq0OzoJN6nkgCWEZa9PSGEhpw7aKOMhpI
/bMg9Dqc3yAZ1YPEkXNoQGRAn0qRbp0oHsveb6Tq77SSxTk+ZxdtjbqfPszMjPc++18pYUN6c+QM
eArcZUIaB1YFZVEEVMqjpV7tnEbOVlUh+82qx4qc963IdQKbl5qFiV52Ztd7W89sRxAKhZGUQ3/b
c5nqwYHRQ28QEVkIf4GvL1yLiyItZNJz2lVmvuhSKfpEG6AgRVTBo/v/kzR5uffrgCe/+o21hlmg
/egNMNiTdTLyoYQldVTk7ryU8A7WtVZaOOqfLhN+BQwEx14aPtOCWriRiNLqL16K7dpoKKPW2FUE
6IDcqqFq2C5bREtNwuSm1qVtsplCKIJQaADachUK8FZCMQ7gh+I+bmrSCHU9EYxh6aYhpN3zaqLo
O5kNhrRYIFyhmcTO2ZPIMRZ0nw7HFh/8N/q3aEiYL0BwWRcUNFDRV8ld4wETmmRgJ5VYgkKwvVGt
eKahl5VqpGbwA0hXWqDOYNEMiOrJbo08jaTH73Oi+Ml45T41Ia3wforMqol1NMF+oMTdebMMjF+e
Z8dVWWGgWRAYUBKQDoI6QUKtntIMrGnBrecKpIbnbhsyY74VKwJmfwR28eb0vmjyEvXoS4vPNQWB
EkvaEnJ0NXNHyL+G1rRLyZxIbeVkRET6khKSoTkxsX+FT1CEI5gboQ/QTpdZp9BSaLZz1WmM64zB
V2VpguvZ+gWwNeGE6mKzNEOXcTq3d8jJGDf0CDUValgiGkVal3+9m0wmZKlqxUbWuvKU7u4QI5Ws
fO4lbDJIYnlJ39Adkm9ow8f/mUs4gS+iUTQs/xdIN7pMuyrjuVFWN6q4pH8KaNqw07D212lFfpwn
1viihsbk+tyuedrUu6hOIqE04UIiIZN/kx5lG6YMn6LtLn0oMNuyPQ9FpqCC+fKGFhXQaJMZzyDz
lD7RZr6wna4ABSHOUmfTgfUBcVrmE23oP2Z0ehRF4pJvTfJtIJaf+xslR34eittPTZIP0X7bdO2W
HYQW0SSjcqNtoggdsxzpMv1HgONHvkQVvIedF0PakHtyQ1FQUY7JvofqxBni2KBTczE33LRL1Oid
TBRKd3v54so8S2D1FGB5BxQcXEXdmE8sQGEfoJWNgo5dLadp2xfZ0g/wq/XN/ammVv1XM0FB2Tl5
TliPFhcM4kw3aTVrlsdOjOkNs0wReffOuTGC8c8DGizlBOWTkOUvYg7e9G8nzQ6Iqbr2yS7f6zwI
czYzQhwEgBpbX9YLfdo6cXnri8A67C8mBZc9ztgDCbCXqT4LsEaABKLPjBXhb8w9ID1SXi7+S/9S
vKKAX9khhQpWTmZRs5KJl6Hmlm9E3NlK0IiRBwhY62ZxAnunaF2mH0S/GLnM8H3uMfGb/OmL7ZdT
M0VPn69IN2/b9OyqLPT083ZG6s4ir321nrG8H0uSGlBYgsXJygjaTxBQhcaAr9NAo7RhZZRGKuFn
CY+fcgC98BzI7ctQCy52RQhC+rU19zv4YnLHqmhWp2FOZ4ErkU60Iyy6T2+6b65JXsEb4cq3kiDi
dFpZzqOTv3V2DcCmymsvnU8tbC+Rk2JrAASfRJ5PSkiHRT4O8IZ30xd5oAc5pSfdn/wMLEGBdDND
FLuJPXBtVTf9y9EH6PdX6iQ2tpSL4FphZaXWNnNvowXjumarN2Vjmfo3eNQwQ89U4nzT1xpTuFPk
L3OOgYRq/XL22Eei2ZiAbJImIh4TBAVoNhSecGlM57x+G/QpFKBZ9l4dX6Iy6GkIf6TewnwjodqL
7EJsUzi7chaja25manzkC6UuwhtVi/baqTmYJnJZ2EZV/W0uUpNu2qrEcrHMd9LcM+smKy0r6NIO
sxdC7Q5PmD6Wi3zZLEo7ExZ79KfR7GmszSvhnOACMnSsRWAaAixkY/dKgZbJeUgRgu+PkWHiJziX
t+ayMWVce4SJp+gdf0prQ9q4vFm364qlzxuBciv1AWT7NMxHoYuz69h8yDacIiNKFvuBUKtr0zgc
f7A1Xzht1pTxlm085QtJc7rn4AgXP6Qd+Cdnd14Cjbkis49cNX0SqjT2PLOJHlnITOmJ9ZnktB2I
Sau7eYRAH3AfBmJU9uybsEQgEZ5m1ZEAF7WQyqAhNrVk6QlrFOdtldIF2Kf5t3YKtNAEv1iAi2Mt
k62yHrJ0xCdyXqiRSrbWcbFW2iDSjT7eylfXApFphmw9Uc88kMRAP0Kws86nD3mt2r+BtXhosHLD
SoFI6uphlcXiuTfMLAXOfdDVf1VeXtK9O3U09yqgIdNJj9IwlsJuSsDojmU66bNA3eIxFVkht+Th
2zH3EIO0ND71lRkwGELAXS7abuq8qIqPQ1+xpTXzS8fVno/ZKgidbpxV827yx0DC1ZAcLgtsT9bY
Fl6BgJq8cENY5ZWIiDLFLagr5ZSRVr/9jS92yVzC4J+44vG0YjPconxyNv77WKJAk8w5l/6WKgNy
LhX0aedLYatfnzHo+fWwTRR+ko1OqoroPVQfVNXIPDi7tpeBAHpnr46aKar0eu0gbsMGbla3Ce+0
zKZWiHnUh8SkiFwDQUjMPvGqA85I0OXSjgaKu/lRmV2NhHRpt8XhAo8Z3hF6ZtUJ7OJh1A/3T0UJ
Amb9dM1VUwQUbOP/79cnLjjGtKb4W+1kv+el3JCis61e3WV1GiY5/XcOR4YM7nvja+PdOqleyK9h
D7S5TLjaP44M2lpjh/tv91sBens8LhmEnBwW8JhdZHBMqc7Mrt3uNZAYRXl4lgINnOjTgQgDlPh2
alOEgHsqvRkVxXd9TZvMloBB1b0E/8HDqpw/++RWHAvaGEN347md2B/qk0CCWSsjkcJgvytoHBNp
pGvzmJM3JfWmGHOE/AUu4N5dO+znr0G4bEdhozPrcq4fAMTcyuT+5Q4VKc5JFnBdGf7JZt/c850V
waOfKFxXkg3thjKcpoGEXbgxJOk9LkL3Y0K7e+TdkV/qVGxe8jZaqcEc5+cH/4fCGeUPTqiBEisH
tmA5kVrOilpqvmGQGySCaIwln20Kvy0mJa0re3mmVxlVIIZxjuFJs90sTJfy9iub3FrbM9gX1eY3
yhhioBCtXAnDNOMRJ/t1hoL/9rtjfBVlYUC/aZan7ty5m5wpS14Y+4JbNN2i9AxHqsyO4ANPBYZU
tkFNld4+687XKvmBXqPkXxB7yzpAvEfFWYQLvVOQOrR5mt9TbrfmdKTnFO1EvyC6TnkIoqsOtsrv
odp4uba0jp/khlvhLYrhacPi68w0xojo2nHw8kuhuHwKvy1EOGycQmfn7U7zREZ6fhJbRys2eeTg
Fr4jLRb8EJxJX+IBqmD63kc/h7tldVy8wi5ZV8r3MplGtXRyv2gyRJQAcufbkuwi4uyeiMri2zXy
YK3TXUGd8zQFOX0W5W3lHOBUEucqa0K9VKwiqa/1b2DjaFQh0DNoP3XOUxKdAYQf+Acwu8VdrnI0
DBk+rkcsPOdw2WxTxeAQGkfq5QQ0dH4cEeABMrF5gMv+idG2dZx/DgvLKdnd9GJMkSyso0uuAirW
tZrd1J8e/YyO9dLo37NR8e7RE8kkIw7yEOLCbDoOGiwK8WPRTdTzx3DLhViaUOMUICvJtnoTJ7ZS
mMJH2h/BtdpV0Pj2A0ZW8dFmDlAVNmmwcrF5UbzkT+Px/nUtLSc+IFrB9gWsinEKTZpCc6P3TN3j
aSHG2jCPndmn1uRT8JZQiR7ZmuuzA/HBfaOhk0XNu++OAJ5dnpq3Qrig+XHGMHnbvv389ZqaYFdM
weQF7XGLbUvwo4qU+ZiVO7+blUI7ZpsHjwIxQeYY6bFnN91NC8XJfH/bEgdJWQqeui82XpoILlIa
K2PA/IXsjIFxXfS53xZoNVgoLlEnfyFfnp/1A09sKnw/9XI9HpDnV8BSpzLzxQwkjBISVOdsAIw5
JG8ZnOaXua2yY5HEgQdK9AKkP6LFazFxc7QZ7ZVDekLakeDYFeFSKB2GoLVEsV8F/NMtcsPdd784
rAmVLYHmNpOhwR5ui0m0LXpP8B9kEzc8mVOBXF5CtXX6z3SNPK1ZbgewPod7Axx9V1S3C7PyOl7A
4wDuJAda6ClN0YV2yWFv8Sy4O8hYaeJ4Ex1OPFXu20zD5xWyfRfS6nDJfkBMMotpBy23zsAOORKb
XGOBrQXxmOnVrUbynuWGmBJ2+mZWgdGaDX2ZrmCDYla8wv9SRARXBG9upOBlf5Nubs7Gap0yo7hG
lcOyAPXOcwMnv/Zp3sAPCheEhiRbXZemTSfKnLwaZ4PIIdk5HYfKPeOigjvEJh3YLL/1itaudryz
o9349+X9u1w3WaXM8K7zOvdXZ4b/+cDCJCAG1Gf4r2pOHpW0Ju/wquhwnWo7nU4HiII7GtRLI76O
wWHzCUNY4segsRqIrs57JOECwzbXSNp5xzoby/9odTgQCMPKSYF9eg5l5e6EiVVfZ4s5S+8hcZrX
srhgdpQZoZd6eaBfmphL3dS1HHUbfYrZZsy62adzmj7QmCzYoagJUPsRxKXy+5+BsnKH2qC44cuZ
zpDbGDXRDbK+KHWxKA2isbFx01rZC1MCru6g5R5E51LCOFbz6yja2OGGEr3uQUqaZ7S6yIEMcjaL
tQsW0xIsSSaNDI97n93N+Jj96hvZ6zv0zssqgHXx+yJ/vIS+RO2CcneIPCX0XjeuzRLJAwtk/DoC
i9BJ1zhWnsqm5WPU0YqXjVEoGxwvZ4NYv+p9Q6xrdlom0Bq9XQB5RhVuCMf5ZWo9kQYQVWwUBXaA
1OCb2WJn+csxTa8+9DYrZ5iXSN6sBZE+kyHTnS8BLt53S3tuq3jtE/oxpo+5S5Z0TiieeHhL6XXg
B9a4Y8V2OtHeFna+gAl86qj9JM+TT5DjkamDqbgzMc8e6UJuwisRZo5z2MVgmgmYEwQlPYR8oHso
eMyeTIFKu/+r4ZmZEqQz/AWzk9XIvKyl8698naji3DQc5sqjA80k96AmuZDkPdEzWQ+pOIGaHPGQ
FTHShYB+lsyyG65ea7NqAqiZWV58nJbVCn/WeJ3UrrOl9cVYzqCP39jYH2GqTRzvcTbknIpxDJgZ
Kz673nH1ccuwlK7fEFnfn+JKSig3mXOhoOMVZZ1dehaN0OZWWnt8yrTKuBz4+7IMhVHlAZDtrj+x
+9C8ukHyb0Ppv2BZCP9hpsjlQDDa0+6meXwOJrRR947BZcCu+JiCf6ntqFZ2Vz40DyAXINEfms+p
ze91mLQVr+XQce1ueA8u+L3Y5OU2Eka2oDoW2feDqSApk+nyHC16Qd2w8VRFq334wl6vBh0RiT1Y
r2SZFga3vh1gGynIX/xJtQ5XGseKNpFy1u8GVmgg5gdCwUFHXoLpynUbGO5OV/iW+Q9uO3qBuFxP
TU79S8TZNvIglc8n5p7GuYqIox6U56PWLqQXmCamD1nhJ/M3QXA6YdeOVBnANf1tZdiQ+lhUB508
x9xqEZnQ3j9dpR9SigAbgJBXkHF8P6pDDwKVBe5gIptRbC9U7x07LrfWtwIskSc1vS8kneqtGKFH
siQCL+BNQfGzbaTqjR1gNMMoKtHXFqVkVF1Uq6gDL9Qj3p5q8aDhV0RfUgh80Iyn0aDXK+AF3edx
wixM6lyNxr7mDtNhAztJbBPOL2GcFh/gkf8GWot/mtUdGTOOeJAbg/VyAZaWF8x9GSIPxqIaUehU
AjdMpdscKiJv4mF5I86ayiwUXwfnDC8msbREZyZyrr71sffZRok3Y8faRCnaT3PGXZR79RnHIMol
8XylVAYX4n0n5JmTJzPAxdOK3p9hhvDPJT+gYkFkCTzgh9nVRfMf762ojAYwQ6rm6O9MJ1YMHyVG
ndqCohYfDWsPaZcsNdUGLEMtw7vY4GHgopMuvmczxCr2+chYz9r7xQmj9z/NZedYuSuejZC2LiqE
H64lDi5zkiV5D3EdzeqQyK40bwA1Ibm//XgoV+I1QlNZG5/57AtBB5MsFbTeNi+jLvIOdQkKHCl3
Z1FltRjd45Q8CPIatxUBvZSizeEWP+bpSUC1WGJYOp3GZLnhmsusyb1MkYKBe/nPUsVmylkARpLS
JMkhElDIM+8k84OkVD7StOgGr4tcZh148yOX1L7gjVr2oRffcsdFcjsV0wJT0gL5noRzk4vkF7qo
zRG/kVTCqBagPtyEbCHr2bXhHRG3Myp8rDC7LpuTSdT1Ii1CtLrxCSqa8XJ9+lpz0NFwRQGWHVwq
TLZbajqCZl5PZrIigPZ/DTLGEQ75d4ceCMYzMaehps4kFr4jqmK+rt7z1IiTloOc1BAc8MRB+4NA
PL5lEgOd+SvAbmYqtx2eLpDZi97tJiVooX3yC4k2S+vw5rugl+B2uAIrZMjqSsoWXkM1eQdB7NbW
gXpNhjzNXdRgVMsu88tV+0rhCd+wN3et10NLZwQYdKJBilqe3VqMl8AFr8axBJr5ldzO2LDSKVGK
DwSwkdLsXucqbY8UtDrTojoNU3CEnn0QjmUffQuWPAaqsGPjk8RrBnL90/GfcW0mM9WWWNVuSXtt
QSpNIEa+O/ecc1nyUZkiALg4Xa9yYGEBeknOEw/agsO4oFiVxYb2WRh6lmfBGooURTZNaD+esnXX
mdB0S3zty4rkqGJjHqPbRpPcFDolW20Zr8ppkZAZexvPpw8tczMgAz3MpTF6GTURcFMyxReP/kCE
zM2mi0ZVIxcXaHXcqsJNPkrv/MBz5td0lcP9aIUcTVh97Z3tZyN1hZL+56KdGuEvvv0McWzkPN4J
pKulyllAlqZLXtLDLqiEY0dU+ZmoCdKy6NWavQWI9sCYwpMnNInJ8KLO+JJV4CakWF4B6Iwi2GTu
rqzBzaXM/9nA0vTxlFJqovl1bAU3xUY/xdnSRQAsQgf2fjuZk4Ii5bGtiYV7WzQ7rv6W0flc7zV5
nyyvtDpwseB2As1UDwztnv4mw4Hg8mO7e3YEqzXZxMzqjVyeQ5B0oBIvp6tft2tZK20itDZTVxb6
XLdnQvfQTr9zK0o9z2U9vnUC2ZrKPeuZBoLkmavSZyqD1Zrm3amIIc78/k1TMK9bjAeX3Rogd44h
pQPdlnKZLZqFk9SNPuGWd719J9T3FmBcXDdaX9m1YKf3TgsCOBCUTPx49WxmqrG1gDjJ2fvvgCuk
gxuLKIPXl/aHOeS2yMU2Vy7C5py497uko5SQ+P0sxZnE+rQiuJQHlRpqQsgo/q7rV5dcciOBeu7D
Byh7Sph0Q79S1T+ne3OU4+wkfCAX/tD1ifameL2xtEuAAFHq5B6PVgsK44YoLdo873Pz3HzYVVAG
3CGBo3Ea4BbYXmUdM0h1RgatlccnMGncSmLh0TrSQ4I9b6Z45rHG4+82EVGfhHOsiMKoHY41vbLO
ydN/QvSzGRCjxFpEExZhgxtBmAP4aAnJ6161j9NrZUzy7FT2DqxuZRcUA98pyqhWnRmFxqlo7VxF
PJDPR2qvnb5Vc7LZ84MywVZ4R/vXPdoHEYU0jeq7DFnk49fMKqJsDWbZP21SqzjdMi2DXJFt7Rsj
aK+MUAgSZ+l4FSv1Wy/sk4iiCyAqFKPPtYZYANMsiqmZGfSLqvkuySgAwxYkr4QTPaLL+Xj7XGuF
RsWlC3Clcn10wYH11Mh4DPxchaEf/1ldHbfNguaKCAKZ6hpB+MFxa0bz5Jz+ecFuQFFobRzr3sYi
KniRjKHoYWckugx8E3hF3Xkdcb0gzjgKCqH+bb1KdTCaWTTuMafjwPMEROHeIF1hrswgtaAB8aNf
bbx3ziqVtUT8C3nZs4moZ+ddFupgGJYIQFkYvAbfeMxwt0SvWUMuLlITtLkhIyetJ6V0xtJ3wLK3
zvLwq5c+Lps3QocqYwKxYo/kVq0KfCEzYmsrSYGrceuIa+iByuzWQ2Twb3nY1uMYlpUf+VEkpArA
6T+3HJtXUKTboYqZw9Gok1FjfWK2JYaB1utCE3ZGdIwnxucRdyHHSuYMq0+ef83amv0SZDKSGyV9
wVLkvuA6eTPgXGMusVTirJnemXjC/OO63S1YMjkRQfEqlevYOkC/3BfeLjQdNBMeyxHctq6b7QcZ
36luWg7bw/uYIELJ26OXzN4N8TjpXQSYESPtmDHJoaGrkwbdZ/rKsP3iihn6mDPa1jx9uB2QlcB8
OcIItYYXE/bdkRl42rjYZBrMLLhMtOXbo7yKuTZhF8Dm/UM/k0icssIAPSUVY9RHMEx/d8vIlWgc
gDgo+p7AwKAJ2YdavT90+b/DSdoqgEitMQV+NG9jEj+FRGE4PB5xDShqj+U5AOKYX0nvKFgDfHql
fyEU5bJBIlLtNarn+0gk01i9jNSlL/KMDOWpjyuifwRXveZIyiRuBh6dVW4i9rLoEKji6MBG1TZf
AIaWl8Ct1cqwtZ9eXaMPxePDL6rp5rUaQ5T2cpDCt4/S56A6IZy0IdzfVOivbrNqsdidk2Fisxoz
PkzprPblTZCVMxQ4gKMymQGQxyUDoujgv4ng5CVwsZqcF6XR5wognvicyy5wWmzPOf1f8sNqp4rB
MftsIaGoEl9Ia3wUoLZROySAPp0GzzxZhZF+gJoD9eqDPWOrqj3x0X7tK1tJw/EJIzB9gE1xHj+8
qAhg4JogyL7n01N0GTPb3hPf+2V8mqNlqwu44cKStYUKyilSeGjNrJfWTufGfY446XkZ6Liq7aDT
sl2yX79RUzh9KFtgnIpTvhH2Lzq/M42mxQJvaQ5VSwwcKRFUIfjkX9rd1VUYAj3SLv8eUJcq9vjw
zKvuYH9i5nBujkdDajYYVRp7xVvDFC+WXFVBx+ltSo6ADQaRmuDTm4GnKSQ/RiLy1RZjoKHp9Gsa
I+GM/gz7/+81E2u1C/UbsZte5YwHQ0eM4UgCdq7LVvgku0cVZHedzzHgYIwF6/tCorY/kIY+IGpi
PTtDHLGcB9OctPvX5XRifIQGG+BST+7UrEKcrHb4z08PlOMzLb5ira3b6EVw38PhiVLxMHWHT3MX
J4CdI1y1adPsuprkpyXwoPPH9iugfwNrRfPparj2+ukdix6ROnZkJjjUCUrQ0fV7AZJhhc6B0FJ5
ePidG31Dej0vPllMX6RUZtdpJ4juZvnNCk32EqkXP2bNqGsqbTg/Q5c9oZIQj3wA8zGOnrWIdTs4
4VRWxcRkNfTkA0imVfogsloUDQnyDsoj6IOM/b1P0QqfI7jN/Xz61iDTq94JBgJktANzd/zO2ZLr
ZghLZfFh0REmG+owkWPRP2h/GMSzWFlAb2NtvYL5rreT3v9cduVC8dGNriysVne4POiMi1aclo2V
faslsMrNTt5f+LotegWoH0h7vGWIDjtIwQb1vilxIppWbHoJqGcENR8rl6IHsX423XHGPBoctHWU
32pFD/r2vmyDytpMpJ0xQxTUet+thuDBdQ63u/7t4lG1afAglvparMI9v7aFg/jWu7tU4rOzYUk3
KGeoMutvHUtUprnSDyHfabrd08m6+UMj1bTRQDLiS5DR5BP6gbRrP4+94Y5/g+alncHdTqCrk5jG
15sppJwlbuwYJdvBxMZHwtChyAlvYeyLAVS8AkTnTiyxBkex6SalIeKFL0EVb3te1wKMv6F0lEHs
rnxr304OhEi1WAMI06MJg6OpbPf4wIP6kWD2v7K2AtRLQ0O5mV4vJ5FhBDD6TTxR+PN/RGSr2lkr
wT6g3X597qi8LFM4LRv3GKrAaDUi8KgG0u6yXIDkH/yTyAI6rDwPDdY66fZRPoIHIcQdnZZpmEX2
W+TXwNvokJlYiUv+yKlyQ7pYzUjcLUaxrWuMs71j0PQ98neVu0THoA+Lmqn+qho+q8ANCneVOTfG
vytW0L6nDcrhEYP5twZNTFPclNKFIDeaFcVnM4twfj/yAWUc2oS/jLcPbrZ7cCwwrvGvkB254rYv
dMFosrUP+h+qNCtyQm+0ezZjha0bYzbGyWp7pBMwE4QcW/gb2cmOypewY8C+4GaBSkl5YTmA6cCf
ptac6elrtL+GYjsI7kFZH5zNsaIPfJSxM90deK7o7qilCY1pYiZU8KRj6ZdxUckx4Mv9j194vFzs
g61P5IvVxtpnf+z4+baRp36GOvLFRr3lwpa2GUWA2fe+hnFqYr3Rl5gYqCigf46bzLQwy0ep2mdD
KfjaTJTwYQ50FuX/G/I3pWFzQ/Loi76KQ3/A6wP2akPYXAi/lMQdsCXX9xGdqMU66Ly87erP2bGj
icTwP9rDD0RdIkKRlY7ydt6dmRE2PUYR5Oji+kEY7zAHPFj8bWFflpNxkX+DXmPAvC+NOY/Q1WGL
pkfSAfpSpC3tFxkfIXQncJgmPJrEoTEE+Gr0cO9UwqrW5Py+Jo5vvl2Na0ZdQKZ42/nnflZwi6wW
wcyP8zFaDPopCwJcgq+z+uXxmMjSe8Q21q2ab02IuE2UTJsvZoEmsFjXmAwvWSIiisbrcGiMncUw
dxclD0CfAZrIc1nkvbfz8kbtq9MTo7q1/fihdYss7IT82XM8T53M+Oy/ZpAyqwklJT9+IQZw8uKk
0E2bL/XeOskjMKUPUnXSol1KYhsZCoW7W9pm8+vp19qgeMClMbwYlORmcdfxDLQTbCv+Ayf1RCqT
zSI/3uRy+5n017WQRv+zf4b7tj/sZZmDwuGXp/HLXUS8UeFvkFRLJ/WYq6/ouNgPoZtM4tD7Awjo
obvLGQkNF9KoWppb95HPyHB5u79UmalUnHwHyruZIqfVU+PuCNfEESQIXQH8y1WyWZGkq8X03eb3
UzYsEL3d3fiWwG/RSyCNVRGiXGBNYRnAJWwYRCbdnnadpx++ZNIv4c/gu3iwf0MclaWvqAr6D3F+
zx+CU2jyvaB1o1ypafd4ZBnCUMijhoPh3lt+JoHbNiVz0mqp5IjmzoMcfNJRGUFaQYCzvGnk4SBR
P8nO4vbErwwNs60U5yREpLbekY6xTwsqDphx9mNDreMuc/cFtY15o8zAL0cja6DgiBJphIUaOAe3
I9Qb4EBZZdEXdj1TqDUmCvpqOHsxqROZEjGO49DOFwS7iYxC+jE4nwfNON1iWLww+TXLK1Q4vgL8
FeUdxeVOS8ykQ/c+nN7xcMa3KEHftNrNv96qsjMMrplbP5q9wUYvQa6R3BCRIHgI/G1mxkmexuoZ
iSf0b8eLVMYv2cEO7f736VOz73E490/vOdmr3v0Jf1ApjeKE42BIc0Alj8o1WVz8SmTUrP2p/rSw
nhBdQktjRshMH3Yw3Kaw/B+DT1Pr71matbW4GCf9FngutDzKH+MPGw9YIiYEGHSdScUGezj6Ovx/
XSCVRFoIkOQDHcDpARYHRWQ/pMJdFbUxHB93Cjon3fcmplUJDw/99k8G9KIe0X++LUWYfGy0PXyW
glZqda8ZPZzXrOXDlaIRGZGnsmUmE4zYaUcNGlrKqWWl6BelTRPLtG+KUqyGEcbHTxzSlL7ocQg6
8oc6zSKRUX32h3fwvpzXwEjj6d4mg4GzQKjO8d9VqZAAyWGLpPVmiGooX4o3K9PrfXWKPdq0f5OQ
016wbaPMyTo1PBMCWPLNjxIh7Qb8Lx1apgeC2qT8O47cptPA+rD0py8CXg1MnJtHpyIp7mMC25gm
N0AoNN3JH//RKInH7C+MBHM8tzjN1rXgjAAI4ZKfXVBNmXuCDCfQKoSRZsViEk5e4tj5JcPf+1pn
OhlKzlJ+9/5PwGGc61txATIW+85pd1bbRPUB+6yXGjffXyRtSagxcX5HoIKx87eCZRODDPdsn52B
+yrs3BLc2cBzXRaFP5H+oAqegTcCqePwmSBVlsMe2PQEfJdA9IpOgd3MYMMZArbKG8rWE5YA6wD6
YDUOU/M526DstEMKR98Hdt6xeQcj7XNQUGijOPq2Q2IAWyALTpU0W8mbzaLyVu6T6R7t7Sy3++t+
I8ukoAur6axq+TmCyS9hmvsraTl4XV7iv++LwjA7gcvib2plrtoTxzSofWQtP7Tz1hEyk1zlurIr
nGWMD2Q52B6qTV1CPg+lfn62jeltFKYGtz6oaFH/LtSDEY7xFThj4dmJHu6vbr+Szo8sWN0dI+SN
UWLqLLNNmjsuwbnDYd7RGEwSf2+gg9nqN/MWw+7CnqdBy5fYqxYW4r32/2UItw+WOiS0wImTooGV
d/FTTZ/QhCFQHugItkiqERZSrNi6yJB3bMJeF/PDqY9gBBN5fn+8vvMuaJvCoKyvvyPUlwc+QHn0
zKd1ujdzm7nfm9MXMHyuebueOzhdbbdx6zllDBnFxO4rOfmw/NluBRxFyFcky3TxK+3SvDpkjPJl
h0zImzm8Li4OM/14C+4v9liUMLtaCL1f+jVLzL5J23ufN2c1zTBmx7PIYpaq1qAt7SKORKdMdwBo
BKwMdC7YltS2Wwo5Lxsae3KHlE/RsDjSW1htSzXQHMhXKQn2qPtG4rNO4s9s9ANEdrSTVrC6APVX
Ola4ajEx9w/NqZ7erzzrZC/VUdsaaDlvA1YohrfU4Zws0VBaGGCTsssgrrO+d3lvQTqDh+EvsWNP
uiCjio+xtouFr6N1+1Ssp+zmAgsh0DY1LgEGDQzIvftGYC/nWa7+DOWG0VoSP8+A8ivOFJVFBOb2
Tw9I8bfZcbdtgLPN6JqyXjMdgr49q8fNMGnH3lM+ctK9qWAR63zdUHSMF1mZ8EXvlut8J36hvdOA
YvnKDAjVe00CRILF7Et/RbO1QYJnptT0/fWVp/41rlpGVTfZN7exdI++kGgNsG9ptG019MF6JXB3
REfGE/l4HIeayTFgVlixcN6W46K5mcXesQ21CUbE2N4adU0HGFN8igS/0+H9i7trPqNX5Sesnzsa
Xu+kG8ChmbgmFME6INMBthGeYscI2AJCFrtTIguTFDZNwng2GIp5f/fVtYz0XudXUWKmiAUfS0a0
vU5JMXl0ZuM50QoOv2LSblb7JwwJyKrEUv9LGPsHbiuS57sWr3OlRXfh4nT5ZljRrxpYLnWhzpEE
E3qDLXgr2VA2BreMEq+hZE+kChRi66TLTn/PrpdFPNHU2Wkt5m/mP7CadIJVQarSjY6t4hag8iSD
VnNzOg4oLZDx0smBxdvsb/y9qa6eqWKAI7wJf9y7JgOuEIU+1X2tSe39Lxay9qxvLmmuC0GWsdfn
uLb7/K/kS6meRINX2uPJGov51SDfQsUXvp6GNQWmOSWuLCRMJM67CqUPpDqqhZrzViVHbwT/v4Xf
8G1eoLkIgfAvd9Brr344A7nhTXZ8gbxmaTV2a+i9BBKKLGybX5U3994VD+i/xVROkbrKyRnhDiRC
A8Z7St3RvbfsMAN/8Yk3T+b0sJu3fpr92UGLLasYzYgzVX7GY/IzZF2liiqLwz/lk8PaachI3yR3
gBgpPqy0TV3synJo+o4SUgSqgEaz0Xt3466eRHR3RcLSUOTTX1RGA5mDWP2paNyt6cVA7vtpyMAl
nLyCS8n4ytdvicJhTsksbmYlh8v8erFbT1KcFJ+we0FHRf5DX9w7dJDhy4AE2JpgxaoEiQtGmzmn
WOXXt61LGefYdBXOJCXiez6qRwc35qNXTP9yNY3Z2JLew+RFG3ympXdeAMVm2eT8p/52KusQOyF+
clFPHQVVePNGrQVJerM/ad/ID5tB7c9D1p2+tjvKoIRFwkvLn4aP0vYqQG5xYK09FzZvPjL0Krpm
TYZ8KmtQ6l1mPnvG3mVQGyg7W6sYIuwHCBbugD82dJunrqKfZ97lBl4pLgCJwX0v3w7ZmObnytpP
CuUYQCRJEER4fdDxkp6neIxExigP1Yv79aKmIv8So2iq5o/iA52I/agUHWpSthHgHF98ADZe0VUc
C5OdBLxKW115IjCOExanHmvxkuS/CAsxMeb2bFVWQCOhM+ni2PEV7W3WhkuQ4W3UOM2YC6qejNz4
N30pNI/sjcoVnEs7nXa4i8yHVPqlFEcggcXoIstymrzSEkx0TH5sSU3IDr2YO0vl95dbSs1bLKr9
/ei4VHVQ6/0EGDag8uDBo3pqTjZo6oRDnWG3W6jHBE2crTtOMIkcF7RZ8HBgR/WWjeaGJ0Og5d8R
TyMf6qjUkbyyXZstqwQI22sWbLfeLNqdMSY/QBKt7CKMhB+Ib20u9E/xSbj+AxtFOcQF3bIXZTx6
9v25raUYBaewSvIXc0cz+MwhKM9cHnJpv5I7M0ZAm9QTXZw+GGb/e0DE1sojclLX+rMl5oAZIhbx
D9OG2zFQLQLHHe8v6U/bubFS1ea7eO6Pv7+hBoEi9k4Cnkyyf8psLxp0yzY5xN5HBXhKAdx31R62
w4t7DI5j/i1xqlrxxRe7eugO77NxzqXgZriPrz18zFRSIHSd4Q9/FZ3dvh9oz45YCIdOhFUOXnBC
r8yYWndscfCpCUYjvxZIVWrKmw8vBQf4CmxnP95+kPJ4mi1nL5TCRfS0ztb2yQNXTtrH/1wogt69
QqGYVIKUEteFy0IYzJ0O6AI5cLjVbXwfifznkMN5ucqtQ0sGYFVUbZRWj5LRkVsNZKIN+j4+7MZj
UNCEEwvG/TbSclEU5sF9fN+ihd6acNVRbKGiW8ak2hrjnWMBxqrtBK7fm6kga6GZQoTqlatpX2B0
1mzSdOuQVIT0BCzkuTELn4lRyjGRHQrredmZRc8UV+BtyLXbj/XTsPBzoPpMbqU3CZbb2YzY9vEp
wzmMnequqZiHjGrQVvWJ0zjNI6QM8iVcETRu+RavTrsNLq6+0s0ZMEdcxq+z29t4D5/jdLyPmyXQ
7Rps6R+I1r6tF0GOrslmvDSIh5UHtwPThZDY2shvJIrF9l9R0utIziuTMHWydScQvSim0LTFm6wf
gtzcOike4UPYeKCLoivYIXq2Av7WSXfn4LQPikbCoaPe74zgIMyn+X8t8ZnGPaKhQFzpfjwAEZwt
WlZNa1/UvWGx3Kdi6x36CFxg4B+qQWThgi22pO3snnNFUf1brswnUHhK6hna3dCAkKa0uguwPVzk
xjxnWuuATJgmQ7tT25Tu9UL+bptzI1JQnyd6FzRBDSuaLkjJq3ggLXHKzn9yDC5+0D/Y5BfcGIk7
7tmjZFiXRdvnMlSyJnAJJbm0dguY/H+ZnB4nf1LRM7AWlFNaWUJ7iCdppbCLjlfHYmWl3z8rTFaU
6whA+FxHnTYmdf80pZGxhv3Pf2O39NhZUxD2Vun+8SWvcJyg8Aop6NM8377OpotnYjrA+Jfm3phN
BeZflQd5nGp+akNFAXOHDC0Xd3ZFCFcOP6O4YfeLxtXjomqR72yoeflYnIR9umJri7cPMDlK4lid
/8lk32z7TVxdLv1qwllcH5DZX4skJjr9+ofoqxWMwnYFq7yFrImufEol7w4hadUebYazf9feem18
cv4FSiLNe6NIX7+cj0KJZgfNgg38Fa4FQCGeqei2qHlyL/vUIjquQfO/oZPcW04Rw9uqIGGxp2O9
iHFsatgokqeR/AfaKkUToqlRmYXET+Ff7/zlU/xa3pp6Qrh3krjMOnPAbqfe0pesYQMccNbSYDFo
bIHtjus4qBhVTTLFI3YMf8Gf+dRHIKxrK91hwTIjb5BKYgmhU337RqAF28ARUfcZjeLEMdt4zee0
IALrn2Qd+PCgydj2Jca/aMcFn0q+/ojbFmBarQi5TTZybm+MCkSYAaoW9By48JlYZzxsCf2fKkI1
ppLAWsrf5CkWOESPX5WkSDIMVVQluRCPwrx0TcNxh+0hkMcujbAUboE3lzdD1BJyMTBkQQXk/8aJ
7+Go7ocwYk1wMPQivjp6A1rLb82E9xf5SYgzCkCDKDooGAtkUvAYkFtEJyO/TZ1RIlWN7qndFUIp
XynMD4+XlEgyqa3je2czjw/7mU1S85PMjrxhkOi30BKkkrtVI7VJjtmpNY/R9vwc5etcQAO2kLvh
GDN+JAgnYTtrdq7D9yaIIbJzJwNO5Bgadfj2tw5FwlIvGvKXFWstBXDABzvkVy+MFVf9Fij5sU0Q
kEldQdrxU75Z83DFOJpdbIsq2EG8GtWIP06clDtkGK/is5ahX6+EZgaie0WxkABZOj8oI/93PwWG
mEPvlTO2HzWdOw94uQuVj2YJwp/x1y2GUp6AdrOYU4MANSC9JIvohmSf6zio6u/mEUht+hDAej8/
Q/TvWKKE/Mf4/STb0SCOE2gcONVe87Cve6Ps2EgycdLMx3X+ivCAchiKFv0cZ+ywAb/qAlxXpWln
uaPysod2S9bXmakNl5vwVf7haH65LpJnVbuvcmskAaxYKKxtw+b6Pt6cqXxMFoyEdtnCAxn7yJaV
3ZIFSgpGQVkPaRlAu+YL6SGbFZpAMjPcOd7FP6CT+OCE6cuok+vZajwTkcMatBxS77Qs+n28sTut
bvW55ICzcgaJtXzd4nVgngA2I2fHHqO/cBzdv74immVzfUw6wkL0ZO1jm/WYoYNSTgP3NtR8qu8s
arZB7IZGib4PcM1zy5cmwc6ZFPu+G05fUp557Aa8DJcTzZ8lFXsM9oiDvTmaD+5VQon0f44VgpCY
htyBTsw3iSP+5M9WUezGdce+6eXLB8mSuITcoTYJ/qZm/Cl9lifggJi3Tb/qJHGcZWocT3KeUP1P
aHNQ2rDvwvuuZQImBT1DDaRd6/0Vb389Hlj8qrS/ftOWswPkqzsVijCBOW2FxL2GLi8+iaZnZPb6
DD/5f+xCe6UQsaLKcmB1wPEECwaTIrFf2fTH/Ofe3iJNt9ibpz+nLAed2rdP1rbm5dCXEmNef+70
P++j9q7i5Tjxe4Z2VcCBTqNsNSjrv+zFrz9zItPaGTJquvKfCQI2oaxbSprcy9e5xOpUfLjY3ldl
sL3BWTU50JiPlzkqdh+qsI6hLJcz4IKSejvCoQWgpYNQLBUmYhHGXLPYTWfEwurv+8u97q5bwpdu
FYYYhB6TV8wPFjbtpHvYRQ4yDjFlRRK9GNaJatuQGdj4LMPvAq+61EgA+Ld94wONxMLdm/RF2080
OCgyCNPpLbOx56iUkdl2h9InB/dz4l3+IZOnUSCexOArWwrbxk4Rs2StpVkiL9S4qCXcZ95FQ+dQ
nJPuFVzsqg224bQRItxD93XZ4XKR1NbK1bNEDkqeo74XfXcPk7tS10Ut9f+u0zyP+zk1ppVSRbSF
pliafYa1pMVpkr3b5mHKNV/jnugiLSO1KHprMoO4eVMvI3iXcbOC+Iue/r3f8nNJQtWI2mSCUBce
noGEIKswOsMsvjfp5lS0nETw1/zfcb+pgCkht1X5hW2JNwGQS620kH1JRedQgOl+D2w8aQjX35oL
MkJ9AQ6zdlLrTM37MwXI7k5pRsZy/8JKDTw1KXAKtOtUVPJQhHa5qLHssRm5l+kxIYbNkJ9DImz1
FdfP418k7+/2MIdFDWeZ/7+Dm/nmR4+JsAuj9Z6ka4rbKzSBKsTGNSfgMwiolax1NS88bAVy22e4
x3l4oaJtCyJAzzNj98A01M2MVXuX+MOBbfGqEtV9D6qwjZWy9hKFsrqEiGfiGm489kP5+nOrrjMJ
+W0pUcfDhAdE2OGLX/tJ+tL3rPIiyd5/bubyN6pd29b0KAGdiLV8nppR8ETqUgIg02oi8dLywAeT
HsT9KEvYsKvFFzw7KEB6PggVD/PWySQWgYMXiWBc6TQ9uttuoshBKtTEQo0eCyrrAqplUhbpbtE/
O73Z6ajNLB0ZcG2OfYBMF44r8MFvi2XPAx5I8ZkYTLAErR7p1xLlMUw8h+VYPUQ6HUiuXA01gm55
1YjYrV57p8W2VVVvCO4gkINPwUbed2CaTa5UogQM4vnwbFDUi4jKyfZuWqAWGPZY75G0dlPtSTQr
Jd+aRKo/h7B1ngFTbistvLFu6V7uc5eHJN+73FKDwKRYTYogjPQf0zF6/6D3wHkLz7r7P3uQyUc7
dsn617k89SSPifeLOkALpzk62YzcL94MsbSc13rVJhHu9H1gorr7duvKkLDD0cuadaUGiy2LMK6Y
dm0z/F2l9dWJOpiTlDDNcxpo7usckGxnSHHHHr88loJP+/vrZvrMNmMZZCUl/smr0Vodq5n7gYym
h/0BYF2P/Nh7+SR6rkPPqpZzAlhyTKdKrZwchBpQ+4fMlJhyO+odO3o2JmSjHnPWr9Ch1vReVp1x
2SPFxU7Vci9NqEVhl8Er4M8Qe4m4I4gsKA0mcEq7w75s7TPkOOclGBammMgGbeDQmbCcCah/CyVH
AtIr2v2Nf/I9qw3GvS5Ma1trmN0mtyupyt2sr36pINZ1E0Pb4GFmAiRBv3ZmVLukTf43U/vwDpwB
IKsP936lmZjeOoekU7ceq+L3svfGX/7uQ9NmHBQBeSgpEizu1bs01xWSe64HB20dzQPQBY7w0i6w
vomlmJ42/iEh9rPjhFhA1TqhVfNkGmA3itpEbqcfXzHZx3VTRr1Sk63zPzQwrFg++xuRaVyJztIX
tTO7S4P9RtMMQGkTpZ+kfAs3f8JeX6gvYqPDHtwiwkywvTRZON8x9DSI9II+AiRleJrx5JkbEKoS
OOas+/jIE/ZlQ4FZS9JAqkGsKEyV6wb/EmqM21CpyZHTz5SR/J1ahWv4d6Oqe1kvXME40kEscNbi
fDl7i10HJC+Fk7lMybrWaxdlcDByIW27kpjpfZum0YKSet30/xIlinr7CtxAojXXTEYScUsnd/nw
sxQmb2uAJD7J+Wiu7ETqg0CKbxfnbgH9tROjgM/bR3o2LtJrZRulz7t73jEaLro7rR/S9qIvLFEo
jqvaKYwwK0sV3ojnJokZrjqUy6pAHe8ey8FO1sk5KxJVHeM+DLDEBXv9ifrhFQkWQ575WJ8F2L5g
W+NikbmXgM38UpuPk1tISIUPE90H47vBF2Nj4LlEBG7wvhf5nDt6M7GSotVpLvFZv3XV70WBMlhx
kOEymP8EqqqXs0vBsA/ejmpLY+i1nxHvfevpAX0N9fAPYRlMw52agVv+dbAUiMezocrkzfmE0aMj
I5Vm68bKS+6zc9sQ0jxZDf2rKxq+HqfcX/A8AYW8mUIRMJKEU0Bdyb6ogr6ryQlHai4QUmXZIbV3
JfcVZIE/SbLcVkfWIFYNjk4oR6D8FFRQLTTZI5ra1k5+Y9WqWKgtq0cEb7agS0Wgeum8IA5s27pA
1PoShJGaYzZgcWzRQdMjJOAUE75KsuCelgJrd7ESVP+cRly6BUDOvh39JASrcJ7n6qadRlmw6zby
jIUDNTuCIf9dkCDK6PtxIdExXVViPCvWkKJk8HnQascgn0BE3Mx8BjXtSECKo6BV4euYHDZktpBw
Hr/Zod2sOv6z6TJzS/CkzpLxF6uM7lQisNglicX/J5XOI1oxkTfbK45s14rAHpfjh0Nuwo7zjsXI
wPJXL43MKAFaJV1jv+qHx3azU8XhkZqoBIbfS5ipNxRewfgqJU93sAlf2NI5410gPgSb8Gz07BmU
rfdZhWVA48MdsWnOgGvsPGComE0BDZBLzqnnJEnKJnv63R0T1yiIe0PDhxCQNJcFol1Rcf52/KGj
DOxr22U+ycM8rln6b6NLPbeIJpVYIUKV+HgjhRRcGgmWjYX7bPe1hiuqWpT+1Bp3mt9JG3h5+SRZ
Jxt3pldc0TQbsfXPg0bjFvmkIU1thENk3/HmiR6+Dn8vTPyHPJOcNANeC1ZfeIqeL69Zqw1ve/ga
C6UoB9p5BdSp/V/7Oa73VTZk0PG1tImsfzQwQZOqlrgfCifvx+CJKL/wCMUmdiV0hYZXoixLoTo1
j8ymQTG+20NfMEXBXhY/IbHch3rRWH4DW+ulzAh8SrGYkGFG7J+A7qUg8l9/vp4+7kY9G4Vt1GdI
j0t1MEsQrW+7Aho1S1ONHkWFtEMhSrlqjgT6fO/ArkoYUmGAJpbaQQgce/2cIx2LBF8mWJtdIA43
FhjEvbwDe3cE8YQY5akAiiLioiCxoS9MaVIFgnKKYEYJq9fvHorhfk+ROC2hvMZ6GvDZ6FAJO0MI
toWQaDGR1G0OQYcP5E1BQly4+7ma3ZJdT0K6nU2XF2rTmClfcImHzUYTRcJgXqlGkdL17DDuwV/x
NGd/KKulOKQ2v9MaQ2NrDMVlcmmHPm0d4y8i8OhFq+YIQ1EUgwhAFt5HraErElTXUeeCyZw+bZKI
hXtrR7AM9ZEOfwNzKJhV+ILJgrswlJtN+TZs54mTmZdo3kAKMX0s45Bosc5z0yCta3AnnA7JU0gZ
rWmzqeG7fqAfUyfJG/+OrA8RjRYu5UhjmiLeiI4SCmbWiafMnN2lYXbkycTBpEBaJNON9vdAh/bc
I4kFD9G1FA+Ql5np7wJOEsE5U+DfHHlzZTBTBLyQGxDUhJCd7vdHn5uGYAFuom3mWh8JvLAyfpoK
xbWtYq47yAv/igZK4cb0BcasonO3ufnkbTfvQkIt5ccqWzm7JrPUCI1eeaNDWG0IJPLrCT2jYrgz
vtNmWOJkVfLVyn6sBi8NaWxf79CE21FudG82pFwFXaSHFXDdW2PkGo3tGpLIedAwkquBmf9l30nK
RJPV+cnPd4gzzBJa2iDm7JkxKeesNW6V/N2tO8II8G0AYWJNcs2MvW+cdQCcqjz2wqnmGVspZR0r
4jwSd48IKnz1lrBHP207ODJ8rHvV8GV6w6Rb7gmQO45tZEM1dqlYxQ5FDv3p4uEU6NapHwwQKt9k
TOC3rghOBerVLu4tMkYlkTibeCvBMUpcP6ttcX3K7s5f5g6rgCVEXBqRV2PNxC6uc1oISAhVl0V3
FLhEkcGIvq3ll8XHQv4dzSX8Qd5+ouUCYJRPdVtt8ksGk7f03zzISaO+3q9PKp8BuODp8JX9e3h1
KatILYRlAjxHrfcjoYuYjfxwmvAJ2jXCLyqSVGorABODGcUe5TqPGofhlBTKUrFZdZTQxAYWyTKS
+LHVX/mxGzVEdxAxNYFRdT7T+sBQedkQIfwv7WCIrosWSAD1jJJ9WioU9nnceZUysiFd6tQan4cG
ZQO8nApWp/1wa1fqzpVsXlP8g/R9k0IJfnpJD5B6FmckqHgAnzIdEfqc9gE9hgiz2lSuUA6t6zKA
udp7VE7zwDbLomAh5bUpI48NhyEYNtb7cC83Z3RlE+0GKkkwIDVTErt5YVv1KfqPcjPvco8TuJIE
KjWW1BfFeJVthsc4i8vTsd3BVJ5fUjXHvOIJJclPnY+dMdnNYDfYjdtWpA3IPOtjNtEiPi6iSFV6
YKcehBR8M2sNeyy3DLYHcNX5IxgZp9bSEJctkiPRR3TEJ5lgsTWaWIUsOHaRszf9MdzqMIuVZbF9
BCZqr0wxlGQAgkjNyqeMPVAAGj/esQDV7LkeeuKxta9nwJPckUSwYCEHVHgoiHeltE/2ZauKBekt
J9lU7En0oCgGnEcjD3K+pKJ1pseVvL3jOthMiRG+r+H3dpWQdSqhNM3jmWWiJmwxB5KgSyJy6gyg
/3hR9kCLkxPoXVKITt1mdgUz5k5PTpFDWnbn6FKD7SZhvxDjnRm88KBAe39T01X9kr7UtOL0WXPo
xK/rtFUAg+v4Nz/jgFTNN2AasmPASsZN1V9Qx1yRDycp/rIB79wARFOcxHtipvH3h80z2n0qxdyH
9Q7GiI66yuS3mNkNFFj41Yr8vs5EFXJU3kvKhumm0pCjroCxwhNtgPjENPsDDgI9CT0uN2v7WApl
vzKyUmRXnokyOLWPeAPJvyWaC8sgnvGgpJFCsSKkQeFE0CxiihQZQvIAbnA9bS6XDdNms0rDIX53
a/9/ZGMt2+eTlV84xOKm+VeDpkJ3P1PhfVOigpuwKK9B1HC03OxxcTdcL+a4VcWizOh7edtmiG7C
5ocgX6MMQ/XxxjX5Uhj5XJg1GHPad18cP/Sx3t+Ox2F5ASKy52WgPkVPKzJY1l5ocDwkNv6vSs7o
qCUQjO6mhvTygdSUdJxJeXqXuK8S7HicSGCpnLT8LOyNAGJgza5+hCPI2qlD0rpLh/CRdDylCnB/
DQdnyU8bHizcFZbixMEZnNS60ZMlAbDKefyhFrh30zHn2Fbj+b+E0uMyowfSxBKbWf3uo0NGJs5k
igSx52vObVl8uHa7rJv/0fVKMEQd9K3KJc72kVmwCMpvMEtqUOpjBkP7UHfPVQyrVvv0+SdjK6ET
AtlilaBRAeRdNABC6PEblOuNNijFUT13r5EOiG5qpdN3lAvLeUYlWq5VDEE9/+wWSzl50cBq6zyW
gs2QqVJX3OMYFhWaI11Vn9yAWSJHLLEjSlg0y08Tznhv+WJTaT/PXgmB45EpseJtVdesekcrSlTJ
K2hZkADIchHuLA1EraGHGTBU2++0FEP/NXEZeRYa5qVtPApnTQbBwoLQzeA1bmprhjSqOpD5ZRmg
dClEbdkqiN87r19gFEVEDboTxciafC/6JauTNCEl2GuoHOWpCIm/05oqVWpQvYI4hVn6zfQ678Sc
M62/1AKyOU1BdZi8XYdkdhJGUh6H+KZvYbTMnH4EnGRT/kK8aDa56/0/h0+5B6+3FFFzSsFnbwjC
DvQcEv3xSyVijMJbEPQ0URs1oaiXa/oliW0wWDdSu9O0hs1kYVH2kU2DQqxet4lYhI5GezJV2n7r
i9FdFM+HXEqUPkSG1h4Yu1V5+Fxs4M+siEe1jk7DmrrpDplYDHVoQzSqrsFdwZF93aND8Xbmuxpp
rCuW7/ah1BksXi3UinSLnO5hKdjLbYSGcyCS1b+Qgx3QoGqd1X+atbnFTN2pkWsNGIT/Psxame8I
Q9LHumT5JQhhGRKN/+Bm4lzxTdrscy0K5JbWOJzFJMNQg29jx5tOHSJPj2K/OvZRgpK/p1FcwcCu
to+HWc76heH+TTVZ84UncwowRPMgx44y3qabkgwCJosQ/1a09YFYyTZ+zzhTWtCE7H47hZjC9fc8
2XyB+2EGxZzuBPqRooxUEGJLBMpDSUeM9taok6BhhTzxx4sWGR9IkL6X3ANbTunpbsISSg06R+UH
ATpm79EqeCjGo9j68aSXa+VF/6mPZF5OqlUFB5InaMaFLmd3dhe+pdyN9RPkyVl79VtFOwiyniVu
J7SaRk8B2HjtK1Vg+lPYoMAkjsHnLt84kVK+z7TAd8c5iLcGIT03HCd54suciGTUGpHxrrNe08YC
5wp2bZnvAzxmx6FVkVViwgXr0u7V56TqG0astJt9dhQhF4lZ7LuBDfmhA93bf7xuQHIkoDDoKtCX
VRiecg3wvw/eVUKeuLa/VA7aUlHESul2y6Z1dUmts/NQ0oo97Ra9tNPWamIGIMGs6+vNI5qvialx
8d9Tu8fMKk5siWINm61FiDMwTD2W1zlaPBBJNu8hmlISfxjYER45B5fm+2yZE6mvarpQMdzqifn8
5uBKa/cvkvYcR5Oa5QG/ww0teofhU4OOrv4wum3SGcNnB4isMSIv/Oj4ElwIVPLSvz2+b++A4suj
5f+dtwX/KGm3wLfLoRMrVJ2na5mLNh2t+1GCuR4KFsQmu2IVZEBsTrS2nbMV1Ths7is4Hoot4iAS
bVgZ9YOR6UA8vhSE58FdJD7bA64+bUivuCivlkiG2q+XUXLleOGa8wt4nuHx3nOkyHUvdBJrYXJg
NVXpyMFg5kaNjNXA3r07Z2VAswAEKY0hyYlXgXr8PhV2ZrWps9c9GPnVoJr3aiH+dDC3/1n99bEy
lsKtxZsV8xD6nTQsI1+WJC6+O4s20TgkhhaaRiVrOFfy8QH/V1dbpcXpNgejeztyeHSkxu4S/D5/
6wpUoDrs0ZyTfROV1vKs+RB6i3rC1SYHM0cs8smaAaK9gRJfxY49CwoYh+pQO44p/DMb3ENU/RAg
y26kvoJgJP7yRdaWesMvMlZZKgVwvhIjpBTw7ruCGZdOklsyda5FL4bNCGK5+S8+E7KhS8X+ApFT
r1iHGtMgVyLB91ozVJ2sBIpf+XlC7DTutRlH6n5m6xdiffMvqnh5VXqz1BZYvDWrks+tUGQpMC9T
lra1HK6kId27t/o6Zm6C+pLRXINPpMIdK1+gs1ZRenikNFtMCgb1jpeilcUBlDYvfL1D0G4CBkGJ
XRceW12NH32sRGHNEw/D40IOZuGhYq3+a62PnlFSS+VbOPV3r2sMkVk4PWk24vjEbhPsAJuU9/LF
7YwQRVEIjGbhrdECivfeUubsdHHWI5lhu2LuZkoOA89wJtGtVUzkfqQoZly0WjGidK880BuaX6i2
vBAdK8aS91Qu5Vqd4nDNuMmq9IgSV7xGpczQ+WHIOs1xKoayK8ajiCTzEEK11xV1iwV75glM+2XB
FU2upxmjeuYeqi2+/5/RQX/3nCS7kfAVSLDpLzP6y3AQ6fZ7jtbFlqA0hVqmEN/KUQuiotr8vl+z
yAgLrkLxZWD5h/ZLYS1S2rYejb9w7q+0Sm3cRwisKdQs+HmdB4p9lhGqR8D9dVRkjSq6vJQK3uVN
7LNgzlih5i+a8epV99S9vN7yVOjefYFYzq7KivsbMr7eo306/FAtrGn9cSErwO/wAroL/QpGGnxy
v3OzfvCdRTiafcorkZypwEtZ4+GxvqaVgGDJXd2iNAQNQ7mqHulVKkXfaL9TbqhVy9ZnJKOSaes+
IW1SaTG+8tVj2tyoxiY+0ScLCPYQadxTBbAjv4z4WxA6mhDNeQVA5KcSLHXPYU0AfyAI9OgNiGe7
5eekV2HQ75Nx4Xhe514ABbtAuWqpgb/nx71fHrtDaAoPalP3Hw5/2ungdEcrSxyt2N3FZiSznNk0
b/zr1weSLdk8/22MQPOk4QkgRQ2zUYIfuJ5Jvn1BoDDTsLGZvP4q/W9yh3OHkanSQaUMgmcsdP/Z
JRszTgqIU8UAX3fG//if72ZakXJTLnvNGwb6A9FrRIi4ot4LmBlJtOOuSayavklYsO9p5atIbAmS
4LF2YQAISl1h5qJ+XdPuKHJdwogVaLtctGcQJ5DyX8huh5K5BIdGIoe0BXeFG5bPFIB3QAtLtPcA
pHX36SQkrz0+EB4HBkm1w61SK7eEWHE7Q/2hcUUVnN+kTtYCcGGrkkvDwuFL7bVF8tYYQtfwBXol
W3wGlUV7kz0uBDfH43PB2k79U6nS+4Ag073Qcxrz7mFyF/6nxvcFE/lDNoi8nQKSr/Zs3avMfWVR
a4iNLf/8xvGE0DWwMiusoxMwvAvLs1UsY5DYbwuEPK81922WAedw+4o0tWV+YgNQzKY9BPD5Krip
vaT3do0OXIqS/psnGZVtf8YKJ/IYkuY+coUmgECHqvKnLHbuqF99g1bxmkCeAiLDQcAOcsGoCL1o
wlxG93j3lm2Ms+GjcDqVsScOfxR0C+VzAILTUfujh0x/1jyrhNRZswkumhW1JEotDVrRPcs2hxYB
0C5Y1GYoQaoW0dmZUVe2qe1seaYAiety+Gw1hc7fQxu5j8S5zIQZez3GQYokSkP1dbALxOezPVf7
HHp8a6X32RxVajtAIeic/NUaquO2XLRLluRCr0eU9t9VdukFcx5j2yA2eatguxuhAjEwCrvQSvUr
jnoWlzJ6lsL32jZSMgZTdWjB6QQtM+4B2aXaO/7TE4kyMg5Kclu0y3Op1/ZmTp4ZOmdaLIzyR2zt
DJkYXmtVsxFZuERTvk5WClHC/JPubQ9KxJCHXgfxrnShel1qC1qi0HMA/dE8ujX04aT5kFdrxZ9y
X5wVzOpb5Ut10bdLqUb442jvhC81109Pexbsua8ugc+k3j9sed5nGx9+kTjCscJtvORa9LoP0EnW
4qECuUSEGIfj580qt/KpyZ4S3j0WUXNpSgCPULvNreoB9pQzzQbXF0EdfJR+l1eZfMS80EKtkAzv
2XwgLYJ7mf1lt/VyYrCY1w0Jl36Rp+wTVgKpnpEgYLd3UX2YnLiMDK3ktajkTGTpWDM1QYjcuyCe
QtAK7RTCJsHE4edx3LlNecBsXou3Nam9UgkcKf1sRhFlUZV7+QSXoY/ga6MnZLNGxMqy28b8jLFe
qFE3UN0ZvsVeYIrhKSoS/EIR7v1sHMFuHUV6JskulgXYXzEnjKpPaX5ZMzOqoHBZzW4dynHmutx8
7MhARsQrU19idHnTQiD9hBwmfVTaUzorxkegCHNBpuTX1fXhUG6iATTtXW9TXsIJP7/x8dCb6ezg
ULRPWVrAwELDl951uVV6VoZTF8kqAFnE65z2wm5MGtWmsAq6t3BIpAD0YgwRA9AJJF88/IeMJzZd
76GXK223WQYjWAyrZPFjXap16sVhvst4uJFJW/ou6UNuQvufltLylhQOTAi1LRxZfXsMDcE/Io1D
XL2V4C3SK4CmLnsvRHwn059yLqCjKmAC1QGdMPjowPW24U198yiFfsjIVSyLYGgDvUjqUC237ZYO
FCnI2wVVhfV6HZL5UgsZ5arBp4Q++dk4SCYW9Ke3zHPhPhrOH5UZ24NP5i9R+6lCuWeKCXpssB1t
b1IIa4XimD3EuJEHITSxB2iFowXKRHXlcuq5rem4ELISBegwXm07HnjpB85ZWbE3lvNQm6QgS+cB
ejdFQBBx72N52YGO3rB19YhqGNCw3oKLysd0HVScuUzBNb9JOvi9WR1kKre9POjJrv/4d4JO/U2b
vqN4lkfugpHJuwXtAsb4Emlpn7fXD749L+AXZUY1Mv2IOYczEs/sxXJezDUByGdp/JNkD6wfe3Ut
/0nZqSEHytTr+VA6woznuCwoaffKbj3SS4jMzGm/vb1HRO0/0cJeeMSBFh/qpIKNBvedure0VpRH
LVPsWElqCnRKNAo+xu0SEHs4NFwJxecA+RS4BFSwerEPcCBVsPlfMJFABQu5cj+pnR8Pq2ztc2WQ
ixdidjNYWJSjDaHBjDOnmKPrv5m6ZkFekDgnq+24iqH467yyyOg+5703yoCQLAzko10J/y/ATdsS
dg2Xyy3umQHSSTh7wCO5AMBLa/TD1FYYtJjmQ8M5GMSn1Y0TsuDfzM76uA56pPa4S3NcusW9zQG4
qIw/SOy/Kg5BGZP7vNiBO0CH1tKB/jUuXFsUQOddAZGcu4h0abyyxYuCc5c7bTZv2K5wdyeaVjS4
Z7eguqs5Bzb6Yw2d0akgfG3MzT/cE/bCA1h+MuVI+/uyNv3JW/a1Ph6eX2Cvrc51WcdVu36PMHa/
IvSQo3r+4Ewy/pX9dBPTl8OEWTf1jrZbJp/CpNCqMhwBSV69QggcomgtrAWRWoAOzlf3gtsZCzTA
wttqqab8rLNUJ3wsif8AkiH6E5kANJMVjr1bp0SwEAHLyLhh9zL+RvpBtjuzayyXjdm0Jq1LFRFM
Y+jrlb47d23PkYlLNTR0BmS0RA6B3YDVHEb0X5XXRK/1IzQInyrcT0+/dI2SHX9/RQgPax0mxTgN
XJMHj2gY+ubGCjayvS27ngC+FMv0s8+EXaSgKppSSdwTR/Gc0YG/6BEvAslnyeeiyaDjL+A+i/Kv
X8CJiAU7Tc/7H9kpIbhtZsV8eh4oUjhsMxygQVN9GSdWjWX/M+39O+uc3p7ycy6QLeCt3VupjcB3
KTHlVNTcLTiepqbTm1+4drOec9e3W/OzbZnKjuPuivWXI0OAmskMskVvz+zLpw2vYYvKEJxUvo70
ElFJW6zgcKA/fX46y/wY8pW2U4/u5pLiGi3b4TIyaGCFUtb/I9A3VHDlztM5fKXRCx2fZO+2prmm
vf5LZffd1SX8XR3vYPlds7r8JF40pmAhEcx/44WT81fKiqYa1yJtFlCAX+1Y5bLzGp/uj/owGVpx
TVq64t9x4tREYwQr2oXdmn6vJL6yfir8/EROJlnXaqi66x+D6ENhil54Q+RH3S9tcteMvSzD66Us
MOrddb/L0Vy5wRLmNqFcluQGTEZcfNL6psvsyWfzjqace4tGUcg3f91UffOW9rQQQNDeU+Mo5MKY
datvLUKtjbNyObiUJFKw+NebJETR9Pi/N3XwEp2T8DwhoWY2e5AAFZiL1LAyQ4gWoF7+j38EuNk8
zG1p2nElXeRc61UVtpY8c1Mfl/QQ1bdY37fxRvjZud90FpoZBYyMEEFQRgz6MwRoGHQMldEHmK5P
KzFAFxLgBvZDTGphUEHV2ayX/6wvQ6OeHTp0wcHp9/614Wm8Pi1fa51PDtaIMCJ0WHzyaO0+4Fv6
lDjTE/RyAoAjfXSaa4yeX+jiOmRA12MYHW5zBcPhfSKngNyHVCzgQb00uWyx4vrF9lKO44LVXw35
mnJKPaaL6HSl1L47TjyJUhrvyem5avARLPBI70tRqJEcX7O+06JJsmh120ZgOx6wSdXQjXn7RzT0
qjgHpw+Qb7ONdUXp85C4nGuj2FJ57a4wNnsc0XA79LDBVogTJE88F7WzeDaFRDP3cWKP3F1Qib1Z
KS3DVxU4rBSU4DS+7hZBmByEuAFjmkXYeD7HDoMCDEM9b+NOCDHDz/4fpV0E06/qnwEY2jeS2jGV
Dn5jG30N9Zw/Nxx5l2VhmBYS1+5xNbYb1AFBnb3IZdDX7W6rVD83U9kAMuyyuwDXAqLCkkVBQwLB
WUbgmnjbX37+7wcAcX0sN153p62GaSdCe+pTSwlD6Us8Qu6JYGc7oTl11EmaXagM5d0dmnfq/7Ue
DxykQnM7KLXerrWVlCJdo+bo0e8mvgbIRX51yTvFq8T+vo1LEI8qV0KkrlHUIiPTCj2YgNQtfvR7
TE9DnzEefIToClVz7ZJbrQK3ZBWCaxGHkl5cuQAho4btWSLgS59hJ2oNup9xROOvLWtvfO6t6IpE
8nkIPUtAAfkW0zN0BFHB8nlAAOF4Bk1miK4qG99qCf0UuQ7UiHFdJ+jUsNTz3/1fQjp32t65csC7
d2ZLor6xLQK3SD2SPFo2wL+OKZcQKd3zShfmDCoARsDIfBaby9xYiJvEg5AcLzfFCSHsdpwTsme2
W5WYVOh8JK9DGytnhVtBwcDaG5M0jXAHfKyWueQLcmeHHWW1UoMaBa3kw3DzY1d4A9J+M1vWd3aL
9qNUaDFJ/6yZyEX4gCjOIBVx1/K717601YFZZHW56AWEJDiSx7bA08lCZhqt0Z+tj5156JEJ6rCz
53yG8cCCahdMI77CPkQxaFj5BCz0Mkv9dRF3tIy+o25k0zssLmNZXnj0Sa7ZcySUaj9nUsuEkx5u
sQu+71GJ6aSBvX9DMF7a/X3zRuigIYzaGidDkO0LOHpQjMB6unA/PfflL8QDFAo6hA96Ji0HFBD1
WbPtHSGLgj8LvA15u0To/LgE4M+pvCIq9+IVd6pL4b1FgJJprpPYw51vcuxkkHGRhdrVGE7cK/zu
PNbxqeRUEv/xeciqqu0s3cb+R7XS1BQJGxw3ci/xDMt0M+QzOstT7AXB2N1d78GlQfAUjysOibQ9
e6u7MEddjrlFboqgbhkb41zBQkErwIyMwyzw56omKvBKh+qpUC+mbnQMEh8siKeWK95ApEoOu9Vk
cta0iglOUHD+4I2VxJxWSoBfCOWpjl7PHtJDGnxLUhopvsKHy6ZCHMXRw5mdRi81aBdM4PY2eZuy
EHxn543I6vZ0NcU83tJdJTeMRN3gWF8S8M+p6TcuLlfqlypmV1YDmc3tLe1oPI9KYpxFzo2j/Vmy
/NwNcSAwb80s/gjpiFI38SdL+kiCcfdz+yEBp26nLOHCBIOZqDGoP1QpVOh+82vFwmI+NL3WnLhL
v6mZSOA84A+IYIJvXrnjlCADQhUOFwOzOK8hJfto704ucwdLWYC3hvXQB7j3PX5IncLDrkx4EPUg
wiCkrLY0Enehc5fcj9bsjSAPUwJeOTbRNbuLD7CRYGLxf1Gb1VbemqzSemEbKKP8Wh0akEdmXFBE
zlw0smEqWiE8PKtIFFVvzRe0zjQ0IKMaQsfnh4Wfo21KyqVWGOynmWc9o1YcR9UUe/en/c9LfIVm
YFGcdOFBak6bBBOmxxPLObnZO2/wLFR3KU9ZG3b6ZAknqLKKJb21Ne8V+Cnd1iE/caRs1dvsW8bo
2ijSdtt5paNA6gc4yXuUfc7gW+IkbZEgc0guPgfwmodxKgGJVeY+mu8OKvaHsGEU7PLqLzIeG1HC
rnBfGHB0ORcpOb4dYxIhIQV/Udbte8o0xPev/1T7PBAqNd6GsSYtQEuohJ+6CUxDGe6p881+ofHX
ijTVv5M85nct/FyoT6wLMjCtYfL0dUesF0ahpj+vTAG0VDAOjQLwKGSdpfzeYfKuSEs7pdWOTLE7
NdrHEZnb+9Di4KdbqHmOcv2pWNK03U/HXsDgxy0DAlgCYQ2SapixmvCoM7vVd66nKBJDVbBxpbDs
8NdLoJXm4/dKBbIO5gZOsjvIyx58AHslKg+dfZQxhUayUfgFEEjwaD09hnCEySVUKIAYsGM3+igk
jrQYN68rUF9b5j1NeHklV38kD2SE2tnq100DsJHKmADejxcZtR8pa8+18J8FKmZHLTSNe3CE6Vb/
OvG8DmsauRghgpkr9WK3wKTHayMT+aBOuNKG84Tr9nL5wzwldkRXzXucYe/12HIvhextRBGyBC/O
ppwB5vNuGnJ4kEt9UOpOtkFGP70z8RGWIfHXVZ5AAQb7DPjRbMsX4jRI0/3LPVjrGmN4UQjP0rZz
npawbZJlzy24Pe857KJ3tIZqwhwSrMaAuspaJeOgzzlZawSY5BQPgJ7Dj7tcNwudcb9frY6xgvZY
qJBdl/EDjKlGp18pYtif/l1jDEGWNPyEKXnXStshrLsKzYtN4mTbs891Pa5vTr9PH5q5xl3oKbXp
PMErsa2LHxbuS2soei1QP++J9syv5PtiO3gIL1ogWQLeDsWT14xk/daW16R0mZb9Mk8tWbVaL++8
iXF/6VqYEzNckWO4PhZhYGYtEsRP+BAl0a9oSDcCMULe5GMG4oMZYl9wRM5RDf4PTyZZwTepZXsm
blJGwx0XR1aK0He5ontmXJYUrVqI57zVTd7N9vlEJfe5kGlwb7zvrIWpugIQ6jD/vTKzR/CjhXmr
alKDBhiFZovD0ddUqzOcqcoCxIFJ2+I31weNZ5CJPwLtx2NnIJnvFjgphKO1Mos2CrT5Su29N1ub
foWzkrlhsfvUm7UBdZYVI4lh2uxIqIrZ90y86NHyhVs89xIX0blz/6Md2U0N5GVWhUSvil3o2A3z
DlUKKRDX46WtXUa5MZKpvol15q5BvpCHFEQrmzx/NWsO3K+WcZXLu30eAhLEVcLGM07iOjXTipcL
J/jtIeKScmggVUdGZKUqz1Rxvjs/843wlo6QG10iTL5VxQoQIZEkwV5IjXeYKd22q/dGEZaAxkNH
GzvvJ1R0IPAMajT92AzIYO+VeU45BUUvYsOFYeaUmjZdTUDXvZOsnNYFSAVF2wqiTb+z2wEnjUVF
FjKiHVd0ko1Y1lJQLAMs2zRhpNLuWtaX2cRyk4anz3CcePVNYR5443mwqgohaDKwg1MTZ+4LvVpf
dS9fcBLDXaAz/pSXZwYjriYnOCEegEJgq2qIhIoSZW+cysZZgm8OYGPYNKT2OWEaad1Fr1OBRetZ
PmBKhUr4bruAFbzHt4dfIZ7tIIueHdynzGIK+XqIkW7mc+kwUB0fd/0+VDwHBLSSEgLSymR3ur7v
ZoKHs9lkaJmrnR53S26u0EOLDQKBk+Yyr7Qg1ZqsRFt7AaluBIl4qNVOpeTx1HWNFO7cZdz9WFnv
gtgROOlGcSAeN3gJ+X/JI83o2XwpiEW810mnOdYvltjyQ7aK0bBoudy61ztZziMVZSP9eB60xWUW
PnmtKbSVKt1RQoKGtC9jblJmtO3ky2JqGL3hMIpl19vHDfMNRd6T4q5cq1cOTpzNntp0QKiGw82t
a/0wNuajpAd/LkIXlOc8fOU0GD6Z3AMP8myZBcIj3jD5+zDZ6eikYReIBKGyss6X5VPYziuF0PO/
8jTYusrMcadn5DraTYfss/UrWc6vUOzhSegScRvFZgXYaR05NIHPbIUy/SpZQ/jvSHOxa5ZfPlpg
N0N0dsuyGoCdbXG3ELWy/mnByKcV1oSCh0Zj8tFmP5zaAi94o8wcQAFegrrmzKkU5CG/B7DbrWis
Ep8J9rn9TMgrAh/u30pcbNpFBHJFHvFVgdoOlZxwKo7kY+qasbWVmlhMYkvKkuQnv7TBHWtg1623
Yy/T0JSaKFU7a66K+rqm5S7M4kLmUF31tVXzvIoCJqWsmDgrePaDHdiWIC+VucY82M4aOUd5gq7q
D3vmLtvyotVX58o/AK8MMFj0MG2WeqdzRGYmTK5tzscI+hz5NHA0RXcIY0cHZ22nM9cPkeQ4jfop
yW5YckyqT+ZfZKXVKm1NCSunv48L81JMgPTbRb2YC0wIdSubdK9jx1LDUM7U9PpJvQLrTh0dz/4S
MnAKYeIT5RUxSB9WJbUVwYnH1NFfTh5oyxC/RotauM0t/2OctAFfmKKthhJ+PiWHPSoS2GU6IeiA
OLmuhX3zXDINMhV7S4zwC08XWdfHXyNWMLUuRBCQIxR9XYZA7ThKTj7WxQj0yRcrFtmwlA0Edm4Q
Ch9oRL/j8uZ0pQoCDhpEPGDqicsR1cf0Vv8cYTPziOmY9PRIZWxCmvbaqidnaYuAxyenS7y/cKZD
kYJDkSf+k1gkvzJjgdYAPC/G1rxyB9r2LcxTTqDCF5nJB6QyoTj4IhUVA7dXfQNkO4mhu15OeiiR
DQyPSs0scjl5enyBtkphJofNsL8TmuNbl39EzN1WejC89sDBGeU6i3uSrwMRVaza1b8MaUSTPv0S
D4A3j1UhW6Vp3xnczZjObhC2Bel/G1DlJT1zhBLSnGwPEtb0+bi0NIUSOVmjtrPOwozznqdBNxw7
txys42NDOPVJF5bMTfHnnARrphLTesxtyS2MHCJG8Cb8pJ/of5vaUv5IsoaG9mdYTZJj1MlCp9JH
Hi6wrRkdTSF7WEpOKUry/Q8FaAyFd/u/L1wLmt7S3Nh2jqkez7mHLgK0uulppFsa5hRBanAgDoAm
qOfEkvPq3twKkPYRRxPh5d5FKgy8yz9TjQ6xFFQk8Tv5CcD9vYEzv3lD9LRcbNnPSumcAI+YvmH9
gmkTlI/gGUNibululsISD7x9utZXAH8pcNs8ZDWTt9DV6Gte4VvmsiHVYWWNmgrVqMNXLDMaB+AA
UipB+gbyzj68NbeMNOakF/n5G0H/vrCFfRF8cr1x21mNg8l6gTM78NK7+fXb/76oWy16MmsCBW/B
IWEIb0+f0Z0uEuQGUczBBpDNTnumCEyIUKxkp3PZsIAm1mlu7GbBaO43DV9hYLnxf1ItiUp93gLE
fYHaY9rEIhC4Mx3AXiX4jV8CaTP/G5I+ZPKuwwubvKKfX+yNSsJJmSprYK/y4XBh5hmuIGI110kK
ieq5BEl2TSZbQP0u0VAGNgLOhf5lA8HZoOO1GFNQCHk8bM1ej9HOP9yaEynPwxOgq91Vc55LZD3l
V66uy8AOb9Adx3/51HJ2HwLHhjZdb1vPodJ5UTxNVfE2oKM2FD13Ez91wooNDhxAurGszCAl4AHg
BrJa4F77uOU1tQ3IYpoWr0hm38nJzjNXmVR17S8v8LBV8Llf0OusOxUReydsphIKn8fxbFuzqu+A
JsGTGT2PkSPpSR9wul+SC35Et9ChtI2v/P6xb0OEGr7i4eU+QO5oQiTZUsf+FTIBMulUp/4skLVU
ushdu1tJdGnNUArE/M2qUkLWdNTbnqH9Masbk8YaslUTO4aEvllmrWoCgPtDqE8wIzWXoga+53co
RloN2B6TKS9ubbFT2U1QF9qnu4X5aKG5KPVK0O7WWNY+gQMZ279a0B1+muUlqg9pd2wArJtyRzTR
3PO8UtKfCoDx9uuqCxvaWvdh2OsPsNkDsUgvW/9a7gnt3RuvsusovpmhZoOmjIOdGCHK25LRV9tZ
kaEDKBLWMj+2Z3ZFowcWrzjGp7EDEV2erxMYWPRGS3jODbAhNoIu9u1ecuHM0/6cbhBv+tQdd8u5
zuhl1+IlAG4+/H7uTwIUN9gYgalkBYMXbrywrqJjGIuI1Knub+kqmm/+sLqkQ5h64V0iGtslpgzd
Gl6swVD5Mabvtlw5Tzwc50B6dUQ8qa+BYNegJqdsX1NCdMVfjNebav4m8udp+JgVD1KTzahkouvm
0BgSxmnnhdIxxbu4o9GHCa4wne0bVy99gixaIaKnEbLhiVis2Bt3fbZ8DI9qIl0IPBQ2AZA+IFob
i+AXl4Jl5EkuG14NjaEVM6/UpuCU2UI/mKxhjhuPnI9HNsKRP7yM6ISJRauTpjek1MHAijRZFdYz
N/OEjQIoAu3g8hpyFt+u+8Gx88fzYHwutxoS827HlbNGuIWTOPZvMJcuRCKJSRTXD0D8gE6OuTI/
2ngB2xHk5UFyyyKl/KwiaW4KuFr1ER8edslmzzAzD7dI9COLVICtQlQLHDErjObqAm9UYBabluif
wyBLcxahQw9xTFysTSedf6P7AWTHc8GZAJB04DeaEpdaWXuAF6S78xnTRy0C0mNqGFtOvFmqPXuK
aCfOZzKQJ/fHI028I71ePXhZB2Kc7GOFQaXr7iJIgPYch7tblBWUSYf8MLgU+yr4qPRzxiqY4MMW
TOcvtDlQoaqeLacaSuX7lgQj7Aky17rUt2b7aXR3uW0BzZZGEuJvZREjGStB1e4z/5D5PCPabWQI
ECAV0q/SSO7Hr7dNupdvSmLthw73NNq0WeRpRizuBAIjYwuaBUn+lh/s6a1v8xBehIOf0VM66K7+
vQpmvEc8mOtuA5eoDDIm0IXz3I6HGUXP5/HF45o2vmDTvXsgsvIH74b8rpJ8wh3Vz+LsMYBV8lHK
qfyx7vAt+NZOx7k/cNBl+4h+6OttComAPAu7dzGrR/YgsaMU9xllmv7MWO3kn19maLUSTMJclBd2
cYQHsD5bOmZTJaIcQmqdraqr+ccJYWQserf8vR1Wdc33qf3W+lmwQUk7UjI95R1agTw9vb7UMaDy
npXMqAFNWyH7iuNFjAEJ4CSnKwQ6GT/MCiMHs2q7VgIU9qohzRb5iUpEAkwlNrDprQgfNWLVdhl6
2jR1HUDriN4BbYuyeZo4loLp5enKp5BpJojsXB1xtNCngwTq6egUV+vElYJROz0eZXgjZ1dS76SF
QPRk9WIutc9bfLrV1ymCM366LUzv7+EvNL3fR21nB2eHxqHJDbbMEoG9AGzVP+yo5By0zY2a19sQ
vk58mrVw2lGQKSahM8tNCYiMUgO48r8omjQ/Z0pSTArvqjSO0+kY4G4ZJkmE+SZhBYj8EcnwjFjD
JwxMBzCrY0YX/xVWNiEOhUrlhgnTUgT1zJziRAVBiQC33wdmg0XlLbg61UlnEaUCJU7EDITeg7di
xFnurIaq56U2K3LjKw/u63AP09qUs7Ik+0xQdxa0jQj7HSbX3lL/Y8ogVYXY7QqbF0cIi/Kpegpb
7m8+Pbj7Q8h0G8OFecHmpFlCuSJhoFkNfgyrRbUmB/HGDnkBj31+FY+nb8Ep7ORDHlfGZoT5/Oof
ZjIGjiSrV/7G7csHhJdkf+p5CHN0wwpy8BCsPjTj+5TybbhUaVpTkhl4kuRVpEFKsBEw+ZzXux6v
W22PzSZFe7f4WbDYupqDpJ5aABa6qvwy7BO4vWQdA8GUqkZew0oU0Wp6b17J+3LW65RL3r4Oq+lN
AKiKoV85I9nIz3UWqDv3vJY5upkXqHPLxUk6QZwT6h4WmATAWYpKPgjTTnzNLZ/laJHOZ7HpFck3
TOQtEFxtt2HUI+f5hTY4OxLvY2VzA3NXStO0hxhZCnC5wP/WG1zxxWl2GPa2K3uGNKTE/Kql58rY
HcAkjuWA/EG6J5LuuXKK6Hdq2U7J0JouqpTUuTeb9A0AC1z7+WkeUBP2Qd1J6mUki2+fQFzqvt/X
ZUBEO/CaM1SG82tsT2suR6CxWiycl2gNfwyE3DslXdc6VJQ/80bNUo85SDTCIUi55Hrouff2yMFY
hR7A8L149jkSdYqIe5NXtbp/TawefK2ujcQ4vT1n+4Ba7pKU+bA5711vqEaJoCHUw3EY8OuOKd8V
yZiGtY5oQjnR25+oLzu8NIqcymETU1H/Zqzu2q+/0ymXWU3KT8eYjEHa0hvlpYzRqsUF1EkIhAeq
s5pJS0yGYumtqq3tD0I6ubWR8COWjbAi4GPujhEju8wJtV1sP9TE9ByT1hTM3Ct1Y0yAyG8L+dTy
3T0pOP6u03osfJ0RHunAvUD5M7TJCOYP8WpxIlUP0PevOmqptMyrMie89WfFP/pdhfTIoY6EQXv2
Uene4WUauVkr3HcjNQrWwHflygkmQCYDI4+ubpxVkdpPS6XpmwFiIhzgL2MPESDQ0cBulvB5dOrh
oAidqhWxNQ7RGYjEj2m4RUDDHOzkumbLpmr+ep+MRVgGrqUyUlqXyPvu+CG6Cl91d3rXviJ9n/Et
HUAQfNNW5jl77Y6mg7xHaP9welhQWcr1Z9MLWaDqiWuWinRx7mcLIi29Zz30BdlZC7kQ04wGVtnv
Vzut5nN42nCPte6BCKLeundkwtW7SMeG9G4X6AQpjW9vEryO+eGEiX8EBPRybtXIcYsRBMgJMupe
oz2SJNxr2rv3BIIWY+U1vJEF4EkTobl2REuD+qV0jSt5hRPGhugipfMn5CvONjLfG6DgXw16Xn1g
R3sdWfQV9SfoiwHTCEAs/baGqT/6DrcrqoQZVplHzK3OX01Ugvdqv/9MY/nvvd2OhoJOlxtxIpvg
aWrEFQGGPWIoLud3Ci6Zk1CsEqodGDfjHY7tAM4UP9NPAHQifGnk1UDidKmrkifh9MHNkD9Fc/kz
wTw7JJ+DHjqOMX5lCDWivmw95CuQj4rRHKXNzH01Uxcf4zmXO+bjF62WHA4NTNUVBaf55VclyWgL
NrqWK4nBBYKYmDNEgNFoqJrMHw0lB43u2jGRIOeULFezgyU1ajVYC5h009yXXrKloSh8o9tRhKjT
rx94F7KMG52GZD7qxXWLaVZxf9uJTWBX7g2m/TP6OYLFCovFQTijW/0JHL2yT465q+vkmlG3deTJ
qlvCPA+wn3z0urZyRm+gaJ+PsqsMI22pBA4RYghlsKa/74f3Kofsqud7IukH4HgyelPahlPgMmOD
w+iNntZ/mELdFvqhaFHwLZYmQUzV1tWDD6KWXdTcRyxx5wkijt4nnzKWDoLwDLa1BsB5Ir4NqtCZ
s9uJFYwR4SVBJROV4GWmgfufPas42sTle3l2dtrDZy9kpFoNJPQ81a5RWslSt2J2d+K3NBBKTMLc
SNDHwBRTiC9tr5CHKf2nUz3LubDG8Q2DV0ygEbMwn34bO2Gu/n9Ur0HiDMZKyJi3XfsVVHXVBS2E
PlSVlboCXBhioJh2UG+dccZil9uj+Dw1XAJHCypXc/gfekmBMf0YmOreZbZMqb0BmF9nYMcLjKOb
G1T6xqGoVkoq541DIR3BOsR32/3MsZnxu+XrpDw4j9d5D6BRiX0jPiauyKRWDVHZHeVGKpkdLKkK
mxj6N4G006KwuYn/iBprhZqgSCVFNUJ2XOsCislY8yZdis8pzzKE6wGOlPRc75SMT/OFCtxwWITm
L3Uh5upbtS4O+M/y+r/k0ySNQdQ7SGdW/DI57tHsV/6lFCb4TPPQd7PKEVMmHemdkAOnbyy5jzEU
wDHgOk3XFSAeew+7lYaZf828Rln1a4Jvoax3uUozEjZaLm30utUoGWJV/t4T7e9JzDf6MtZuJIUw
x3f1JZ7P/oU+8AeWN/9AiD0757sd1BdM//Wv66VlBYGBO3bEUPHuvcwEtTjlvgJcFUK6uWl7t0qW
cw9W4IQx0gVTINunfPVMeEcb32rpXXoMPYJr7yWf5fYWrqW2ToGC5ginzzkhgDazTqLamALNc9yF
6p7xIe6tCpWc9INw6JhVUBTzxs594ekk/AzJUN1oAKLDnhuY5T6WtlEVUeljTMpUr/oEFCX3oVtu
KboDcw6L41E675S21G2cBULDMgNQZsSAyLKiprNmrahMr8iRzraMNuWFJ5EjKuW4+wTY39fjMRdl
CN5ZFKhqLM+FgrBSdcLAyx8JQfWcVIX7BcY98lgXkEa4OhY6QukMkTqNCPR+XBXewfldoC7TGEyH
QEFy6mgXQwajXbmsuqKCy20Xd6iZrWJxVEksDQrlf/6rKiR4BwiVavLQeQm/2wk8m2KdB6wVuImM
phsvgQG75Wrmpv3nJIfpyFlYoMEhSCdmsSI73+PXD7TFuR098RjhEXNPtZdzccMcjpiRnR7tH3i7
0baNAW2TqfWMjGFq5/YU7GfKLvrBs7br5k1fL5fCHW7GFRs8bPaT2+0lAvezu5EwbVlqqck/Lvae
p6XqdQ6Q6i0qyrXlF+u4JIbPE+Z+7/JmWTd2sXLy68A843oEsfb7Hr2a72gSm2vuGJhH8RMkkEQW
jLerNJ0HI9PUKPfoQX2FxOL7gppTirKdzeLGpbNLNL3DfWNjSOXAgXe+IU2dfXz54SzZ1tkYqgDd
Lb6zFGp3uOlivVmH+1oCQkAUiwsjlyVl9CgpX0Vf3pjanzSSXDN4p/aIsoYNMGxo/ltOiOAHZCUN
owthV0lFFCSyLHXSxrHR9Cu8Yfnlv72G0Kee8mwy/H6AcdwNrSJUxO5Ipzn8dAGFSuQupO/bD0QU
uFoOQ0QEhdzSjhL5+otXhIShlN5hwbMwUPeQTaXEoUfGnWmYDy94bXCukAHLd0180KJYvd6NKH/P
E6sxyf9uO28jfAixzYAsia1Y3rML0kINdFGKfeUeiGuc0wd1E3MvQWBLuYIoS5UIE9oourTHLU2B
rTnSK0gQumalZDHDLUMnf96ifYIQ/hksk72ZXOlzNMqbmcvp38JxV92YiCVgezwgY4Yuml4IrAKp
FAH4tpT40JYMvqFU4RMMntSwobzXwpjSc9jH/hbMTfTJd7q0vTf5cdugO3jhEPb3y0li1xN12Xl6
qGFE+6oRyNMvVjOppPMJDt3oBNfcdWwzsNGyB0rxDU+0ffUNVCWyHenAeZcEQzCcy0Io+NhXDTmk
qPKyjD3E+bD5dVOXqykcFjwYNUHB6iV+V+Ozk26i9wJiXKNYlcUS+vlN8zJ07jqqJhfpw09slUko
bOjs1yDxuTlsxztwZ9usQYAdckk1oSW1vZB5mxAjfrp1KTLDSwRiE9PnGZX0aPJJbFdDYzzRBAnw
MHsrsfrx6pbkPHWcYckLm+R0svSeK4kW5ergU4ZO9qWtrxYNZqkKG1LxrP/U6is1fIf4zXA8BLXK
6uCdUz3pwTKZG35EGf0ZDEIckaeBsgwfzBEmeXHg5gDj7n6Sf41KAY3EG5M2u1CqJ/AcGLeWheAY
gTyFX5C+/Bphj90hsjTRL4mjnKSflyEilZ5SpJs4k370GGzH9WWmk0hw+lvwKLxp3FD2ixy9sdu+
Ftew+x7pFSwDbG63sgZLPLEF7sPyDbWTHMFt8NAATdYIZHjvdD6zq0uS/24bZLUNtVqSleysXHed
8xxa+TqKEGNrCjeTjQbQhqX+vjmSZLxQXiDguDpdC5+PwOn/jpVlOWQxtQrzYAY8TpfQ07GdvWsZ
KMs7nB+4LxROQL0F/os5NaFp5Dw8WfbQwRUCti5mdlNdcRvY7VOjDM/8VmiW/cepBt0Fpt2M7FWO
SvNgSJD+eM94MgpaGTdSQjAgSf1F+OzVrg5U06C5rWyuYIIwJA8mig6R6wLFR/TebsQz96f6MkxW
j9YHIwo3ePgWGUvE3j+/2/YWG7ADLxIyCsQVG+zyb3Hgi3oAj5N5HIPw+OB7J0y0SWfHM/qYfQDu
XcO7clejusDWxCmyIVy7P8W9lOf6FbkIos6x2ip+FrH8pAWEkXQXT0XeF/9FoXs7Rj6TJdu6AfRL
Kz9GgGQOOXT8lB3FP7j7ymH5IZGGG6S7SsWz5fpfsQfyiuN0mvMMeAAV90U1SJNkdW9NJgaD1Rjp
1JLEllF+R2UtrAQWZf+Md5bCPcGQpz8MWruOhBw+w4ijZa279tIkGjEwBK1TEmpXTX6IbYWNJ1h4
GHcacix0r77LwewzetWge5SIBOnlXYviJ7Rrhxct3zcK5FkH4WutagV3UxGB58X1EpfxlzKTjxg0
k5zYQCaPcCxkF5q0OasjWmOEyP5uTRU4xtBnuiONvzKRqN0M3MyUk4J25EOS4Aix3gAgXa8GfC6Y
nP5jwbJsWNSrRvOVgj5VBH5KcCMD8YIb7bsUX+GhgpH/7dDaHF3asKDvW4BclVPMz4XBcq+iij2K
PoE+XVtykzqA4iMZrOQRhcv/L9fT08r5iw59VBqy/q8BxDViC6TcBeTwQ2aM2RkyNUiqay9ewHWT
R2DkGZg6jcMP4qaTON4F+jKZPjwbGurOhgT+VALgic+EMZLB2++otZGAD1xzbWerHfrB9RNdrU3R
1Aca1uqdy7KiZ8I6i8YqOWBYyucgLNwwj7GkhIjPN8R0jhp43JnZjLyp+rBFJXjTr6sDCS3GPi8u
k2NzopGsnubUiD5EVmxb2pmZlAHHqLvf1R+o9tQFHWMlrq7i0NfKbs1gYmDZ1AFNTSfmH/QsBrrV
iSqxKnkvQwu+tpLSiPIEoI7I7r3MDD8dgpQDp1iVxrivO2zE4qv5v/dZ65JspUGyFmDzEP0KandU
yyJcDNFf6cDu5b027BlXrs/prPd1QeEM7lvi/Rdt3OWH6DCxqvXDntIONQnKYTsKPZYmKLmI/wKC
Gqot2QlOPQcQZXVVbB0N6KDDz62nWmZV1N7ztihQhbQAmCa/fJtZqlmO80wvNWEhAJB5ZEyAT5xR
KL0+kHEQcIyu55S5G3YaY3wDeHx0tM34Ol0GX2TlX4vf2LbSW79pOGoO1/7QXoZ3ubDl+9Zv0Imi
JhtJcTxzhgh165aZTw7bBhcT9ube8cFIVsIOtEM0+KUO0ysJUAGpYZxBsqVLfNX4pcJ6Ky1TMzw6
nNjR33/X3bvbsQp993VpLWappj0mn7ZX/7NgTBR/7YD/LnrKjtxm746I6sH/B+Xi6slkvkYhsLJu
5BfwqD7QXghxPWX+RD7lYzJhkR6muf/WQIQtNWJQllPrttfz6R6UgbL2zd8JoXaN8DVXnAB3NFPD
I4qBaZ5mvNnZauszswm3aVp0Nx8lEdK5tyfs6CA/8EcVqRt8zdaJ3aCZsOruC8lYfqu1w3Tz7Ogz
s017y8rmu/vcqQ13/dHNjP4ad99sgN1hMnXDe+9ai/eOD3QxTAvqx3xeGhyJXQnmFq3K1yaLfoHH
qb+vms+cBEdDbD2BLJEU2ksLYhpQIdC+3i32u0nFXIfF+/ZN52atRb2q+6RnZcCYifJ+ru0AKreY
JR7T7aokLUYT4aHGKv3yawOfTDfu4jQ9q76QFGdMAjGi4Yj1qzBdg3uheYiiENUzNo4aiSIMwpGi
bSDhUcyWndgaCZ1s82Q07voNdBwubWT7gVcBPOEwVjqraA13cRWhP6Jaq2TekM6eDQEfgxlT2fGd
3u6oV4yHtdWb4MwqGolO9xc3Rt5kVMPt+F3tiWLFOzZ2aE3cqHTrwoRk5Sey4S5ux3mygb4ixQQV
bNS0r6HVuuZnIE7ByG/yrT9uv/szIFd9zQ28PcpVDfcxEd805t4Vn3OtTBzLAY7SwBbUOTCZFu4C
K0JNT5xk5/gR5BcpYsDmaeok1SQ8cVzAhuCqOXlcDxF3iwx9eDIreArivzS2BlCla4m5sFddmD+u
n2lSnctaTOdbnkwF2XJbBw3l6wKfSCyIh0sWbE3ZSk9IlraQ3NYNTu5/Jv8bUn4S663HvCBpJix9
Dv1pp/7efW285nNe5ChOX0edoFYbC7JolgjV2lGDrU4vL3l6F1G/Sii2hrZ0La1fXyiHbNZ03D8R
+tzC8OikhsIGuTvgsiog1DYrKX2uuIwuASXRyHq2XvF2FMmxkqQu7i1jeTKtx7hUy1mnBM98peM8
Gmdz+XJ1Deb/P/v5/V21efQ0CEoZUfELLTWAaA+7iv6bji3tm13GW8Hu0h29hUV56v2jVPdXFdB3
zsPyKzeBBUbA1E1Rhv0yGMuVCGME2piZyFI2mLQXFZHpuPOe60v6BPgPrBbgoyrlwjy5A0pEnqJj
BimK43U+5mnOdbwb82f6wpFljMl1ClS3Vbv67FcNFRRHXzMZthjNZh53CNc3v/v3t3GwK4+E//MV
z5BoUBLJwbeqX6wNyBbIlH0BlJcQTaQwh/nPHf21piwCbycjTjJ2TQN6X39721/E1T0Atsv/MxhB
XHFKizCgnsZXukzFOlgHdAQt3rVfGrzK+zlM/IStElyEF4USn2r2ThV2znGvuPT3wmbSVSgVDhJZ
SMvDCXsuOXsavVV33SVSfw7otKViCo+Yd+vjqUxhTYoglTCc0nmSjglEPMH9h7WlEkWu6lSiN6Oq
XWkosSAs/yKJVjZF0YXfW7ywM+YhXLI2FFurjXX+0j6pJ9SdjAF7ziKeAhwiO1hEpMph0IQPykPn
VaJVq54I/nwjCzhlQ9IF9DMUW3G1mgxWROL/pmiAKQyUdcU6Ql6xtk2JpKg0ZKCy+PwCCEQZ98mZ
zQmYfqfZHJ7khGnziR211p0toxo1TNRb8/CxTTzmkBVDamFVd9oeL2CBEjylrp2hfafmEvLwNeYw
MVZ2WctwoE3RSfc8d3zQU4Ib2WoAFsHgyyYbNnGttNQ1X2PABjSCCBY4czMWl5jqC/xaObI+79Cj
dN5WoL0pgeCjQHCVzZC85CTSjzFZ78Jx6SIvzzKNOmRqh4tpwJyF5E6jHxLUg2GeKCz6R/6h+Unh
aRAUl5/fH3mpuLUKUhz46KaripXwXRksESrnkCVIkfy8bS+GCXcrk437ERgcM3HqY0/6LJ2Q51q4
w4MHPs+vY67xEGoIarIgrND2QGkAirB/ou46STDSFNF3dSzpl7J9zPyMpAimJZyrg2WaBAJr86N6
QcCTqNv/jG7MqBmkpnU1KfI9uky9tfRII4tSmQNW8DT3TytCWODct70ycTwqlHoB2yPBaqPcBP+l
n7Il0N1mhsWU/yX5fRXS+t29jusji2Lvnvh84aKC2+Zsf8AsdnzyXvaY71/W/+4/q6IeCw7a4fqP
5BOkuVZuMr0VND22F9MUH1GhIZVN3JZZ2oBK1Okj0Wv4ExRYU0pr3XJA7rShNosXKBwand/nPEWq
tkhPtrVjWfgboqofgaJ1Y4+DL+ScgqMMI08hlAqE6soEdYtemxx2St/WAGRyUiE91mpCFs9TGsIU
y1VtwrZjlinLNBvxjlrwiHNAingPdKHvSeNinG4779OcWyT5IuK+6vGbzv9sEjx4e/yyz2qikPeK
g8mUxj8ERTBRt8sfbC6nWhKkG6n+mqaoeubeFvqrsybRorJXPC1/Gcv6tjqKRLsW7d8JyPPZ+jaf
hTYdWlYlV6wxBp28LhW/zP3Pf+Iszd/S49su8jC+3vWZINo6m0uzzYHlZvPgCpmWgghHDwaGwxp6
KaYPVmcTAuBwqovUrRagWDJ276jwPvkcRsFvUA7Ki23bDa2DeoOnMCWPbOJeUCGFSsv5mSL1Ugjx
CJhNZLH+XlhrLpGnMf5tYjHIxli0AMh1A2xjytBf3jLKUyzFISH7vEjniXjL8HTkXokIRp8PWWlo
CMSd8yvHUQriTWbUnqFe+Jxj5UzJS+I7GfaB/T62w7egx88JpYureMuODl+0rQ0ZrI5qZ8NKykIE
vKcS/mEZWbKBov2o1tt5hM3vy1AGHcdyVcuRh82UExF/DtYYeJrHdTCF+kxc9pQHzkZa/WuhWuJs
8hIQc42cs2i+kcGxP30TT/7sSi+t6kQTJRegOGKDl2JR6AJdqoFtT0zJPX61B60tsslOy5B56gu7
KJHLk0+es1j9kSC7uE75vs6mhDAmFlVb/v4f2rbzRILKkYEjFCsM+4Bywh2eD/3zi6Jq1eAC1vv8
JwsWab5SaUDt72SVofRPhywkwYeYMinvZc7dpkUT8gtoN/NCMLhPRwgDwocFWQ3yIbR5xQjuHoe2
czxsCE+N43BRzYqnDaI/5MpnUwMWJjATAHVCDa7mN3wi8VEdw5iG/yXKz1aVNtEiurjEZ1Y25dl9
blDmy45GP7RluxyKXUNBzYBoSeIeteFN7IoNgEBuUO6tr/MAHq2zMl8ueyIvmDwP3j/GsTydE+pQ
3FDg4+HXDAuUVMihdLHiwp7xK0Stecc84L6f6gpKJKVHHs8A7CNDTOm/slz3OiE4d+MrIr7zVMhp
+VvqNbwiwrk9mo+sQbU7BdTUjLPVDmKnWQVbYepMiRXsjUrv2jY5DT03+LTrmTFAfhm1z1REYflz
aae2Yy8MFrQp6Ust/5aQk5NLsjChJ3qSklQ63FEXJl/e/ZA7lykyq9/v105YW2bFrrqp70HolbC9
PF9bb5imJWEtjz1aXQzsbAix1g4jhdnzgr9zi1utL5CI51fNx3XNE2UooWz8Whw+07PH2t2Z87Iz
btIlvmqFnw5k1iWpt2YwjSrL8t71F8fWw3GDUgrXAAH24QcOabKbvTNJA2/n4W6NRXXox1Tz3xEl
enKxvCwdXBAKooDykNW9mlO8MqHrC+TBVDAiW6SfPwp2FsqnQnbvY7e2/DOgYrlet0IcPIIfFhuW
X4XNIgXHqw9EY1fgTvSfsiLb9GjXq91Uy+EG9R+Dm0sEj4PXouxYJo5992TskiyhfGrrj/u2pjKp
5I9KnboFK0+QjHyd92fY0bEUw59lhh3K6wvjZKQ7eDw/WrFts9BlbXkFutsG0Z7k3Viv56wFbB3r
VveKy58HbWsWGM2MAQII6owbfa+xUXRuYkO9q1kkIqu3r2uEjvN6UJpL2iv5SZynX4TJ/17+JjTT
OMN7K0QNrEGDF2Za6L2FuVZufcodPrRlCpDmoDs8sTC6/y+GtF4kupANU4RHqUW/Ky+FVymYMAwr
rp6N2MdX7O6V0vnrtu1da/36tYi1OBbdJ0cBAb1Pe3zeQiO5VJjGLf68PXI8Kg04fxKQOVHQOleg
nR8X4FZOy4h0SkVf1jiE5jv2mHMTWazUHFlpGGiZBGklj2bFbpTX6zKKow0l/1nqliiCYx6mz3jt
MLO2DnrCk+u1zSlWTK9Cw2kS5STvXJ3v7E4yWCKrnN80SZNtejrSJTRs3t8LnnMEFbInlK3BYFRd
5vIWCLQt2KaGMuttyh7nNSOnUdxL4oppSopF1iO0opjhs8DFJrnv8RMUD7ZX52zbWlh++7kuxFe6
S65ZGi6tEC8WN5f9ydO+y0C3kj8JX5kMrU4BVb7lZCcA5fLq09/T8TiR025MeOP2erTIkmylLRAd
35LoUaCtF7/+FnNi6912CNxTetkockJYI6lFdJuQoBKviRAzjkXEqRl1I9QIP+q/jn39KpVlHLi3
ka7TNPTSbdAXrsnyXM6pi2I02omTjwTicj2wAWtY+245Vxv8dkrpKx8+kta2UmLYmqgXxD5Z9TAc
cgoYwHXffyUQcpo70hl2eQWvVwSnRnadrSKuoj0/8sSdjSzFSPvei5tNztLFRx7bjSElvKJHKhRJ
eQhOKAOItR04VfEZWzCi8s50p8A5La3UBE2DzLGAbYG8GpJQ5tAMgUjE1QuwYbXb1f+K3B3OxFKj
E8E2YwgQiOfzGiJcR4jsDcuQwtDYmDp9B3VvHId6trS2MF1lF1XUG36T6j5wGransFcy+L4WpfBF
TtFUhegLgwd9ston85Kmqm7iOQcpITCG0ewI8cjMnRyGM2ccPr6Z2gjfAuebfvWt20nEwJ94fems
Gb/ta9p2m0cYr903AZdRZH9YADhkcXa/tl9KtSamibc1/XoyxBRyGIbdt/ICUEp4SV1zzTMQyuMQ
StcE4P0zwamulVZmI88eBj6QhKryp1SOBE5iinU6lYsT09LqVHcZ2g6h55/K/WoZjk41oxmDCKvh
rwl69EJ1oLggJl4SZ53b1+UBNn+4hemxeg60VEdoAVlsPm+tZcFS6LLSgdrYZLSGEyTbXqM23A97
tAUEKaBkUPUCdUFs/kkBaAwJvanpNblyv8AzEqfuBae6VkDbvwb7FZ0lVVoaQ1LxRzw9csgEELnI
/O2uhY+9wi62DdCSWONggzGKjkDIf+zQKJGz04EwFPSN3vyh/ombEDXTUqPi0fRMLmNK759ptM/z
VXhimU7i9gyoVFPm4VoQsk1HQthkacu8flGWgyjS+lB0BuzfAgL6x8DuDbf4xv6XNwoJF+XkluMr
+mAjBvz4IBCPnl86crJFc64hb6V6pJAneTqOIvcVHG/ToYKZ0RVNI98KrV677F+faFV7Nw438mIf
oiiOEFonPlG7D2N/K2/WEHIS10mb43H22DEzGUyHUqe3pAIMTevvMJeVF6dX1h0DYN59VI9OQT+G
PFLpN6qp8ZWwQCM16Son0QZAxmYa0OOjMwictt8gx43mVM8rkjVsPC1MXc03bvX312hjIVAuJtg0
Sy9wYjLUvatPRfHXazXvcv8lDV5oBpcnypIkaLNvpG4lnANRZHF6eQ1a3Nfg/Fva5o+I5ifOReiG
s27SfEpm/3H8YWfgchVuoAo0ut2a/H8paYh/xh5px2qcPPke2qUDMR4sTVjV7DR+X2HYLaWZBZFN
N7SS5qKuoILbv1rKAsRffFM+NTEqkEmdVn8iQYBH/dHUfpWWyQDgPkhEQnr+FhsUAP8MWeHwO0RQ
XxAKteAuiZI3R7/t8M9vRoMNj5WosQWYUwlY0AvjztlYmJ+h6x0GymV9u6I2PK9JuqhdEgzbuL8C
RpK9JtXS12YUAGqhOiRuFoAuRcIhVBPw+3uowtoX8ZXgQt77mEwwTzOMeXB/b126IDFG1fZPY9BX
RxJi2tKPP171k3DA0uI4WPF8HLC2X3Bx5mpTCIUtbEWpQ4kgSfMfrThbWAHn6MnRcJxkwPq6vzxN
Se/kq8C3vsOJ1/BBBfxvcLidZb2nlthzuK0Mv4C2EaT/6g1TUutksgJmh2Acvm5t/0U1w0yIpBAn
wijj0bxA5pMgeDjrLZfnxazTbaCuqWOe8RLPJfkpVcX+dRXCMLwiLCiJc6Pflk9n2U9d5SvNaIRa
WsTYVMUQmuOsxeAK48yeQJ3gwHbusn3sSnD4BuFjQyhSGy0YVVN3jZQ+tuH/ccRvlAMBSpci3Xin
E4bgKz2uC4yokY7Vdzb9LnUWkNv20bLYQABvanTMe4kOzzTVwXVZjgeaYfoB+TEZAulwcrMUWwji
5XB5oYLxXqvwyXl2fgNHgHDuieSJSb06e4rcRNPjVxIkC7t4u0fsvpYYaFfuaBZQYE4haajQ5tcy
cf/1TkU4G8j4rd0WltlAGbKP3VKx6zgp09CGj9VI2xLrkfI01ARYeo9Wrz4FreIL+9QzLIRt6WPA
29TxrQyaWkXXZq6SIqCyblCnhNCafH7VKVlYZGrNd36Nm3tDlVw9fYkw93MTPyzSnL3XGzyivMw4
Evg3ZiPPs1nueY7oaWaOA7hx7FK2GTBCS78iMKJw9j7Qio1c/wYwcD6c+X4Y9CejAoATC2M2V0t6
vqHcoJ1GzW2saCydbS2W3+jsvFEwVyaXO3NLI6rNSVulvNg5hGSsDDVXDB9sFy4wJ1hyWGSFJ3YD
lLP7GK9zH8MkytydnfAvWAVkqco6gzqLsdEppVaLdZJFJmvTbE+5KzrZVvBzHPfSfh9ObIBaLK2H
aBW9oG41Po0AiCDI077pml9J6royE9KBLVjV/YHNqAab9Oj5OexCwn1c67po69IyqGJs4DT2+lJC
CyJCLUojW2egE+gWy7L8+uFxEy4rlWPD4XCjNlBQUo19JLniih/t8u2yPrIaefUB81je03r1FvIn
XiTEj+7T1woBemkqwuCMWiw5f+1lOV8/Uh03xB/f8H9cMVIWupNuxewfVwDxIvOaxDR6rees7zGG
vupqpdGgm2lX9GH0okRqbLUO+bgpc6Tbr9j8oEjYXiNR7d0smse3i/VS6HJWj/YkzLXFJw1qWTsc
fM/JQimrvY17ZoNKinttgwPEFiOtboSiU9xgjhDUNXTx5l6VUhATwiJlb9i+J/1hyrdWKKfuiJLZ
GIqAzCwcecDJENzED1+cY/7a3449/1YECSxaSGcI3WMZJ3yiQRW6djzIknuTck8du/IdU26tRIW4
tHHn0eCDGsLTEKWap3UYUqcLc1mVU+AhHZvf3xJTFKCnh1ekOak6qIuLP31Ur9zkZs62UVXmgAuj
wthQlubwibIQ3Qk12UFV9aoeF8qug3rOCeqozFu+MHio46Y3fbiulF+TpVc5IujYiuHFXTBGYbBP
HnDD/8dQozYdhQtEO9iM5UafEHkmgVV1LAWsjERjfWvzKLpVsxqgu9rWzX1gvqgwNcTJMPQx0g5E
kEgwDhtrwoKwHt+clfK+l/N04GVPipRi1VVtqmSP52qphlAnMDYu+aAduh/hJPg6N4BjZZEocBXA
J9sXG4+ntJWCiSFh45GM/0d8XrrOFRs2VBhZHsuxVsDe1FGdmO8l1m9UjYLjCGiYk62KzpERH0Sb
X2FbTpboa6vKAGslILi7gi+SKwbCZ3c1a0Is7s7TBvxQ7kBZin/ntBt/Ug15jp9/CkZ+vW/9u8dA
bwW/h7PvAnQJkgzJVfxT/xr0bpBDNqWre13N5n7djaO6dOxfB4Im7yiWYUDNacRHGVTg2uX9jekj
uxzfvnbqN/yCEnAS5s28uJUUWDDcxgNKkWAq7hjLrP+feR6zn/uUxau0U981XHMbCsWQDPBqpe7c
9AmJBnDeIq/8Fyplj1aH9wi24AOqJJXvujRTnmLlMPg1sxPozYPEghSpPFrIIJZinIIfT7caOLAd
Ai8c7NtFncfygtJH+W1xvh5Mb9livNasmN03B59Crl642YR1fDKhujh+M0ExZtY561bxQKCrjwj+
4P0oohQwfhtLyaGFtP7wEoeDzpy5OE/c8oFasadyGkemy/lrha+/eTuekag/mLz05XT+Kw4oaI5e
gqBdKZ4OdzCtuiRP7pog5ZR4rVZZv4XtD9YNWuKsqdSy86jb8eLP5BSWYS01rbEGxD7gUzTcAzrn
R8U4uMU4ViT5YkWOZNf++k73aBwQOwedpvJxb/SxLO1DPOEfOzd9VwDs+0G0D9Ohy7yKptcRAqs/
dhYHpcAtY+o4CzlRFZB4rdj4kIp3aNuUf3zUGp/tm6QCPwtx8Uv83he1Xrj/J2JXNVjWv5RkklXm
2Gx+iuNxrQcztIp0O/pc0dE8yMYgxkJ81QGHtFABS9K4Yl07ykwrvdYJBJSbSxvfpf2dll5DMgsD
dg+Q5wTRBxxgp+uzQRctrmp7vcZRPtyuP0zv5b0KpzXwilo0mMzUCo1VE12/TuBmW/10BtdrxEXX
ewu30OFnPtuDSDHzm5ILUAUAynCGHvi7FCyyYYoZoYT5ZEHrTPhTsZtcZ3vMX8N1mRhu8e86o9ur
RRHPNcE9yccFzizZxprxXfy7vxmInvFFjq+fBsdtBx75GFFaXFaaRJ3TJpe6kQlf43UTL8Y3XWDz
2gqY8f9AfxLUM28WeKXbqx31e3A4MeEcpESbNkCM0KQKGOXy8ZmlxQg6QXxlBqwtxFxNoUXSv0lr
mDHlMKcGypc0LYTj+nwwLR8Of23Bt/gl9MQkhN1lQjAXYEaiMNqyrBpT/hw7RyJEsQFOwtKLWOc9
rXHaNybG4pcS2nMolnvwUyrCShtedjiJBgC+cNwb37h2vE1lRAReKuLz3BoCALvv+ksrFjwNkNJr
EslSY63Ugkv9vLIWdCWtz+u0aigkVPncZG9NzfckBuLINbn5NmDoaxJQNB92P/+Nut7uLkwfkf2P
FSmeeTfsRqCvtHKGk7ezto9bTZ5ugpIbkCWLBd2hreJDvxa9goi21dAIlFJlr2pVTONyx44iDHWc
9gG/9oYn778cGmFoRdyOd9H5fX09E2BoxeVFttMZJH69F9IRhoWPRzLMWgDlgv1ygdNjYZnKcV9Q
iRi1wc5KVEcEq9jPth9l5x3jahokfeO5JB7tEjD+or3RzocZ/0GXy03E1/meY9dhfN6mED33uuEl
DJOQMHE+UTyqk2Kzp6d+F491ClpBXlzXx9w/DznuRfsP328JYpcZyLMWFUJQLUHLNEBLiCCJKmjK
9MxFknNzVX3kjMj1DGyMif6MdCkpQsBv88RSL1zwvLyEAL6taETUmKSZEsQqGA8CSU6XVtnlAOdR
6oUDVSbl6VV0yj3ni+V7PE1Ki5uJCckkKhpCEzJ7vO8C4QmZ8cx7iuFWFttGK1nrf6T/fjSGBan7
LX1nTN5hURvxUeVOHHgeKF0Zn1QO6Ii/1eFViFGHSOv5u7BxaWD0nCVQlNLXWQno5zB+NCRj+KiL
ag7e2tNEFwlk/65838VgINywXQQbyvha/h50oyL45pwqaFGs+6OOeuU42hoRHx9yp0dwMFb00aFn
yUQaTEw8f44+B5cMRqlRgzcfyAZOI8P92lTob6baOItWowmPE8ZiNPcpk8QpEe5T7xLa1rhM65k1
qUYqq0n2mI/6GPPeUHe+ctJJmVq9tbOWjxg51ZYAyEsNpTjzDUOKHDMcZZp3swOQ7Ow7jJXymCMj
zxqKZHPNgNMtng4k2oot+uBGrqeBA+l8Ut71aEg5qo+K1k1vIGEL21JiZpFtONkWnEzC5BPvyADR
07BmZ+g8CsHu12HzaWUga5rK4ynZzmB19ZlAY/CxC+GtqMg5mSwfSnsY3aH138XBejcq8f3vj1e9
feJmxh8y2276U0BTBJCZxsODxVIyJ6aFPv5eHSqYsWiRQ2ZyPbTOnB1OHmOkt4KgoIMnaEY+vFI4
W0adGl/eszSkRIkxjeqDGKa9V6BTFx6wSx4WGfsioDwzy97g5Aw3V/nGbJ4WTPTxdpCkNvbMDNn7
vvo9GhS+wqA1S/pDgA+cHWSARy4QjU1NKptihzjBVosw4u4SLEftmsBSGe36aswdzj/z1i/YDS3D
uYC0Q3n8ilrW8k8v6/1FfNpy42lA/XNMpmIT3Uka2Ti+wpvFrAqumiFtNG0OD8QJ0ISIqxbOahUP
Toq2OBorOZvFdlHbFbldFItaUBXRlkj+rhc7X5/ygMblP57iz6SgObzRWapDVKmJav9F8Y/xovF5
myNppmY/j2x6NxOEl7TKF/gt4xLmBrdffJAITHPirLBlkTROGDGtShWlp4I4QHLvshaRuZCee/2f
BmJ7shi30tNy8k6Aoz46Lm4BTUo2hBxND1U12wxIXXcD09vllixyHLbhK7GugY7pIzypwPDbzqed
lmgaFDP7JvnjyGbFIl/0sFIj3RLPYPeKdXZwkk/hacN/+TsYj5y8LO6j5RRDAGBySMDox/NsuhPB
qIQqPlqQY4rJjZ7KTq4bn0+Tfdn4/0+JRMXFxn12bxP+AmMjKFxX/wKLpd/cP+zDUTx0RrO06cb1
Y1rMjNTFse9WNr7tsv4yRULuVRGTsondT8puGbdW0BX5CipTTpiAXFfE3CU16IWNdHKGnF9YprOk
G2qgRa5THDT5Y8kHku9+4/eOpH4q/IiYtKOSci+FbH4BhyzJKZrBBspB1FCPwcmoVsjm4Yg1KsHp
f1C9JNXzBpQAvUjtYgp0eE6b6L/hXg1SzUZ3e3yRxDxpym8W5vhGkykPuxU3PIW1AfLrgo133+PR
knsqee8lQjKweGHmxZB47KqEWPtqczQXz2FssnpXoFkP+9r3JrHUzCsEtoQozV6HlrEUZyHvRtPg
Q0O5bMdkqnqB3osbSztguJSmawJooqmcKqLoiTBRf4G1opgO2QPNPR0OmDTbYeiII7BoJV/xK+5o
N8kVX6CNVFdvch5PagT37liWzzB2/4qaINFwxe9E7wkuSsbhwbnGnwinkdtQ+Mr3nowqnFsfXLbT
OpLMLPM2HFoow6nKcLbGRCSyfjaCYqf7bGyoG2cNTE7JnhnyeH1xKPV8Re+GCCMrTH4mSxR/L6lR
QGxjkgVzIRyjRzCYHlP13pBPz3fDeNqC5AnKC57ZClIOA5d1AnD0WV4EZLns4EXKCfsG/bSseamm
4X9ePwsUiSYJc+EYb9OQGe+px1RJhTiCtMKICA3tkoW8XcYYanEObSGqWdVywB+9ZdxWO7oB1oM5
8Xd3x+jlOxnW+JRMDbXB6fb5FOnbC+GOZzigbpn/YesChvoNx/tObIpjY5RE+mYdsHPmOlR6tXsX
7rRng/+BG/LxbIaJjoFOriFBeZOpErseWcShnR2o6pmKKjh21Cf3OW7HeYB3Pg1/zLMBC29NsPAG
7IxI+3DyNJF9FJUTXAGl0GyXfkPbkHsxsRKGlCN3YK4uqpCPwP1tRhNRJcH9Kjy5Iqyq/W91NFZ7
eX42jG2FZHuPdIrhQwaxp8doW45r5uXz+VtW14XtOSSJIfPM0g2pWEZLdx+4hynIaWlIytSIRCdW
QsRNSJUJ7npDoGC6gosTyo4Be6auJj4HgmlG64hauonCjP4v65oiQ62Bo4IxEm6SFb7WInr2H3Lc
zRubftnn4dLNrtSfVcrQ3lSL7ZCyJdSLEV4gENMeDN9+4z/WLc45FgGv0HizsUv4dT15STZ2APEu
tsBzD0mK3PBAISjGE27e9sZ0z3HeTMSVbIRtuqvzXfo9hRF2pHYkoV6hpiyVN8dKz8v1x3HKs4co
TdQVDHk7eL+eKsKl3DA9oVxHmhye64I//GOEqcUNpIjRENTMJk0IDghgR5qsqO0fCZb27TG7JgC3
8NzG+3UtIQR/8OV/YiZbLlStJBHrUl+OS8JLxxWeYGU/TtR6amxqmPUkBz0S2ttX3Ru0o7L+Lt/N
tgeWoQA9HV5JXaf4aOJ7J4QIE46aAGiNRcRTkqldCKyIIEAy2uNtmD9jH0MGieI76LYQnyRrqr2w
1lKQINlOIpk82uNwskyuBSxhI2Ni2DkD3hxj8j9MYDy9apqUBCtkBGsRijAM0xBYlFVbM32rcm3t
C3bwyAIeApyHCQg4JD07JYdyewcLYjZLOv/5BWIj7fJC70rDm/YvYX3puZwInFKMJuyelKOwxE3N
Y54KiLcceMI865OdNe4VoH+F7Y/ZNn+DS1UAspGo20PTwD718/48rZFX8xf/c/6/X4+Pb4DhAxdw
9yUbiY02XjeLsBbbEaFyAWMJORZcQ5dqzANdyAH6reqWWn5ViaoMQM1z9cDg3/I8pLhOVIOHt5MP
TxP4reySUqsXLjlw1maE8p2gQ5rhHEpq3NZh+HDjfIgnHQQ7wIfKN7by0NnlNFcLe9rLnJr+phAE
G94LyILFer+akLXecGkUbE658cPkU/q4BH32u5JjfvtF+MzpuadLYW3XkbmqLcfdJt9kqzQtDsnv
JUsYacSTprY8Ap4xs6tJf2GIgnNphpWG0Mi0aahWoUsXzQ9esHEB1ZCQs5/rLDSewF7ptGTwKeR8
YYkYh1nG8WSp1aIWASQdVpPVC1pjLA7cbjxKBLBW5OuU6Sx4cYkMm2do7yq2rhQODzWxbR3IEegS
mtwAN+f/Dw70Kt5jSTeE+2yFdAFPxBt3fVdU1g81/iNWXdx8woR6XCrTN+LxZQ/+chOu1IxouYHd
IrXmP1SQBKihjqu1lO93u1EMdLQRaEiyNuhkPKaMPu92L0R/MOm+iblrH67JbEE0fRtp9ZKsRVew
5UGiAXbLbZDvwHvytSvvPz1aK2XbdrpUWctsqIyzrzChg8U5jkGwpx5iBXWgiegYQC2CLsImEU5E
rsj5L7zIeGdGqq7Bwc0UDKpTIXSvx8S3sxMx4oIGXWmrIzoR6h2NBr3zn4WFhkQdpLxtcJbgw1AK
jOqxS9i4Aj8u0wOr4t+PuR8W8guZByk73FCXnwJbFtR8Kw4cicSegFLXrsDxNjKYYp7WmXe5da6Y
S58O7ktAya29TpBGqOUNfMPIsLEIN3kj8CpfWFgJvNdHZtqTFqb5ldH0so//zRttmmXgzVXu4v8J
zqb73pnAZr24iERTRhYFjUEwtsL4FDoOOqJ46CKfcQ2TXqir455XyerXm0JhptNRXq9SUB9O8U3j
DqZLHV3rM1yYIs1YHWz7GKaEgqdRWhayGBX4f9WfRKcON4WENsqoj2TuU5hi+YZ+qplOwB+TJxLU
hoPzFZVjSiIgajpMfCUQoVXAys2byZVL06TdgyLaSWDLF2iH2OugjhP7Wqx47S9oRhdeg1eSZ89i
QAzaElnh0lcnmpiUyC0D68agpeHJ4NFuVacyYkQU8But6/VIlIKcediGeqVcynAoel9GCjdj4r3Y
WEhL0Vo207CM/f/XXm0adWy2iRKRxi8GEOYrleiKzZsmmyusR1kDv3hzKv2KrfXhYdhhdpG9gIZb
U4LwGFMsYZIKtGs6nIfBVFDsXVmEwejAqPT3Ja3Omzb+yCQuY7LtI2L9Yd7JXvhF+labxQJURToL
ABG8M4ZrpRmcGNxrz9n5b4TxF5zKx2ZzWt6Gik6isu4+UnxBxsIch4SKJeMZAy0KEwqIz0E4Z6gE
EKLjOcbrULWBpY8y9jN5RTEKwV2hTAYPKZ0UTqIafREw3bXKcdO8MdOtWI6iNa3ssUPfxWIkDsPB
eLagD71gA8/qV1im+qiEhCuZnMOYNBUPHDY2IRY746C4xe4JOkMCMMCLme9Kiu26EBwgWzpqbJKi
E8pdathyVDqUhxjrN8In9Jj7qTevvS01bVO4Xubh8UVKgG4A9tuFgda5sGRugaiQiDM6sK5Y0SSA
o5tW4pi5oPbl4cL6AQO5b3Z2v/YGqZD2cfYLcnlAzlHHOHm0k3Qj3I7P5ff9vKLR/elPCc2vV1z9
gXi9Y6fTvwUmnLT9m03DgpvPCOe3fjwqJqfakbbFVSRk/Xn9r0/FdPQxcIpwXTSaui3G3iEa2aXl
bpiSusJvvS+ebmAr3faFTOmbZE2lHktFFNfcqt2BKwjzc+u5XZuluqjXdVSXaEaWYzbbvrwSgKzD
Ge9tnqKsaoDTXKgPAHCmhnOLKAq3I67wS8BXBY4xPU/Rq/DOY0U9thAI+SeZsIKOHhK8TRADwTLJ
fzWy0uQOtmdkCHjPcDjaTGJhChoaq1rcZuLXgJWWGaeWZQ6fz0ACHM1Qpf+PrPVohRpald1F3LC+
vg+xE9lvkftYnsStDilTiLPihKwHOWjtXaCD944dTpjIkViz3aE/Gp38QNXKxm8cPgBRVHVvVjuH
10PFveLvKBUuOaQAg/1SNEJXZG+tlPJtRo41ZTh7khE9bZiAIq393kxGQcPw4s1yAgqyhBdLQ+3q
d/3m51+Zlbxc3k1US9fL4yE7BvMVWBOdpqCbkRcB/EoZY2ZRSjInp3zR0n31ILlWFr1GjUE0/X07
9NZZ98KnAXvS4SwF/jNNLfGGLK4gQg7ynPU1J2mFLk/eTTs3ooxQA2pRYzyeu+6tsSxcBAXEIIY4
OLTtPKvarD05kFiCsSMgISjFdk/CZz6dQorTfbgqDe7hFZchrP5Fxb+8d4I6K65nm97p7kzRubje
oJ4ayAKLaV5hHTzAvT/wgXJuYWjdHjPzGQNgRO73MEOfeTajOnc7wSDny0qLsvj66NAjz7R8+KMb
HkLZNqeoqMMRSiVH45cD6Xz0SmJB+ruHj0etqTP7jXoV+8JjIQjxB6wN0leJTmy3y+kG5dEn8Bc9
zFPEMuNrM6s2GPgKBLSByHfeUR5P6ZAJOz0j89emE7ailxCzFJ0LvuHrMO/D71OdOnDvCGlsonag
Z5xySD+9uQc3panFI5D15deDENAwGe/U4h+KKG+1/iLK0zucXHK5tMu9ypoJLUXJ9d/AbQ5WCgNT
q9iKwS0GiuQIAZWxbAzM5Fe+95GcG1BT6wOStnJIQ83M/zyrggB73erdnG9iz1ZqtCT1eYz+37cs
wYOTmNvQxa41IZWxp9F/S6W9oIjPW1cN7b9P8m+xQJTuese4UeYgVqC6AWQdG2mhG7jhr/u258sA
txdsjwfWl/wg68dHaEpwliOP+hFHCvPhSmE5rUVF7EDPi0/GXMABV/Tun/HZuUXFtLplkKiDv4TX
jY/5aqKlbydsJWSnV2HB+1ncRsbfMjuTu0zOYA4en1+PAL66VkC87iuyMr58eRXmjfEUj1Wrhzpv
cfESBreReRgX9zpWqSjI5UpSR7lQouZZfwYdd9WMMelMBbx8HL6MlJaFa2x4B7BRySAzg1E2GrUH
oe71wsr2+AKVNsuyt7gH+jLp9bwALtBLQiJEWcrv1HHXLZFDvZdTW5+We0g0E5vPbPOcltp0V03w
eeJEorbMnykZIqR64huHtQZUoU+ZCh2PZyOoVLGu8aa/qpb4lDl0xD5pq/WPt6ZJnmqRoBVWzsOi
SYKq+dsLEnTijt4NDJd2F8VfKTd00/VUmLmNwLqgJZjEzdbi1Hv+4uwW57MQlc6NV7EM7IU2QOhx
JWbgFOnUpMBOGkWmdn3tFfRjl3fPnyn4VQ6ltSgdpd33wXO/anc7KySTFzDPPDwpzAfsu0zX+PBI
8N3qLe7PSVYF75QNdsr1AVp39r+nv/IyC/tsZ+eIfa7LwZWPIqLxa+44g3C1q4xfkwAFpckslWSb
MDCoY6Mqjam6aJIwpp52lZhe0lucyYq5oJPVYHjstKWRk/M6/+AzlOYExPaDLGWoQC4vFIrgrFZ1
sKNjQx6FO11qQjUM/osoTRk7Bx9qva3gGAL+CebnDD6zs+fBUQ6Rf3MA2Z8aQgPbvZz6ymoVpXHO
Qg6ZTFrRCAq7ceNfWCJKIiEqGBd3PgmuYO8G8Okb/1woMzxE+GkCK+SALHfWAMubQsxzs+IF02zy
Qk3UaxGdllfsbY3+6QDKQ+EVVyhQYYHoo8Th+GYR6plEFWCmoxZmnB+bDWjB9v48cGtQcWlE1EnL
Gn3WTHdc1tEp4o5xfDpj4FgpFdXu68qg3QSvuw9whRPy7/b2XOUgrck6q/jydtJZtjaskA8I7YJg
JpeZm26R3wQLNUfnbICkQXXRpULMfc9qwbd2ecR41hH1ZkOKFwq//8UKCbxlLNks/vKBhmiF8+RN
DqThgO0yXb6R/JrCJqZvIHtz+QtTGYxI+ELVS2/s9ohi6Mz7yGwsZSfLXtRasQIw6O2DSGEoVVqJ
tPtQ9V+1UFNZH+ZaD9gS9eC/Acy3JCks2OmO5J3ngzRmQ59tW0eAJZkD501Wv8s+eaBWSc2Wr6ag
NQ8UOKi0qszMcIQXYNEoh5NmHe8V15h7hLX4hgB3HyFbm1eaVD14aFt3zaua+D60NwMc7aPgm/q3
Q/3Rve2Fl9oX7XKYpcGlQO2MPpewAz5CLXe/vA3todfLcRi3RRCh4hw7895Bo5trIOVSztLW8rFK
c9ftpFF93rjZk3HSiaCRVaUpVFX2Xuhs/5qiqzlUF3MMqbllFBnXp5O05J7U6JBieEojP7LlCe36
8eGKB9SIR809pBkVXukbERPJcGlYiO8/0YLuw8cHG2OYuANVOKv+bJl7lpOzj1sA7MVsuZNgPms1
KnqqljJ1FcM+DFoz7Yp2e+Mx9muysbc2phx603kBpftZZqk7zmhMkCwWJPmdQLCADo+pynm+7+tr
f12TtMmTHI5AO3K8rBuGvDaa7BbMxJDO3DYpOiMwozo3huGlgFZU11Pii4/Eo4OLLaI7DgP1rh91
2hrSjG8sJ9hLQC/GMA8RuoA+ja6q4MWA1B43aOLPAIYxuKjLYiYJMdISOfjWnbZiUus8hSWjiRnI
Tb/LDSempxRcb1UiL8CuDepotW27JKTsiBIxaM1Q/fwXiAjUJ5VhnjDcc5gpW2fdiFl9c2sfk+rv
vbJLC2n07TYbfp0Ld7wg0LVSjX7qKJWvmgIEV+IBYgBF4a2r3fYKmRNGuu041spnXobgNedVqKS/
O23XPfXDZpzDOnFQ1J6ADcWVAiOKWy70sIuztr4225lUNiMlRh9jJFUK4P2U9yRkskVaVr11APWM
PJUI/ZAaD1envpj1hZntpZnLfB1YySXP7J9+oUI9qhs5RveHE+2YprlXGRoaUzWL5I8HYbwlH3cs
x5fUJa/HhdOREEeD2A0FlSLYxqPyVK5ehMbirHBcsT7bqJINHYwnYPSWO4GTRQaHDX+TDbNFX0wL
acCYDIZit/foVgY06JlbqmzBuMg7sphsiIHVbr0PPsf9Gg73PQyn1wSXyWHkYWCJN9ig7yH4fhwQ
XmVGh+8HDrJTzM9pbdGsxsWNnvd13mIXWKZUHAmsYl2P3BeKocvNgFy0AZZIj/FcXSn4+tm0Iva4
I8Nyc+Tx2i8eadCPTH7K29yJtGXOBs7P9fJl5jQSQxPxnpLSP6e0KthvO7fWIJ0XBMgYLHcMgDpA
XJajovKNSjh41aZeOO5tboFoA36uIv36K/gqatCXohZBycXvziwETylgyhH9czcm4nEQHdcjB7Tz
9+27sN+SBzSmedNBq8S9I2+yimqRSR0njUdBO2OojD+H1CNSDZHzG4s7n3RvCJeE09Ao0WQTQ0xh
MIZSDhxtxJILXwc23eMBvt4DM2cFpyQhDZB/PddjvkVE5YEdNVFuuGerhuvHlyyuPbGyEeqMhU+k
iW259VsHttVGJfFJJlqSuTmjq2s7xGM7V2SHeN9dUMzTazhu29xE0hogbow9UifuM9Ca0jSR3cV/
cJRk2M5l5GGbgcdvHTEhLhArOX5MQyvc61T8x1A/lqetUiWh2AOlJn5REzRp28FcCvmp9RbREbDa
lcn09v3mEWCUIV43vlDMjhyfmxnNMQKDailc4PDTYp4JGAKXtPDHfavRYBNmeVMYZGoChsIrm7eu
BZqZLeC/TMXAl4tU2i1vFJAHhx4T0LWZaqY2y7wgS8WrU5epGJRhxX/CMrDJJZvzmZ8PnvuzUYos
+Zg16x3310CXhTjtzT6PzSN/Qu8uOTpPO066qrQy2iyqnU6W3T6oxNWwOEhzu1JeZ3EuXuC5lklC
Bl81Nrookv+58TNlKH5P1tVTrgf1BIbrotZiF0PqQvQXP8l7JJGG4Wdr4v//l9z3h/vislPlbaFx
aHscm2G72tbWuTKQ4XgNVFWbTdrPNU/TvWVAV7Aq10gLtPQKIEdO5EGFawTuY/4WiyumyFbNHBld
sN6J6sIgf2tgFAGFYHPEvEbUicpuaUMaB59uZ/qa/F9oDv7Y2fIQihGRDJQpyQs4w370zYXkP2VZ
5o2PFWjk3vvxUv+9qT6c6TJHYlwDAmEBvApNYMkvFFFkU/KdNdCL3xm55SD7rzXQAKxK3uTQVQ3Q
8JlQc55W7MJ2McQfNQSwpPz9UeaxFFEd3b2wE1rxTWsRfQXngB/EnbzhLhRhEnzabl38ctcioWJ3
mIidj/XCI9BS9GAh6ECjY74S9oHqHtcUisTcmjcWtY7u+e7GLmwgVuLJFo+fCVySLS9a0OvC2IyF
P0MAC6kWAz4BXzLMQ/BxaUCHBAOuZTzA33RC1VR8HurM1os/iCibC+z3sVEG0+QDdyB1l/bnpdJp
eqgFQLTtaaotAQUzkY2SGW8buQRv66wYUvUYEnAo5RwOcSMu2eT+xDHIZSiaX+es03eszdZBwv4S
mg6+xr4eAwFDivSB9sms78h1bqQ7gVF/TahpS4rWNcwOp3naQiagOV0LfA3UlQwF9VF38OhBIqXV
Z7Uu+yUZCjYwMFB2sANly9XH2fkq2mMVp53b/Bg3Bp2tYo8uQB5L8L9aY4Sd+Zp+ogUAcTFOGexZ
zpRLDhXLOmlNHwUat/gYPlyheXN9f0cxRnYu0fKYSml1MtbFznAaygoO0eiUw8LJbDZh14rX9sH4
gj06jZA+7pa6L9eTSapVb6QOwk2Pkd5+DKr8snqrnTkVsoQ377uKY4QyP8MfWrnGmhQUZA/Jn7XI
u69jEQj01EmPzon5WwqFTO1S4mr91/IjeGJoCI86O9M6FmUsLNm5w5AkiW8LUIpjvSGO9Sf900BN
5n8INw4hSQPdFOifauhi40WukzZLqq3UOiGkgMmU1wErn17YNSBRvEkHtdR/4FrDHulWS3PAks5m
6dy0MVvoI6s73dtqaFUl1xepCIaZgaSOXrSIqJlgfTvIOWR6rBa2eVs9I5R6Q14iCtx7tfPEPfNs
4Y30Jf14gAJGJQWvig3Wjkost0e/DVGTPbB30ZcnUEztEY9iHkaTGw4NdlApZSc4oouCcmeMQxgS
/JvacJGwvMMixULWwqVkYyQqyF5XjutdCCXt4s63Veh4gos89JrfTUZ/w56sgstbSoEEfgz3eZbN
lnnYs+2rm9Qfm+JjebGaYFGFmoX4ZlbMr9GtmW52PMPqe1RXpw4CiZ6pNnfUVZaVwreiLz7KMnvO
gk/ovGMjfRwGAhxJSHutu/82guWkoXm+rYbRsjSuNnJcEWAHpClJiZePFo/Ixg8ADlXVq6v+epnk
OF2g+EVDR4//NTCTLpMVftCBJP0u1J91wBUjXkgzYPGEZn6Q2eVIqPMVMz7YRcCOK4S9b+aUgq2f
LMBu/EjoS4AkgILaGLRJktlaj0sdMQHAZdzNqXOgsMoxMqbzw+hhQsp1GTr6Sh0zx4uTBuUy5ww9
U1v8TGTpY/X5KbnGZh5CYL12c9el6XxeiUc2M6Hc48PSAqER3hANgcQmvhyHs9m8R2ya+JR/1Ss+
rF8dFZp/u4L7iRSa7Ruzb7xM767Q6xOS21gi0ukij2emOevDQ+DGMXfV8pvI+tjJpsEHDWI+7ZrW
oIKp9GaxnGVzJakVNy7g52hn/egU+vF3aNFaMgV5CJSnLalFy1WFeS4N0sptWlEkfR2bdxlOKLAF
89tJAmusbLF0gPPuacnxNsKGQDBViLjOG9vKGwoRMMX9gugDmGQwHBlp8ShSvB2xnt0Sci2qUKoR
Gjghl6Of2cccsYGuegphHc7/2lNUFot+ASc1AQMlwau7z88SpwDH5vXqsUs3U6deBPgqoB0ef62L
oK/V5KDEhAb2EbKGxgWLar50bP4sCSUqJ70VBSz4zskCRCzjswMZIqtWzko0GtVH+4kCYaHn8tzV
fTvQ9yezYJWR1nf+4bKiADJV0pEy6BVJnpT9mHx/TL+ss+yQZcR88fTTbHp4iwg82wvFDyZx4G2A
oXQxQxOvxPTciAxXIHb45UT5nt5zhi0W1x+Hb5U1DeLn3YkOh15vR7v31agGzE3vAmeKM/BXQGal
35ZFuxKFUX8Q6c+fbLyG9cgfuZjROTEqPiRUAknxebGZ+7/bhxPQLiFneoEi44IL9kEqbeNCK2pk
DJZsvorZJ81mADuMjNFAmOHA+8A4Rx7zfnWrrIMvTh2L0E2C12hAMO25JHFWQaAMQlZt1509UbGa
HTPAAUCXm5w7p4yO7iLHGoj4zcxPLVkmWAizlCM2DLN+Zt9rmT9O5x4cqy2Tkb4gQmU0InOMhCYw
J7CBJ7qG4SQz/X1e/oT40IJV3vhwjAUhc/Ec+zllXIjoNV+og/gmuhf+KuwJ7l8q8NZ3K/202Oh3
I8JgvXFCdv+0qBwwf1xPzJxAunHUAM0FCOvmjoqy2JXILtaSyc46pOxeUaaLBPOsyH4h5by7MT2B
jh7xuRjO71UmUGN8mRTw6OiGB3LoK0ujFrQntRmXwZySC4JClRTa8pKsYxVo28k/6mpuLn1B2wZ4
OCQl1dYKM9rrSPfXrfFo7y1N6YRiSKP3tesEHDTB0A35M8zGtP7HKFqhAT05nc54iNajSX1OrqYP
cdS0PjW9/iHg4B89KgBjb/dNrLdmdrfryPs2XD4r23MYtM0E/yjmn8gALQIjxt8DdQvParDzAGUH
nBUGNq0UlClbqmK+VFKOJHVwPW32mee877M1YiU81AAtmo8Yp+djOoXRw31jr7/lQ2vOM9o4Qxtc
OT2iv5PEecUnEPLXaJhNGVWmITWbXEJYhxKyGldb/YnbYziqA8Njfy9D6lgG6JWQAT0ee3g0FCdK
rQH95CaLqEApN9y/h6twp28Lqntcg0BNdQWQ9QoB1zzYsGZ/3RdGA1ytP6RGgsAhd2geEEEbys6O
We5Pgpgab6TqCPN275hjkDpVjgNA+0D1ZBuS+DUu9kr/Kspz54Vh1bWgh7nFvrLFha9NFhRWSvuE
YfMr4fSVS6EkqUNMW3JQgEGLrVwBwOLREsonv+h6Ys18yzIwg1lRm8MKtohyJNUaZyiBdH74U/Cs
yzqYD6QhXGH1q2J4n6kgYYzJVVLQopA2asfcBrXVVRxgS6AOXdj5xuWqtoIMCZy69mn4gs0k2pLp
ukcZcz3YjgX2VUQs3TpVkctsTL4OjOAfPhcJgRj8Pof5Vt1670tHX6vG5bnoOQaCsbSzXpMK/ADj
Ypbyh7XnOTwarylFGPXsCpp1fJtrW8wESCCOsdCOIVskt8bsPpnAyoLPZPu2qE1YNQuc9knUUBen
28zGoQdX/CYyAwq3UBKkW56vVB+Q4IEb5U03TYzFddiF8ipZdRSMpUFhqCfLkPwovtErCDvfKqZ4
66ko43qtzbKU4axOKMI4Lr6W5ePB5IqyadX9dK4+/lC7eg05gt2aaOAgVfqravHUb4WPwWpL1Zdb
3gsq/5pVQ054iGT7zLDr45NP6bPHmM+wjdUmH/sgVgxgF3RWgYInZmsjXKHy+QRlsvKLtqdSYA0c
U3sXZaLHzzsZk6kC8Xffznos/rGFIvD+82cOBcuq85FkBM7T+LcV9JIGMSD05PYQnQrl9QonftEV
KEmtin0gy1BIS7BXAOJhk2SrtpWUmNpP5VJJ705u+9d/6+YeVxqMWd/4ZoFkJoXfDrPSd6BeTU62
wOHXbSMOw1Pfjjq7IZvoU/wyWVJmZDSH4a77IpRxGgjde2xqmD1NTy4X9tx0fGAObS3XCYoulEVd
sjSV6bu03xTLnYRN0k62Zyruv+lDq9+POZQfpXrloJIskecrYrY1/tfmF2A/wCjJ4Igvrn66BdMa
p5vnoXLrFqBGJQjtFsVwBcllxJHcCsx7QZg22k6duHcqKkFtgAcGk2u+n0UT6lt6AkXA7LKbvEe6
HuvRqrj5tnjT9HMmwDPkC2Q/ahKIgt84Wf716Oh0l7Hu7qQibUvUTu5Gi/nd6ADT7n25PkUqHbdl
+2JaIhb0UwwAvZgumN5m3HpRsfKuX65Nqou1prOzBT/kyH0vmcAq1aPyxGj39DH3i257WQnhf+YB
RmL8MMs4e/SyWEvrXVBWdRgLO+/YOBJqSBXV/ZaHxi0ud99KcB/VWtkL//jB2tkCQEqqbyr30cUW
88rk3Q98+oCTbD8oTD19qqjSJNCPnc6MeUlm6HDC9bf+gVBBRkwTbG8pAjTZmZeyTao4okLwPnl3
n/hjodmUq+von/CcxuGafRT5FUHG0IiNGERbjHsCuNVpais9uDVw/vA6anzYUALiDqMJD65eXH3g
zF0+mn3sGemf2JHqgdYsUUFFH02rpr0sUVtnJnfOXP2LjwiqpS+Nj4FtivR5tatD8lodQ4dmxQ8c
aeiq6gCR5FSkfD3xYhNKZ/1y+QZGwJEjNnUWGL96a4Fr2NHKstOonEcFqLEPl05mghQTbakBhsXc
97u8fIcX6fvTRxu++paidq40NDvsS9XXJ2mAuuMzwrrql7Hi141c7STjVm+alnDjguqgBrJ1jtdh
vG/2PXtL6tesylml2DDGUkz7A40/j8cSOcmHO908tw8KOn2oHxt5i7BaBUKRL+zZbX0y6WVAEWI7
G48aDX4uazu3HrDq+sgRkXrAHZ+VHHoSUCB6Q5AlFcZnPbJbuv48w5fS7k8N4yA4MxFDffvLLqit
LnPJ+CndwCYHtJUFCZg1g9J5UCbi1Ef1mDm1eBPoxypv6D4Xc9ZbtdjVE7TqkrjeUuMiqTOLCaW4
D4Hudl2cNlA2bK4TCDZzRdPBY7cehqj4nzWYU9VPYbhiomGti09D3uwKGq4hRRbQz4U8xUF2vdVP
cua2Rw03W07w+Us+YUF+eUev/gACrpjVQU5FOun0QAmonhrtWBW4crQJ9QqSBgHnMWHdqwSacoPO
jLQGB8NIiau0OPld6FPTAWJ02I/ekYXm3ghZBbXmtHLWVFw+9W7mNGuVekHOeBDQs/Tm1PTN9ncR
6+xkWUaV57On1kHXWKeMUiVbj1k2EzyxBLew16Ogn593+e5p48u/yHi7BnLk7MCE2KETrT+4OrEn
ITSI6sTDYPW1QdxSSBDkVUS5Xeh8WSTsXGKh7Z6Wy20+EwBfXNep6jwafqm5TDdRbsYBCfre0u14
7KNyEIwRBJtxvkCwcu0NvUnpO9/C2SIA+m0+UueZnZssEdkq8u2Q9y3mGxJT3PlhxiCY7laPKr9M
FZap1uLOw7bioSiCKqbyWGi6pnkFpn7zNUimdJutcJV81whUdG7DzTaVipyAOYbIrpkF0Wn7Fddt
9DFfhnzkV7SIKQ//YYCatekVmnWgdoscxUz5fvzXhlIVzODi9XWEAkPf/scTYnJD5SGmnDXW0t0P
bwwAuy9YTxdVDxqTKzCEsnA6pWWAaQSi+OipSfy81jQMc2ZvrFsRkzeOMRKVHpVXuJC0ZGASnsFN
9yAui8goYZXrbDEHNcjFYf/5LQUeM7qjX3dFkVl01DURlNcHo0PuiQE7iXJZR8d/SJjym8BFSlWd
DLNYtXfzOmV407mL8Ed7fYUhnVzcLrAYb2FGzca6rm/MiHoBjAfMiuL1ooHwfSulNIb5ifvl1BlO
j9h/AUpBmcl18c6suErBogJ3fM9FCuRmnZRhUZACTXjOdm9s8L3GUIWqmVHVqYZLoDUKH6kKfqsz
cLY3YGSpygmKZfB9gYu1KKhQEsA+bZFacyUOWAA/Bf8FL/Go+odtolrbWrAyb2AyaPuTlZc3JPPS
zjt4WKGM2Pi673FJKrS/2g7L6X5FUDIoxN9Y6EP8qmCxW829O7CSKCRI8IOx5guMcmZW9virUkLo
ycl+wTt4owkM944zglYePYGo6jhd9Ncvn8Fr897RxQOIeQUBL23ESOEwYHs3zPMCPU2UWpQbgfcJ
xd/UgHBUPeInYbi1bdaTmcLAPrGVU5ARcfpi1+eji70Uit244vMGu3er/hb26jWz0d0ok8cMb80L
+eIwnRIqgOaRoz/ogX4wFZktH6WOh5C8A3RNJ/Lhc2fuLP9hWodjgD3OSbW5Ityin8EoeRhcEC1e
iQWO4pjeT/4Y9SRyDrz0pmoWN6/fNGRSI1j3rhDV6ZyFJMuGWAGlkV8+QiW5qHa26eYy7cE8sb//
X4UaicagkStWaO+E6BVQ8kxMHLaxZQ9YNqdCo/GMVMc5LTAolGzYL6tUzWrO3LS8DZhgcCiOv1M2
n4kvQLpJA5lRL4HKMFs51ymX6Fp4cpes42pSjZzIRd7RLBoSAa6uv/P1UDKy6bcFpHjLgvX/8PBl
9x2JBdO145S3fuIN9yvwiS5GFA+eBTYUX07ksuVMgtkHsbdxrxZZMGCzAkziGFJgpSjZ9Hu8EFrQ
esoObr9JKL+VPNZTuhde7PiAYN5wWSosjkaOrRHN3AkWtEA/zEx8eagbKs5gRoEmPso8CkT8FL83
8KQGCphUmByGnq/kM1mOcIOAt9XxcI8UicCQg4tKgYSn2nSc5SsXMhQLnrz4S61C0zIM/f1wQyTI
bg0bCDuIDSnonVNr7+gOfITxLd432XPOXJtGBqkpTGGFNNnqWftqte4weo66uNdFjWSaFh8k4OWk
tgwmDgnfrF7/TP7HgkGjPJrNNbVQof8z8xOIYAIi+bI2oA6d7LjVbeRFaCL0es06+XW/dNs8a8MH
3IolqeGACMvZfVvSulAwFUd/06SDFruq2QVdoS4iuLiPCzhQqR7V/dEIHaHVnbExNY5mWEjijaDH
xSNnMkgrohaAjvAVxq+WJpY2WwZVjls2J+KcXOznfsl4/FwIc4Go/6KlvltN6b/T2EGQM8He//dR
9Bj7+3NfBjhpr2RtC7CALVrDekjuF0tLxIFNCSzwrmSm6pqqgyzSHseZV72WdgW8mNjG7Wa9UQ77
TQKCJVQaM42gvVsr5gdmy+e4nH0k/cA1fqfj5J7KH0+GEpysvIggF1H70v6Lj3bVxU5pROFZwLGR
H7mOxQqc4nZbFlh2XGCvImNjyuZ29FVUu80iiSmNND/5oGlTVFbJAre/V6JqOFyvNxUinwexeO2y
/SS6Om1lb0cfjr1rB4AVCtHgYj+va1JeZbNJrUjDKoRnXN7ELA2m+nkc3jpzpIcg7SABQALt+9FE
WBuS+AELuKvdOCNdAx5xKCKajaaFlEqz/xSgr/DCVp9zEzhe1GeiAs+SJW2QT2ghgkG335aQUsky
PtyekYp/4k0o0LqgBMX4Jazh4WhIEHPl0n0gXLmra3toage4FVge3o98Ahn8lCXAimSAZzhkNtif
h0UtWoKM+Tz23/v8i77WFIpyNPbD9BEjHHLUjjC6P6B1oWrZzRa9TgT7o9aZ7MSjJ/L9lkGygygU
MxuEfS7+SSOI1HTLBFRgGZzW966zM3dVEkHY3HVZxsADqKWm5QgFHhBoE9a4Au42QzMYNrfsq4IE
UGOxtt154Q5/RlQ7kPkMcO1L3xG8rBS6ofY7h3aEdo48/tzQ94m78q9cp+kIP8vhVoaLQDbFfyYl
pgGT6sBAFhaSSpQEYHqXwjWH+0srTHFJUa84ufSNzkpTDq7z/3VbINEO4e/xfuklOL7GJOisHBn2
8u5LjYq00zUOZQK9crLs0zSs/A/2BDfUZfLurrIimYFcl3W2C5gLyPtYlFnwaTDlGQLlkeOURObz
ETmQjsXbd6trw9h45B7EdCCI3EOzyMHYb+RmeyyZ0fzit/6HalRdilQAPFKsMtDh3RGiUwDlx877
LdDQ+W/Ky5V2aQyB4wo8jMvY6/Yj6pgE0Q+8DFat5vTD4p5XcXTiqwfDzaM/evG5O6OaV6cQyf6i
/bDdiK1lJy1+5WuMq9sGLROnGs6p5cEMQl/fInzshxrjWxqUiGlaB2YvFv/xKr5hlrGNevB6Vjk8
5EThubK8T760imBIIvOJXbqJzIiVoksjwkITjhrG9S9z8PRLbtUHrGBe21E7ce+7Xtt2Nix/LCov
CSfjY89Da2QlsAPWnyZoesxENrzyglPT8QGtx77PimYW39L6sJD1WkatbfDCCQhAu/S+EIYOG2N4
H79OqnH2SUrviWdYzA7rGCi1fqp5OuIlni+lK8BD/UKfROoeJNYKqLql+dedDk05srayx1VYz2vm
Cxt6gAEebXw/q0ZQQRl66nbGKIwBxyGg30Ap/ux25GyQYB7w9sS8cWcH/VU8kpu2BYOUjedQY7Zz
CHAux9Jv8gvcSqYAbr+AdQdUwbLMRcvehVP1zPRFYlkFLkYNb7jApKQPOqodND062JWxZftlEhk9
pyPwnjnNkVKyYZ5lAx/qXwlFNJ+jFqSUTW2NFFQetqUu9hAQjMk3XOsZwNC2OAK2+D1xUPAFKUJE
WJMYllHOCLXs+a738Teb55iWvCRY3719wd6guyNUi1q4iwInkUNsbwd/SRs2D/Ju/m2ea+HatArx
NJ3lxLf1TrWYwIbx2iItQ/qexKfuyw6bVLjHiyGLMyxPYF123it/I0p5cPOB484ybAInUgZ8qwQl
E0Lt1k/XNHLSg5th7HMkh7ybmgHagvVcSa8JrJ1SeCkjfKK4sildwe+dm30OEifi5GFYsGBs7vQb
w1W0fy8LhMsiiSN7A84K5ACGFiQDUBJy8I/QyZKkHVCUwgN+JqnKexJvZHd5TK2SWCVugrpTE4oM
hpMUe21uJQ+ETenp3Y51kkhATWTrpB3EQHnXFq99R2Dhpi8iZimqXl9JrrQEIx4UoEezroS+RnbJ
ZCR3R9uK68gmts4b5lgcoj6kTa5mXThEvLvXGUM4rj9PhC3g7LavfWmcp8wMgnC208rbOrqi5xc4
fC/LXGkiyMxLEvtqQwu8Id3seigEs3fIETFRI+5jtsL5rl7gTEdCACGWXG+9MuQW5efi0TmmYR+L
/novMPSLEiQxiKLlYVTh1g6aHWtGJXdtg3oDV5ijyqAZZBI0VxdhBAxy11lDLW9n44zxMR4Zr0FO
WUDWo13pzuRchM3pYnofh/BUVDESpOC6m05FJIliQkDsZzSvTnNtlxroqb9iTYMnCBZ3UOsNQP3W
ZcYGdaQhgKaFBqqANDRNUdhpxU7MSwgvQeyiaXlRhLo+fBPjMdCs+tWltsSRkZ/MhgqtfgsGnU2M
qxwtptPNbrwS1u+S4Fwy3ZSqb+ltdds5y4Gkk6ParHDXJ3fiAeBYoEzzB4paHxIblRw/h3MTkLoz
CyCj6S/mw5DCpcorF2lp1KVLUCg/giMeHd1jbov0/dj2Txh38czXPlSerBax+8ZDzx6KEyLtTtEg
mlSf3VURuxxnPNGsNOgWhsXGP5+YZkABjJ6lFHy7WMriSxTTFeSYXzQDvZEw6GoWvRrKETr9kWzu
3jTiNJ2m4yhGkDcx+1T8pTwWscxknaFvRnfzrvNGPNsipqngmPSH24FEAVJAySIfpd07SV+rVO2N
rHKSaNoI+Ged4+WwZlTX5KrglHSFYYtSD4Sq/bHEBeCf/Nhv79j6NtHq2UluK89dS2K6OYzKmCBK
RUQgEoAEUaAry8SV76/YMVZJ7NIQ4FBhWKLcY96wzpQA2HSIuwjL8gas22jJuFWe/skF5vKR3miD
zwXlFfQTtBHZsQ0Z66iVaZv87O0yhYIpELt8uPyEGSc1IUsmywm0OQyn1y8qdHvOBhOh8zTCQVPG
BRLFlPbF2xUiM7U/eCzCPrvvxe2RwhLLAdp2xORBtGp8dtVSHvXS0oHmXytCoTFWsZpBjpSup0iD
rtFdBNffEZGFgjZP1fwFBzZS1MF168kbYSGEDWkINYNckUSLQ5npPpjPuDXQEYfwBJ54euHNjdhe
DgaHbHeTKOPYkmoE1UgZd19swpS3HNBLVUSDQawhRsdI6I4oI8VSzHxeRB8kWh6z1a4bIy41CK8b
iNCiVsiRRCd9gVWLOTBsI9trks9wJG2c+1H/PNRTokvYdm3I20IwKVJvFc90534AgkKBoEW2EILr
nupFvGJLPFn+/8G9NljGdl1dEp07fGkg3rSBaAQWpJOn8cvJnRjyQ4kI+O3isRb3BVr30Jxa5LeX
EqxzQ6BEQMruDjIsrE3lkyJ2K2qb6j/vTps+5yyfMIpGcRVr2dYufuoHjj8cK3KMBkgE1j2sXThC
RvZ0N9liMRg+gYa8tWvhD6G9CY31Bc/qmRL2NydT2dUXQCuDf3OXF01MSsLH/1Ud0sQ+B2fSK3aw
wqBPeJnZB4HGtiJ9pyrIm8/In7OoIVHor2rDSaNxlIOtHmqwU39DIQKoaaMZc/p7YkurmM1d/EnK
lk6TTDzst3oIgCtq3N5xhcyNa7Yj20O+sqjo7LqzBNDMJ/2M5slPa1CCEj8lKhyjkqj8//Fw9bxR
T+//eedTwQglz8ATSBEDMMEduXuxiohTyNUjldTEFgN+I0NCUuM+25amYVECCsdGtJ/kqnXPXp+p
PXop6LbL4DuH3RC1nV3P+dwl5YnBecc0WFMdBGyUCCQuVZC9gni6E2dAuVLuZ8obh7lWd2l9lyzM
NjR3j+uOi5Ov0sTDogXHm7ReJdlS1/pWoT3er+eNZQo0NB8+QA4ikIVHwoHCMc21XD8dzNuvdrux
RFB3aMphdllNvaiKG+WVsIuRsVcWFlR89Qd1bzED92jv8ubqiJRYZ+Zu30xGOh3xmcWrBhsc2qJ2
RPlBoCx09AsoM0ztZr09pPZW/gZjur80+18Hil+DQuwvhvYRdCG2RWQHs+oH/KzQKYahRU1k5j0+
el1SHzqJYUn2knz3cNoB9MiAf3YCP8c+HfaHK/GV/ko08PhSiyYIGGMzAZqeaKT7hndNHU5S2Gbh
O0nM6TFnAPBUbRqYqKRO8jLLg8tFeimpzjsYk5IXd4xfROtfgawrXXRE3uHsEJpElXTzTh1l8ALX
9Ex7dSQ/+WKV7L97wR/BR5WmatOWzZzM8HHa3xl6iDZBi90jXPVXvvF7ZoV3dM3VONFIzjy9Wv3z
fkVngrhvnbvzuH0L5GEwxoEqVGkAfCfVn9CXfB/H7v/5buuKsEKw4AtTpnTOdbVvKViQkmeIIGkZ
291HoLgj4lUgUNxwTuv88Qs0PNbdsPaocOt5RgYmkvdbdfb1KsTqoSijRPiNmTmz1omVTo+FngIw
9aWNs8zXOXqM7xE57wirhbHEGlBv58Bn9blYGdclJ90/GPZnfRXj2ge8KLKjCyglDABInyhxtIKF
HYZPhKd3CuVLD25Ezq1PacfDJzEodUUymGcf1AWXYzYhHUCuvmB3Gpk8FO0LDJG4USfvs2CHZLXW
2DVscGR3+0eKzeorbUI4PQFgATTDCGnkCQh6seT6b1rQLNfxOMzZDpcMBrNE15J5dZa0At/vmZPu
0tsC8lJ3ADhqRWBF0C8xdJeGJqoiBzrpHLK8pEkG0bhZ3KPu/190R17jp2BvBlfSHQatW2V4Cf5J
pClS1zHAOo9oqBY3RiXxOExjmA0naw9PhaInoVzZgAzc6x/C3QLZpo1aSv1mH4jQIomGYTaDoLBa
vr0l828dmuWoxB/YRueiUKV3a7x3paaN4LYE3S3khA0YPtxFfx8UhiRhCKKvTswZ1REMettErwAD
E3E7rFeJx/ldzFy8ez0I7ZBaJ8iemq3AnWmBRqC9SdduGFLhCKfsrtPMjPGOJ5RsJGqf4XzSzl3S
bDM29YGFd5nuag6fQFW0kWUZhjQCFfiw1Y+rk/raTRQkT2zarlD9t5v4Wm7hwrAw5ZYI23H4EQO5
oLlIytdabrfDb5xTt/0kKtfeSNAf9JXxLck3jeolE8v9XUADG0vcUPnWGLogY+SfqznBSYdo/W27
UarqfQmPK9apFaPYmSn+Y1EMzWxtzG1K8To4dWmeYpb9+bqZM2J+JN9Z0bTTFbmnSpuyNuU2mqxb
Uf1RxQanvIA4llnPq5mCqOaXd11/YzCm22yyU0QrmUdVlN9Ru/hupBVC9geX0l1+55fefYDgerUO
xuwmXliVUDjYRxmMtA3H0nyO+7hfFTUn8F0tMCCdU3J9whbBmt90SiGJZ1oBH5bTOK8VWQRzOgep
mVTNKa+jW1eI5ZZISpg8tsq9QluNV6F8XQarmGVg0qGRp9ICs4t+zU0ZINMrdlspzsbSVfUtj7BD
sCIg+44i1ARoHqpACti3YPrBOYbIaX+vY7c9iTY6dePuj9rlNOi6EwMSTTrWAQPqhDmfxDkOp05J
ZSQ9DQXo98jVwfstjfN2ZM2/lr2B3tbz3LjCi8w2xyzUwFY6AJJv+ad6WTNbB7sbrDxGg+fyUYni
LTIVUNWHqSh5hj8u/JDIdGt84WMn+YIIspaR+sljfa+3CPB6E2faRDuTdqWeD5vbCci+7+DcqF86
Qtv+GVTEcPisRc/u4NTGuchDoHltuZ68oZV7h5OOltvsa4xlm8tOo6GCOla5HPwsCok8mqS72dCt
q9l9XXTNWPteVi4jHh+wjIujtpcL6HcxgUH7tedCBhCC0UztPN5xrbP5fGy4CxESw1MLkMS8sPGW
t8uapiJmZ6hEmPDDOFN1x+4btN/fVlGEFq0WFlhVgE6CGrRvP9SO8fT+67U+PEjD38Zk3ls8NIcG
8GEdvGXgj6cJwuftQWdtzeEtvQuxRnScGwN6XF4hMt4L97xrchqdJoVUKTn3+Uh7MXG8oeVNQlMd
Zev/25qS+ZC/9mal8BUpR4SjlALBeYioYGoH0CHyV6Wiq0BlsTCVXLtDi/7ShQu31gEKym8h34DD
5lW7PIkkt7GzEZkLUV4QLvffYnStsZTmf7kDrvV/ig8Adr0Xu1IpYxqOJnuZTybtQQB6PQHvdU+/
3xZZdBygwtqBghBZ36FVH9lw/XjsUOU5xtTZRUre+3ljkJf5xHPWTbV5m+7egZtUeVqdfrQ49uJw
JOFEy4D/Lr/mLcwJoL9r4zUNKdCi2rwGv6K94yL2p+yJt/RcObsT1+Soxn9rkMPFt8C0kwlrhkfF
aRCyXkt8eZpzc8zYkPJGWUI/vz+lLtu4kXDaEawoVy0vjO8ODXI90cYLh6RzWctGln1CejI34Kby
lHd3xMcTka1G5m6vMWYNgRFTQ8MmUNzldkFBYCMUvn6qjRqZ2w0dS9j3Z3Zc2H36FJJ++YAVtdgL
Ln3c/K0Rnt0oRrVVdHwrehTl25CbQggOK14h99POnm5VFbaVDQ9wbAX5f0TkM0Ts0zirAKTCBO5h
Qwt90/HxZC7qpER1M3SXVNhB6n+VXqvlBwQDs/8AkdW6xZjJ3DLKk60RdFaid5dewdSgzZKmjvCx
atQPmffG4V2dLeLWMlCseYVeuLNCbadaWm1/NfoJw5ElT5KAcHqX8A9mUgT89ZwjVIzRV9b72iG+
Cdwpky4F4p2V7pKaagxQZ9ZM6uj06RtTA0Ia+IJmsVFBZTQzy7Wf34w0ubNY8Hu4wbzMlSG96bBR
L155NX9LNEHeuppqjPRstsIOi+WA4VCOJHMS/wFNjlhwwMDqn4Zglh6UN8mwqkUHDN/4YotAPFM4
BWf/tP/o6grGzSD9yGTeOXFszurOHfKOs0dbBjoeI88kQU4Hio49dv1yi0niRNg+v/pGwWd+s46u
FIFOpoo8oUG0+QDY7xlcMc3kS4mZkLm5o03C9Gk7blMrIGD+y+Wm9guU2FkjPpQY0KvuKmBb40v8
0JSNjX+4/Z4cEYOP2a6NA25iU7hf0c+OmIBwyWfJm8PnvOZouUkmuOGh3S7Pmg0b31ld6ZovOEw5
RrwWL+1KJGNUADfai+CPCL795NlJbBySysHWb9rP8d+in+lOq2OkeoEYExjgAk3JaTgue23Uh8Wo
fwPoORXthNGzSZh8BhRAsZ32+GVqoXnGQAZP5V/PKMOV7PVBzBnKRV/ojh+feLCxuhPiGVbGL8yt
LDl9IUa1YonQ31unY4/aazjwd9Jk8wVgPq6hlFbEHxheBv3EXLWA5LWLQ/KQEsI4/kjo7edwwKS/
U21pOupFZqRif+9BocxXtrb3HdK1u4CKbg8e/RRLhwu7EwLomRAaDINmIQ1OePvmcpIGOP8zQb48
8YstqtUFBZmVT93YhgL+rmxl1dSuOi1Q7D0+BADFxmTiHAfShJ0p3BX1L/nZ8MbZcEi//14E6BNd
QirE5SUXk+q/R3Mc3J7RPJFXLg+4QVVMWydKcfeL0T3UFV4txrC+ISoNLs9YlxJJV80FVlBKEpVP
HImrQGcNWKfoYHR9tWjxfoA3zMKJ4xt7SdvCvYKY6GGCc2GLSFiDwLKgLIbp3+1UfML2oSJ1JEcG
BqW31anjq8wWKJaBL31qLo6No4Ex7yqGb8WRHhXR0Gi79A1cbBYdzjKVU7gZ+1+1T+Bfv6RXHnrN
xeBFMw4xDiirV32CtFVC7cU8ZQY/L//4+MqqjnEa4d1Y+H3ihZ/wETX2h5EwCQC5ung2nWTB1HRi
lggoST0KJjBAWyGWVLPv3tRIl5VEqeztWbebxHTPEYzEEfGAUNDVS3colroNBxDy/fO9lmGayaI9
c+OBnDhns2qSHtbk7xAaFuRz5s1ZcmQUmtO42UMYvdMSgpdF117FP2oTMI2y/f6ZYE1Stfa5/1nW
50yRaMrGVczLl1+BAQUGdUoWdhfxRBEHEVoGUJRglYOtWn63dFfaCDActMuYzAmAWSiXRXzrhJCR
wTWCjq0yf/ce7iR+Gzz3Vgw09iknIZgHYWzJq/EdWiNCvPH3GDMJdf4ykN5WgVFD7WJ0XeWJxy9L
vUHxQrr+0Mb+/0aomQorLeiDSdGkUXPdVnu0Glo5seCsslWp6U1Eanave2iGfE+qS/2PZYWwjeo9
0q37HitFlghDDjn2tx4buFBrGqTkh4AfEYCgTQbGjzUEM6vTznGX8oOaatq5dqTwnPejZmlBhsdA
MtIUz3jycZNgPod7iMIa2X5rUjjxi9MM6Nl+Wks0AXQTQV7kWbxfrsHPzhC48+O8ROIci1Yx9ahq
N9cNuvgfPMVntTeKSQkny7yDzllL3R/e7TKByWSRZDftVgJ+GjSC9ELZ9yXQd9k2D850aEg5D0hR
SvaJm+BNxMPWH/adVyeIO4vibXB1wM4WVgfXYCcuq+/kjaZEWP0khcjniiLKAyq2iMtijEoVbqrS
ZzdkUu10Ez8eS7uxhCXuXdizckLi35N6jbJfXx2LjgEeAlURGoeICli6Y+BJk//Dryfi31tRZE1f
I3miV1KzktfCIFctMlfv5cI3knE41EHGgqUZpvqlqRY90rD5EGvHfFn6dfzbB9UvPhufxZ42UKhh
Jh5+fEeFCytMjpAzMXAEToBps3n3yXZxXJhMSeaaT5BU4A0q43aZy05VNJJSjVLULLrv4M72lY8d
9bA3OFVtHN8gdq+96YNO5JMqYnBQf9LacfGjloSOLgUxMD7O3G6z7IL+Gx7YOiKwGpuH2HkFfErg
aTJcJ828jXQadtipQR+IzhnzmTPr5HtfI0Ntjuv7ymTj5hf5HWkqtOkk1UKuL6QlLmN6EXRTLDoi
JF2Io6pMoVrSN2sGSOn2lFFaANlG5URFsy41+Ywks/xqHb/uxUwRpMNEcI8uHBLMdNWn1sizEJmm
euJbX+a/lpMUKfLYTeT0eTpfJWWVZX+FYVcAjT0sLMr7HCRTF93sn2k8WhMkltZ7O0AomMxUu1it
iyM9mAbUxmVTrEgBM+PUTCSunte1/HbJBSD8mufCgvUHx0oHqBIcLUDi373IPswcf2/iB6YVztOY
peMQZ1iZmEiTsn31Yi4LiOLMjerxbaiVPtRVmX52CMDhpd850ak90NkggiPH2xyKcqH0SmHTnT0V
tB9zwTaNj4owEjNA3PVmR9tNgtTcjzuOT8eS5mNJrsKIO6qY/BSZConAj3DNPlrUvDhvmsrnxjX2
/+iceVaorXZBj8XsBlyaZ29HTGYGzMR86uxU9iJZKGnOxykedQVND8RC64+7SxbbS30PJPGmFm4d
rXFWT9Kb6FQXET1ZS2SqWcLKBCnrAdTTB43AHvkZyPscfP/IkbQcaHSm/XR9EV6sBvO1llMUhHY1
/Z4IA7puWAELwD3r+FEf9IrNfe6fwiJcADRA/OsmK9AQPg6MbLibwC6UfbTBePYhFystbj3iH+TE
FB5Fp4qNL/U44wwTyv4LmgHt0+FWPuwB8U3DqgtbJfHbXvepa3YU7p4sxiyaQqpAsPcl0cka4acN
78JiE6ieMBOwisaa1akmt+pE0ysdsPAXB5GcYn6Uzj10UWO7sqC0dL8PBXZrF2zZq1a3Boq6utjB
EkIdroMGF302xQVRgT7cjl0MI1VO3xRVGBlfQsuYEkX6ypO/FQoWJX7qQ8Zz9xPdV1kIDYlmS/8O
+f4C7dGDP8Ux51qhr6Bhu3ubC81BbcSqKyEItEss3t/bWX6Gf8Mxi8izDK88d/SRTiZyu46Liink
ClQZDQ1VHv9RNNCCD6oh83TqhD2s7O5EtH/IkQdHgqmVOuYcQLZwlNi+DsZkyHtMuv54+OYjhxHo
/4j3FrwsTAPZR32WXUCanlrB3vhalIkTcGQmZaqFQ5aY4t2/VRGeF9Ucl9ObZSC6w6CCxYPA5tyW
BQRuL/5G5x9+vNG6d75g9jubwBDB4cGVhYXn0zPGKLLzUDzirpGeKyQ/IKVS564VaoEXoxI75WH0
KBRP3pxwR01OExd+PBmxkqxUnP89vOdbvAMD9Tddae/l/oejY5XlyIw5hgviTYM7I95m+j8rtn5B
DAro8awKJF0GTTHhBQ+OoE3L/i5mWwbAUJr3dRJucT9f80gEMTDXzNRT48xu+w6ofM+bVnhtCl10
84HOUEswClktQw4qTvyloOZbOnJHSsthnyLlgdjVRdtD7IMTeMjrwOzoFDBCCRbG3RxiEaFakEQo
pdFgBFpNsObohU9oSG6niroqLalr90CQ8cxuXnvXcgOOnT+w62c48+yT1ZirJR4QQdhZPNEyGbt4
nG2i8qrhRdJjBvGngI88O+VMd41NAGF3MyNu0CAEUgjmzV0ScvVfrHxwMdDws66ugExot6Egs/gt
aGy+2V7Dgklxpf47rG7dUejSk4ZYUcRefnYXkQy7B1LufNReJZEliFrkCS9+dR/lVVRqkAMQnyG/
OzQJg9OPlhJOHs/9efosqwqpgvRbzzUG2aM/f9wJcBORlq5nmMgnN1ClMyjVkjvVDWQkRb3eqWgU
olZxvaUSNPlKx01ecVtr9p4h5vTrnuLiG2S7NwRD0Z30bikwypkb8Kh6q82aZJHBnpxbHDhvzDAb
2eimcyUb1eUKuCHEvS2wGI2KgI60zVjpPSJyg6wV4tWKgi/qTUgvE0CIRlP7CGZx9SONT3uo3gOL
FhHfr6dI+1hYqGfaeuiAMvkinmHItnaymZ+fVhsSNT8O0UL05+huqmy0qmPMpJxen2lZaRWDUdhl
qyoDZcKmUdZC9co+udaBzZpZWBMSnbEfNiJH5SU6D37xfvGdN59gIi2BsiDbYI+VpxlBKcWCoDsU
2rC3+zd5+pR0ZOTejmDTlBmsG8QcberSoTEMCOKVCr8OxOfPN7kkBjyrFy8Rrp4dViU4M+mfgFSl
jp9D5Kdv47CJ6MyD0BApvwNsAOUuoKphG3gwGc02iDuDVTEDD3HdpAbDGp4bmgfJIZJvUDxplE2U
8xasmu3eLafD/N/wEldv2G9CUFamhL6Mo7yNXxnvZue4wGwAbCr8/MSDAs+EApIzNulYI8aOOFYJ
snPwkmeZTzcbYwH+aFLZnz4n778hOrY4wOzfEPyuTzBpga2BiLPvSlw19JXm1BZv+GwPcmfSQDs3
zuQgZPbrrhIYkgX0LA7Hk3iFvPOBvAtLh3efFn26O+rYkilVD/JNFQChRMvK6Kau9Izst0dXsTcN
cV7n8XWttZDvpn1o6jZHbfTziG69KJ4g4Zt2+tnrgRE4j5a6kdne3OzZqfn4gO+AbnZ3/FLt4eDX
SQ6g6PrjXYmkR50Npz7cPn8QbmyxbBaC0tlZMklkrK8sjDIp0LlsqGlKAVvMBOxvSB3qQlJ/OBSk
cNeSZlhoWyqiZQBaVeNGP7m5cnNy+0wcG9msOv5RDNd+FhsGeq2oM/NytvZcyKJXP23e6F/xhGOa
3gMMwkUxq0pvmP0i7nAe4dlSpO/+mfdSoh660+yZaTph+t7HuegCZvwlMO3vDhsDWQ+DyHnzgAhA
s+EOYlFxi0jGnRu6oefO81vc6MYPO7LElsLq5sHSrGyhLTox/TCIjzNX14fns7hFlrHY88eVzu8Y
52CYua1YVfxYV+EckYMZHxQCut+WudxncZ4s36Sp3FD7Aq0isKrkLCi8S8wl8yjk7ZiTp0NOZjIM
wM67Q0gvf5poDIxQjbjOGdRCmSaTTkM8qQ1Stbd0XD7d3V16SnrC3wwf/Y2oFUyFWFj3OSY9WSbF
knQrxOi+m04A1E20Vl5VftUeqC3YzEdjGxuQPpMRgzUTAg3ukPh2kKtHvZYaWeY1PnPh5zEz2XTu
n7/hE6EQU7hFgJsS+8MbLeNwkmcaezdaePaJT6ttfH+ZkaL7Ubsqni/W6RIJ46GQjA0atet6p8EV
o4F/3nfdBpkCVYu4uhHvXwp2F8pxCD67miRx1RSvSEky2uzlm+mfM7FSnn102H6rzJb/UjPrYOl7
KExTAFaad1PZwJx2DCO771gviUagCpcqpbFcyduSGWNp7gDmVa70nGCCdCxhBDstrBW2vNjTeB4X
mNxHeuV6QiAjTXcD6pHsWgoSNbGZNNNmr1EoQ8iGj0xTNyVw8+8O+5hcRpnkdzBMxRqPvNBT2m3v
Ph9MoMKCun2UvKMcDsJ8vJZNwwHDhcKKWHfOLf4civM4J2e0WaiJgPYtT//bLe8b4L3tgZVqeWT2
6nRmsOTmJjBh2WSA7Mvmh+QHnachRceI+/CUPefCaful7JUdsaLEBN5ejJfgpGuDy3BGAU7fpXt9
RFwQ35/czprGL7HFa6bys8enFWUS2bUUiQBzPydYf36+ZfyDx7oQYbQQStOfeN5iyx9JMKjOlcak
22nCZHTSOqDG3gG7Y/Mce07RBSKyfvUdiEB5a0bSHrtD/rj9TFgSLmHJVCJ0mptfgHQY9lJSP6iH
02IWXXZ6WoG8hjTlUur2NLX0lH6ZfUGLX79w974HPLwD/Y76i86cSWYcAoFM6UPTxgRmrrArFuml
75sQg+qb5qMD7sg0avj0f+/vlPteghIWriW009aF8bWBSDLiw47GPeFsx9DqwlIBY5VEE0R4a34l
8Sifb6DvxLV9BQrLZHKwMiAznGF8jCNjN3g7ykFQie8Ku8iX/qqVi2OFNuiNt6YrMdEiSDUVZe0s
PEs6rDERe/y9tlFnBkaK0r75LfranWWGimS/ZQYGVnvr5ITpk4/hKQnxQI76YlyNlWU63zyTjO3h
nl3JpABXfu0pFAnVxgiNwGu0GuzN2A757JjytSedP/RPWVa+QLrMoCpWRh9Q6D9O+gzz/L7hjLyA
G2IIo9x6aaxrQa+uQH7FIIOo/U1nPIHt0RCXcOWAz1O069J2zgy4SRWkDDusIFaVXSv2Mobh6tYN
zOLMpa4FqnFsc1hdP5StO7HDcez604EQZ9vsnjnG8gzngko85YKteCqh/9qZe+gop6/mYg+LE+yo
JAjG4mlQwH/jpgNgv+wGrO3roJrezPlLxtHtwW7wvyt5HcnZugJs7+rYa1GE7Mu4+m2b093FdREP
Y7Xzx7PhW/XyqaIPgjlZqFzEuIo03st6kDaKVal7jSgEg1XDTzxScPJX6qvaJQyrYeOyslVHg9OV
6az3Z/GExvMmv9JCJ9fW4cZy13IZzc0oHe3fqC+wlm+WcnTpOJ8qdJXqmMIXKsGhYoyUDlCc35M+
1DTVoQC9WDrb7/M0twY3CQaIHzL2Nz1x0+IVeLygusvAZcYEA8CmKKfkSInQFzAtSjDncfkt8w8U
0sUmT24PPInT4Clz+qW2VFCwy9R6E/i/NbWKq0BblLRDZ4oDhAt5xTMuprOv0EuLcPFN2s1FklQG
jmNRpoPZ4pbQEhe12qGcdA8nS/iyzGFSa6yKJZEiB8mqjja2YWz8ptfTpYgGojxuJkoLZTDFz0LC
+udP1NMN6sLntZpvgcfmgBp3eMCnjG27eHJWuqLyZ56juSSwkqA9Hpz1c2ykB3RLdJB5+qyvogem
EugmoxHb5+eSCsI2jFPmZi7nLwMjFTSq3Je7AV/Ddyszl0dBI9X3YyzcLQk4vmyRYg1zsOf6UusQ
YbsSWGEzd31LNPW4FMUZQrzG5qHqNz8988XVxepMA6Z8NT9AKNwB4jCHev0E8KROPnYQd/2C07eG
9GSuuPS52/PDE7iiHBv43XVUUNCZsS1dKc0HytAzSiOFRmJdMsiJ+n3tAWKMcTZb+roLcmeq1bHo
eso7IyVabkWczQXcqLO1ClvGuA5nbOfFCO49vJNAcu4W2dytNQYeXHf6fhiCROYHX/CEozcV8in+
TaxbdgcCxoTnVJ7OM0WcN2yC8NS0HZG7nk8cWVsmetXJ8r5BBj+3XvYpmMUUWkwdpQABgYe70sOQ
WhUU5b748EK30w5kDdarZk+u2SHaV8gf2EswMAijn/968jANlitQ45CinXotE/n2Cg1EzEHQVSSm
GDzVhAzCrJp8caXeCiSKtt9aT97CBzrsQ15Dkmxy+yGn74S29bBwx3eWkjcn/bacHhv8yaMBRlym
Gb/QzxLcKmz4FY9rylhtZz/yaK/l/kBazmsD4GFacOouaKhgDQY51Jzga7R/jrjk2XXyNJvG5XNL
jAC2pvzhtxbw+KkIgSWKsdDR74Aq04UNB6Zg9htYoWdsrTx0o7A+c4oM/0XhzANSANzC/W79FXdw
4uKRtgRTWm6BGr/wwZMwsM6F8T35uG+sfG7W9JRkuSVK99kEqprj1beHxWlRuhcLUgW8IQ13Lw/7
U/Amaws4CoFTF3gWkphN9eMsKH54AZMWsKB8Z/O763ZWXp2ZexLfI41Xh74KMpvAVLRtXDwbBtlk
NJmOiO90oGIFfpDPLfnmjC0GwxvxxEwKzk21aC1F/6UtyPI7K8DSZBCFaL05lAbo1Pyz0cynVZaP
GinM7pXp4dS0PR80VAxwyOCxy6njhc6hu6lfEucsttCWNiyDo9aU4HXlCRuBKl/oXo9k16j6agYq
54Gh+fuYtkuYIuUciRH6NaVy4Qj2K/meo9Bp9iZ6GkMjDzSravaoanDqmNQmgjlf8cu9WGBkcGsW
pEAUKaNxSEtfx+eKFE39HrB9pP5ihM6cKXs+PkH2D0CA5P5UlMum64p7GHVGfm/27tmTKbiWEcLl
Q/ENmRw5Dfbiyqqg1RRGit8+V1NT8W6GBvjTq9FzyrnxfMbQUiNFvhdH9bLtJ7Lkozi1nY/N2UQs
E+9lWAp4nurz6UgSD+rxabIMQvgKOPFW4Dn9cSBSy8dfrUio54VK3Z3ZHz3CUTBB4U7l0BMJOcOg
oFT7XnJha5qvRFOzjE9V+/5g7Mr1F7YaKxemCCjMV0O94w2vc/60Bc1JO7XkVJc0tfSmWpe4cj8H
y2oKWAJKC5/gp7ZhmNf1/8fCh8YlO/biviUDrf7mwOs3dmk4zAMtAfuZgYCRZEpbWMI/eu1/WOJn
LZUTmtZ3AzssXloJxgh68IWG9FCwmexbnoxFU2jpxTVqULlpGGY2m/kszZMkAlxi+nhEYxQ5jVrh
v+I04Equ2hssdjdc9F0ovciA4qb9+kK6LDv99oORAmt3PerHWMsmEx1qcTK3Kqas2kBHAPu2vylL
RKqo2Vlyng2Bf4pTe0Me0rsPkffq8H1AqlblMKxaWm7Vtap6wjmdeE/uFQkoVykMiwTnV0RRJ6lk
66Dw18erhKbk3oDOW3pAgdV22tn0DsJuYs+4KJWuua58JKAmn/NtsFY9Khv/1JA8vn3w3myr+DL7
/EVSkCq/td9VDCAzZ8oBjRJs66ucdRjKzQ2OLf/A0z7uzhYlf8JjbkJHyctXSpEO2Ha/QKLdaDaG
88OiwIEkW9qGfyO6+BL14N2ISmQXn6C4lETM2iWhQ2EINTWcy24leStv+ntS+aN1R1WE0l9nGHgT
lwiS2L2cafNdbW5gsFDZeDIqM39jA2JHwaC6bgttSoVvyhbjqZXa2OjeiM9jJgnX6b7Nl//WecJH
PBIxYlCW8xyAcaizoxFeGWxQnN2rXKY+9MPWEunLIKlMtusMmuuEnVyrRE6ydnXboyKahRYc+s0v
fUHdqhibKI0wSZmVNRR11dIwUyfUN7HXaHNdRYdx+m07YTRNsoNGQp+hzuo3gJ7ZVmd+ZczpRTRw
yxjaBy25OE+2g6bJUR7kdhouKBGQUWgA/CtQQN6/uy6PcstLRhCX54s+vgB7V8XDNDVBo3UudIaJ
Ke1GhqhexJIQdpqUcmKetlki4VUL2QSiYp/RyiL4VIxWmn7KP4A9pn0dYZoPofwbOvCylRlvpM4w
hpuVBfPe22/k0WOrWo2jJBy/y6BiCj218TfJXfSIpGwMr3nt7axTbmMPhEJxyyBCNus/GxGmdF5R
7IKbPoe0ITXTlNLkLEhM0BJHfVbNMY4qbAzuwajedSygn5EFuOHFm2CehiwbDf5eLmnh20nWjqXO
7ILjzMXVdGeNiqkMYlwIGfQGP4R1PXInjxdj1e8BaHYGmW7VXdSbJyumaJ6T0nlGXju2lE2rNrSv
m/6pAAJIW7yVb1cqLMmPt7SOaF7Z8ZrrL0T9x1GlHtWkEAnQE7ykv/6ndBlONp/BFF7rQ2fmB25d
ITfkXeZV1fuZM0dZCU7cNKL8Q8jcb/Dgse1Ps0BqOZEPfESXrYbceNrstHC9SO2UKyquhsRf5C2k
R/W4vY4q6hUcAUWOueDpnd0eYBNRCO27hWuo8ayX2AvKF3Xwogj677TirXr4Iiw3VbvcHogLW+FV
ixUASzdaUAey8fyEFFL6buy5I1NfTqAA5SNC1IU0YJ1ePoWSfxvxCOANK/meZjgfJSPtQ+70mlWm
nCANrygPVmHy8/aOpDbG2LfV0X1TOOojTB2Q46d7GAIwD2kOS6uVB3+g0WELQpyhLlcNyGy1DoPL
xgGckUlA/Thq+FLatZfvso3nVzAP5TRYCVdWvk9iBiVxHRI/OSdLndYlf9R9YXbavcmmW0zJzoEj
IcqVLbO1c7ffsYgpqMGmNo+CpoqHTjMtPx1WgnY5Tevh6NLx8ehdhO9Vat94Jg7VWVx9voxB63M5
uhxEeO+QWgy08bIoumEi/oe+dc/4WQEWJm6lFjeLugig6qp187w0Vng9hd+0WcbI1tLRp4lnWR3h
I4DwWlh2V9zbyCg/Ka1doZtm8+KZyYtuc4XSZLhf9d7d9XizCODQP7Ixn7jwmt9vOPn33u/wglw9
5hMsNxB7ywsAX9mpW0WbSTBq7ynQCuAw9gXa4aN7dF5IWfMbLjhQXThEUYx7OCL6Z65a8UpFlak9
ruYCc+2gO14pYrqNYtFlcNGT4I19m5WWlQCFi+0NWHefzApPMTURXl/rH07Ca4EV6DqAds2BgVK3
YScrGSTH2iFk73f9SHZsj/P94ScE0ExkhDKRy+myetnt68l+gVpLm5YOf08UIQ76yyoqmp8OYYLf
aGbmN+mqXTL2qcQtD8En9pWSyoouqfxudrTfR1dMVwTKR8SDlia8vbPDKe88woChwUzQ2V3u8272
IcNfO9ZrkaBQ/N5HWQRZiO8Z2QFejHrR8wLLUxe/GhcqMolNPPWcbCE4XSo1NykEMMN5YrSLRjtd
Y8M4hYs/5YIWPcbM0/Cj0KaXbhtC8iBTpyYBRb6BpN748hZwNlbceanim1vzHglURrEBEbSfU+DV
psjqOj+QJMKYW7Nwn68AGhZjOtbYeSmU3AFAm6ZvJ1SkDKpxZ1pr3+JFJCRwb16vR/lv+UztynK2
DkugalqE7e1sNr8xcyPj7zbGfo4uFbBu0flmmorFhQHzv53qcPA122Wc0CpV8YPikn6CgtAWmVrW
QcX3LPBv68Y3rmbg88MkgOJdH5Kmjq9lpxgkJ+c4bbcgwHWEMvktN2NKYR0u0n3puGn+ieQWVUF9
6ON3xFuqLG+sKMIH/5oQrRAI1Q3aGhDztpLVD5dlfA57RrOgGfXPsz/skKR0m7zKGEdsTqKJ/uIX
zezNdHthbzVhEHMjNdRDP35B5PP4o1RTwJpxoe75rXeQAqbDarhy+3Df0p7LGq2PUFKPvy2QWKdC
bEJ/pBf0TPUiYjUKcg+iJvPFPQRVjPj9LIpQvIdrs5BRRAxeSbwXbD/UVE7MCa3e/P+P8duMCvR6
K/9KorwSalyARI5hCLCu31P+g0km/yMgHSiWur2zoBC6NdhvIr0gth4Viwv+7c8DvQft6dJL22Oe
9wb31yhyMAX9iDFmwzAIsZbRgp7wM0doldgcrDuOYa2G1u5Mkh3cpOSdAs//XRyCpqXuvpYLUq3r
ei6lUb6Tf78FE7trz8bJGnSxP9acWWk3gzVPCoYVcnGVxuYHkxbqb3HnB4RZ0DHwfpXpWB6YsfSB
zlHkDb7M+uod+lukbmzbXPlicb8lO/FB1KbWQDmzvsJ51hef0YRQAV9WJPsF0e5ObYibXet3jkSQ
WqAdqkRGD/XUkQ3CN2tdE7LtsN/7uYRuImkLkWS9gi74a1PNiLcbf00Qs5M5U2zm6HhlWawz/JcG
ck9+ogdk6dSBhIWZe/bAcyIqmCsPFk0AcMXsu6omFPpyDM/wg4qUQwSL0yDsWyJ498VeAojk7BlI
H5r3CXZWws5NptQ2ZgXQyDjnSGEblOdtSoAPANJzYaRo+rEPHTdP0ZbieBDCaZKP8dAT6/qjiIOM
ojLLKLaSR5ER+CplNCT4M8g8X0AcmLtA9ktZCf2fKkQXmCcYXu7ACd4sZZOW5HPikuTrh50hC3ap
n5E36RX13DnW8y8ZojzHcwgJJ/hQynbPnZZV6zb0dBAnf+pKMhSzP7By7BtEwxactOfCN70XvB5J
mOX3I6sZVb2wnRAO0lRQw2U2qnq8kwoGGOwsNsPn+R5MUf4fkj0rcyo6GV4KvEMb6ugvDKaIur9O
O3gW+FAF5V87cAGRrNn1pvqozNKNxc9DOrpVJj3s0ZgwKZKzHf0m/pVcEC9thiMDo1rGo7Y5OSac
8l7C3UdZxHet+E/R5sThlRe7b7PEJClCt+Wo4vqkm2L6IIBSL0qsmOKnVQQ8QUlffvopeqEQY+mD
IfpBTxf4OTxFbgJTakYkwsT8xW/cpFsFwFTrkMrPqBea5PLisnE6s+RsSjAZv61uc7oXofmanQJu
7q4gJYDpQjjHDnKj/+7UC/mwgJsnG5v7OtdOxc+XBK6jHALfn1HoH5MPfbwmJdm70p1SU9skb3Gc
TRlls16PQTVZfUz3eOZ8THRhnUFv3WV/5v0L+BZoLe8o4l6tydGMk7A7m3e5tFnKNGygye6OU8Qh
Hq0WqSdRwRY6sPCi9lVzHY8sKfGAMu3IIujzwy9G7kVQYOdBtzAY7Z/HNJHRkz4hC3pkpOH8TXPr
/m+LaZEPunx5M4j0neYvvUAMzepAyhacoGNKhkhE7fP56Q8h4Qy90jd97YLgDj+C5eCThzx26+Iy
5LrRPc/GkCXq7114Vugc6EdjfsZQij1WiLIfexolN9G3Z03XXLpICN7ymsjK1l4dnIG+nFp1Fbxf
ibFF11ziAqbsEzblhAGJc1c7l6BrlFRI5Ai6DWxPhjrkke8NC/RHrjnhRuUh7BEKelLvjdI8m2uN
V7Mm+GnltJqlnD/aPeYc3lMy7QfSJzGBAwrACE+HCl5bSaE7ZcKFBh+yp0eSEphti/jvdcKdLEPZ
6e9HkUl7Loonl7AzaUyssJQIE2HEYYC7q6SKGnUawfEnjOtFTyVoQcCrsQF8fS2LgeoJxIJ3BOz7
QM4mzZR+kTNmHyeXd9elDwk6LWjINyQbei+fZUkiT0cCdlOqf3qPkpWaeMQ0cnBEtr/EQaqe4uMo
3yQsSckmNUo1rxzj4dyD2chhktRs8PnwAZZQy8L/hGrGbiq6rW1kBGy045nT2awewItFRwRnhYmb
eR+sF6iEYI6EfHGpCxVOrFilbyNvXJGsId3aOCJdcRyFsyaUr3C7+QdMzgSQAbrzxyns7+eb9Fw4
jjF9tNJDjBWAe3FbYg6Sh2tOQMhdsS+olULnB8q31xvVN8WbZ5lpRaQx0heAk7iS2w0onVwAdrG4
tapwPPLEieN9hHDx4RiOm4m51And30bcrEN7j8EmkIrxZOnrdpge+N9hToTI/7NhFrRz2MtfK2l5
OZKGhxrmVGnQIlu32C/cJTXQBVRw2u/92oRQzX8A4alpV/t/sUztScjUeq+V9xF3njYF2CxW/Ihu
ulgR0/mtSTw/FX5OWltcKb5DfvWPjoS3hFO5aVSIYwoDHJ2lOoObEe8uIkWVsrkBf8RRgeZ1cJLo
wdzVwxAA6o/07fJ4YE9lNfORbHX8jcFDBWTIbGKi2iJwyGjfu4KOSUNFEnKOVKyD5hYIC+aRp0R9
gWAR93VNG2dqNDQn4iGIjuFjNKlaxoceNQgi376wYSYeT/USJIGT1hcpyFlhgAIxNkwNqGStkymE
4KcXgabcFuOFamQziSCnlyNLmMEZYmvXsTgjhlk0lmg8dtMRK0A/WujEBBtJLapuSpFHf8iAXF1V
Dch9eUaTbjO6eqtInS9Gu+jnXPPP+aW7bG9aAK477j+Q7Kie5mY4yiXV9/TbyMRAsEkDp8tqFfXX
lpQWEs63wdeaHl2HZrx3Ug5FqrKOfZ+b2dyLnA9caipUO0HYfSeUhuSeqw8+EAZn6kJYlrW1DqlB
W6TIzxX5Hp2zz71G08y8PTxaXxhtRAmvcdVIke5fENG7iB1Gy+7x4Eyf10dSZdbFuDoD99hbT5H7
54S5uw3ZnvfFYRdv3ZFSXGHPrWHLVh7Fhlfj3NeFXnsN2fFYv+RjOBmyEIRLIyABPGNdKRCCtzkB
qIvM27r6OlhYh2aDJNdr/ofxtJsmyjg3hr3MYRKmSgLlpcY4kGDrC57uKQ/ETjf59hRrfCnVwxnP
/iQ8VZg1NkXbP30Z7fslylafV12TE8Lu+9cxbU15SzJ+Bx42cIGnmmIuXPbG8GaL//x29ILLvuLE
UT/8l+1Lkc/aWtuk5pAAQx+mkQHnxBHX7Yd7kRKaSWgB8l7PZrSHeIL7DCrWm4iT9dnfTkvBXXmC
ffi2rHVTqOVP0mAytHlFnAdYwIzVOSzd9ifqAqhdTiZRJvgwM3DMQaH6oi9eLmBBQO6j7D0R9h/q
Qy/ibFGK9j7gNwPkyoqAytMXmBsjntGK4M/Og2LNvrA+DsUz2STZ/Im33WLYQmG6B0AXz6eLE6oY
BbAxCH2mALEo0j8+AciWw8KTA778ILHdcQbrLz3QRW5M1z4c8y+fmVAmupD6XXxhzhgurEzW3mmo
JqWsa20Kz9nBpoqTLpIlMbODkvhW5EUCpIOf0Zn075J2QWJwWZpnx6yLRYNHK03VTqFg2Wd5Sqss
WQ+s/iMfM7cmkmN5mEvKDPIT48giT+YGsG2/b8uogDhaulJgvYXqkWl93V7WPY6jxf+4cKtqv2Ro
GP7koz2peqHR8sqSDr7MD9DqufntscxARhnDCAlzxEEqUcqcyjY91goLGjGFtFgbQp/jgkBHp/hz
VbzlspcJInxH0SBGNxUUKfY3CMCFOAjwAQRI5QuyRNn9I8/uUj4Vzms043iA9iTpEXG5MB4GCvxQ
2yijD0EG9odVrsyCdg21JhKGcaNgbeb2lj/8c/E8F94fb/5QVTdBvK6ewAgxxCNd5WyXvuJkHWY+
z/apnioZzdhQZmMtSNkzpk5qoARmO0TEARICEMydolBBZEHN1tKS1Pda4NNx9NGQDCDVDF7hrsQb
AuFWQjv17ChyT+J4x8R/4MNwmV5aw0ONs/ufq6gMRx1ycyk1goYZfccdSYaSYeKSYA9czwTychgT
3F9TrBfhL8YD/21t3WRlWE6FViK2wgXpRo0uz+rE/RlQaeK9mqYoJaavGnGQksvLt4d15sy8IiBx
oY8nTN/NrkZ+0EKDkwu0RASF5S7/GAV5nzH1oEn//cjI9y7n00qR6aE6Fz/CJ7jJEy+lDPlNAo64
qPf2IogU492YUXmIkQXgS/ZD4BBXUS5V+DjE8EFAvJUsWLAYazXXxjtJ7Cca5do6IAkdPzrMiFel
iA4hBwUt9J41rcPKuOzS9KHlNmnA2jA99vPLyQ7nPh/vDOfYgKL9YPLBHBgnU6Gz2jw1uNHSnFqz
G3xI2OD00HMTB9+iXy3E8f/9EkQkFYN1FlW5k6dsjm8K9Rmh+5IyuqVgXB4zYQvgk8B+dQFtm450
KdgNTiBjDm++hRiWbGC8teh6ZO4b4RmXS6HIUoy3S/iq5vK2fJAdhCK8Nxgo4QG7wbJHOpcIPxmF
KyCn4R26rVNW1lqs4JxZT5KuHQL4jdiWXG+uA/FhbeI2z0c92T46bLlByXhZSlE5ob5GXF4Zf9Fx
+fPeJ0AyE1HW/q0c5OYIm4U+MHBqwmJSSO9TIkKXityGch+pYU8uvfsJbMCm0PfPknA+/6ZpGGD1
79MANetDIa6HXEBAr4RiNOSy1Bnm+A2vn7BO0Z/l7eGxdC8V91KbodDVWu71Zfc+khCfcxjh4QWn
TKgleHBDd1CKGOiJDiZWeRPEyVj9HsXU5TnwZnd0Wout6ihzWNYJolSvUoMjOubi9niu10U0Ms9Q
SvIfki8t78ef+hvNe5c5vW55/TSj2oqc9wtS8Ta/JFrgmnGm2yAa52f51tjVd6wzh6hJEHm+LWjn
egfqHKu+cE0oKTOMbRsoPoDnT92t/MAbw/jqK+crYL/IbUNBJ/8230fMZDYczB8hFqP/WLnl2O/I
8kvBnbFtBuHXApPOjQR0NNq2JUGq1Wa4gKUjbY1o1LSpkYoHYRMrmQqjIsHKFtgJsfQ5Z7JoAOkH
VXyKZ1RA0x1U78MSmroDgKT4V3DY6sYaXXSIQPwCXcvHnbYAfqJR8nwCr6WVK1/FKnQY8PRFHPiu
Z08sm/AiQZ24j/16HUscGQhTCUl9jkaPdVdGdQhUd+zhpl1AAFzKe0c61BHWcTA0GQygHyR/+2K9
XmNCCNb675iTSx8xDhzANnWnd3LHMNuzvAZLwvhFb7zDHNHOJ/VWMOC2nNDqm9c7O7q6KWYtOZwd
fy/yfX8MwRV0vtx87AoSgypGBkfsqXjSz97XGiY2yGQt6WD3ZtBcjQGmcHDrnsNN0dagN46zKxxl
mkXMOdpIjNQq3gd9ruZdP4nNqoUClTg/yUAytuRbPP3bST/fbgbkmfERNnreBCXVVXy5MNbarkf6
AmE+YkFpF27ObLQTL3lm8U5Dy5ZVb8xCAeIlJ7ZKNfyw4NnJVZHq6Zo3OkZapmLgmS39oGEdvi09
0DkMF2EZgT6fj6g1jt5lOqx6dsiiPdfC7UBOSKSWkwyrXSB+Im7oGK+5zShw4/5iKUNFk+GPNyuO
G32o5H8NpDmwgAo3a6ig4AVj1ha6J/ORqtLW3bgz36drsjcq5yjJX0dO9fNCZwYg38krXtdU2noy
iubXEEJ1R1a8weByiEOR6Xopjg3ADL0bKwOwsas1eLVYHJYAWepmHl4PTyb1djUXB3/U5LzoKaUJ
BHyR/jrwcLvrr6jzjj0Xj1bcGg3VHBPW9PHpr/GLdiTR3kTOML6zWaO9Hr0Jqoak8w1yNBRviuWt
qeZxKbqekH0LAyj0mPwz34SwsPJp/xxAB1JCYfrfuh6x2tHpB7DmhbKQZZRZPlvEdgZLYHa7/CRm
Y2TVJBY7kZELKmcA6HLLZMQONtwJN6sTWQkouWQ9ndEJSJ735LxsZYO3V6ZjOITxNvjOs3M5yySz
wY89FQ8Cka4eIyxLjZbvlJIJ3yaEdNs318O9fjCkb+0wPPBE76ugjGexRClRNKvUonv6D2BP0azp
k8pCc9/JWydcVFnXASDbh5cGH90VoIbgXSPZUl/zjy7U6XQeHkEp5rBM71NG7soaG08HLxuXhjd2
LWKB1fD1p2nDn6PhMuOUK7ULR47370iea61kEMmdmyLiUgo0Wyp8H7enUvc3eep9XQHG0IfrHkzy
VmyysOw87JKBiLb1Oqz0/N52Wf9Fz6rL51LC07B1iv//C5vkBK5sEV+8a26yJI8qSuFxHpC9BvX7
PGobYgrH/ytBUg4JXyVU55Z0a1ORnlr5MzAImKl0Ec2y/Zi7xCWM9lIwiwaeyHg+ZFQGAegcJXtX
F+XisnCkFrPtwF5AzjaMpJtty/1v1Z1WfZohfCA/2HOkK0t6a1MO92cy8gxk09aRMJxBYAkVquae
8gNTXDt9TPPJBMW6WvFrIV4bBELM6eLLaicuc31xp6f1E49g/owDGEjyUwXyeMQ/Qz91Y3ZiV5fU
OBLUcwGYCEsflJRSy4qHukW1hYheTMmN4YLsEzFKxzGp7hWpu444XIsKCAIti0cZjhnNi0+96lI2
UhVsBC++3J3gikB4dNS9Ngek8bgT3i4p96VZNmMoTQfbC6mmJFmD30Kp28RycofjWGBN0pmz8Se1
rUMRsKL70JLMbqtM1nyrUqB/H/7FSWe+Al6WGH5Xz9oEYK6481UoFzpXxHf+xh8QMxBHbt8ygE4J
aRSvMa6BclQxswmy5wrZecWV4Y/cjKTwBZQxQvN+L0Gl/Vhq4o6iT4OyNHJg5DSdpN0aBEMrr23F
8F8CehRFz27ufAffwAI7MOflBgfK2/bbEo7BJ8dNIDqQD1ERaupvTeLKsB+fmG0ocOien2ngysBC
OYG//fwiosmp0R8U66Z6o0prLe6TrnNjvdm6tZTNAO3sT/RrV3iomSjqjAp0fxKnzH5bCq3X04U1
qH6ECUz2zibjtWFlVhAe3qO0wn03iCv9wnTdiWh/+W8BcRBIXLj6Tb1Nrc910RztQH6M4NV3an3J
O5K0DsbXrisEdAz8xnwTMtINv4CNA4tGdI9Qi0Oo32hpIXR/ILPyX+slzYZUo1fzULF9zhWZdKjp
eeFIR/aofB0XUkoqCxiSPKoFwhzmpOt4hMnlVKn/33E+pEk1QGAZ/Jg+7ZPKKaRWzsLSMHYuoiE+
YqwXpFoQkADDF32rHel7bS/bPbAIuyc/Bdc/644gCCaE01jSCkH0yDNnFA2+UVnpoT4jlVkHX735
NHS7Moc8GL+7B5BR+Czd+h7XqxSMt/EkXId/gWcpy5ZfAvPMHAY9tBBPgnYnXG4BtQd3qtAm7fOh
Vm01V5KGSrwRjFYIvHF5D+QTDP1unGjtG1jswdQRHvtZMwTlYZ+AkMc2Hm72QM3eMRjd0X9QV+Bt
/ddTMhTw9DDWBtXnSgFlzbCx6UdWAJpVDuK8rKwS9OiUS1g2U1jQ08/tTp0dLMglnVdcfPjGLvpb
eQqAyBm4FMtCGvKb3puw3aYi1xmBu0R68z9bWHR70F1sRH7ZJNw+Vt2+asLGLcdO/WbuD4CX4T+A
bhX2aEUWUVmR9N18MFPA4iHOupuVCAMycD8BcHCKkkhTVhU55pdnlUHM6L1YOFyTFnNrv99oEE4p
BnfzcWF2Rgqvqp8p9CzHhnVHX4Pab3/5pzfLDH9Zg0irZqWQPF7tJYq/b+HDCXIydK0zKdvlr9hr
GtH4sfqz+oGFUF8HU4+2L0QQU19br7WExD38IccCFy3xkgpEIxO6LQwdbQwtKJtZ+0gm761395Br
g6CD9J9Xc/OtAkKmO29EM5OHLyRR02OzXllovYtoDR/INiMxaL4rWZzv0j/lVCCMzUQSwAvzymNg
imsROEo0VfztmiewkScnuPpBUMVt0qRHegI7dm4q/V0BN6wk7hqsB7PCogqDfnVan33MODxwWjPH
otNNlM3kHetClD6PFABs4NBrRlowAx9RZObrKeusEZc8CBaKjqoebcKWeVGZCenqVk/aS27z866u
ZgajNFLhGMR03XBUQXA71AZiWx7HMprqhrr/GSzVvEZ6DSS8ryk779kV76wzaWQRBW3ucpVp5x90
CvB6abUSCZe00FxZHkVUur3YzsAu8l/G51uU7jJzVnjBhiIPxmT4ndE2dDYhiVejUkFGsy7lxlf5
Oftke6QEoFzDTT4abya5N5/CzBcoUt30BrKJcPxzcoD2ZoR2w3ZUw3S5F9N4dSxQm5r6DzX6lZU+
8E9RJyUVOnQTLdhhKD0CHLE6514ADwlbXSucRHmn9IFbCfz8E+JPaMeO+oOVXUAOa6vNO4UsoCwk
S5OcTVhgfhLOCX14s4pQ42U/mvVPhsfViCIlXGXSLGcAW9STbYZI8mVT7Xrd2n+H9BTcO5yFuNpk
nNQJ7QVehaaVt8VpYqQhOH7Ju4hCG1QPd1yQG5vlhSPxoCC8627Utiz7m7u/WtuTJnKxO+OyRqd1
VHi7SNdMV5mQyuhWTzox+CKKdSDkXh440vj9+5k0dA8bV3xRq4ro5nXn1UckGG/LyfszxaZHqkRj
/x14fS9ObVGkncfG5nCuPD9IntHS2qHL2VniHZR4U+kcGBbNplG6KeUU3UFRGTGC1WZAfMdtawcS
Bpvdakt8gj7OC+4TKMDABZNi1rE13ILJU7Sfmd4pcB3dp+oMf5UfmC6VrUqsWzVqU4Zt2MuC0wB3
WSAXBr3xEY0IG36XLnsBbUuH0qDvy07oaSGt7ZltznYhxjWMJ2s6rGNNpzeFBzc2MqBqhmDCKtwx
wJXIT7ebgjVSJxeBqZpvpOQ7fhuO75AM8vSXxEDbopkYgYL0qCApvBc1lO1y6XltR96Z1D0uASPy
F3pAhzToza/J7jvbNnJs8FOxJKg6sZdK7yLWuiOMSIha5dVi8gY66cIlDGb4qIg63d8BblYSbdWx
wD6qZIXRUSiJrRh6nrsuaTvCfLK3YjkccLdftIaWvOARdqIuLM11i3TdP+HpYBL0fBTQQfBMQ/+/
snxz1y1j6WjXZZkB+GPknKIt/yGarRNiqG5I9eEcLGf5zKsNf3X2Z/d/lzhEB5TsGAelJ8Nalcew
O9wsgxg1msIBTNCjMeyFkNOqh8MZZrLyt/BsYuVLODNc4PI/aoZKnQRhxOGUKttkQfrqsEJZHdAI
iiY6S6U2n16POO1mIzpi4hoPg978CO13oYgmSY+GMq0/3waMiXkw66cr+TzIqIZW2O21+5+ZxzHs
S14H2bHDt5TS9qeUnHCIMMbBcyqhQu7ruith5CpuKCSfEtNPveWSSxYr/60nD7CksGYvIsWyOugR
gcOvB2ULWHsKHpiXNboGNVqFOf5epfWnknRZaxqLX+j8J+9thghDqDSeLEd7FxCUAWFyRrLoT2SB
Vuv3G/gWN0CjaVsC1Ehi5jJ7BjH0RY8geuiukkVjRHiwnwRqlYFU9uE0Lu4rdHc5ge+dsVwUA7HT
0RKp2GWkvCmd732b8WoR7Ot6n9BcRhJJmCxK2sgGKM+mfi3Cnpnbx2tCeB45hzXnrllt66YZ4/N1
NK5JuSvUOtkFbAc5ot0oFrF1RDg3WNVg/bESqegYQLsfOScDe/Z+pLrBxMLic08X68YWCyV3jgNw
4c9CKj1d0msdnVnL+31fmYh02i2FU9R97J+SB/8ZGCf0A69FxFzu8NGcHTvvEVZhJ504RmHUYFlb
LN+i1SHZdghX8mPgBbbhWj0HzT4sW1D4K6rU6qZSEat9VhZtIjK+GnLEZTwP49U/J6A9XsxeBNFq
6xYlv2YNnwxcfrnVyJFIj1dds0mh0lRAPXKEiXdxhQqNYtLbYHbSmHoplyDmKay0AZG7htY7PXeX
JlLNZdkwGumP+ayRUE64Mv9zTMoj1jt+TcblB1V5B/ugPYFksvMciVqpDjp1NSNPuB/ItNLrDA9o
Qj4jiz/xTXG2VCslgWa/cEYzD0Qs0M03bGr1rZADh8O2vsWGTXDxEGdL/j9ZUFbMcHjYhyHoqZLJ
sEyNvAJcL/LvO85AaGmpmALDUoK3nqIqX7mvOCp54UwSQbq9HyKd7173oShyvRMy4AIWfM+H6PhO
nGsC/hJYC3Jp0/CNqoVz5m9nRdnGVf/PQmLfIQShenDXFe34WJlgcg3EinfZBd3QxbmcK5VqBxo0
WYKZdGwVY2FenjoBrqnRasxY9lvKceoyg5fa8ccoffFjyei3tGTLNC/7DwI1BKf2QldGIFOticxK
ImDk3N9pOgfyMY7RM8d2xDAmzBKBtUw6+J8VzvRR+D37poWKgQMUfH9QVJ+/jnJjh+6HUB1x5FVk
UPptQEddu5X3ZdWdkP6SIeRHlwTlS+b1oQO2ze9HG7qx46IHXgSoxK1FuppWMX0WlWV4w8hRVurd
8NTydgdcrHHGW4SLzBUjfzvBnx+qUGVtlSvfl7KoPXjLqnPDvKD2ahwt4exGP5ZcGsPVOAdW0FqT
b+3euQmTY2JDGh5j1ohfs9ogFVjO5bKmGtSwTkTylxCg8VBD+c49ZMVhANHkLpLjvA6tktbvI65y
0SVT9QQM4Q98Z2XI34nCX1x8q+Yxm28Q17jIr7jXVOKqdS+kQmxYLAbbsu/hbGi3s9XVxkd7hINt
a/lsWpYE9qxjdzcPKPNbMSaQuFUEvx1syTGdEqTm79EtTKwOeHZtqfW5xlcT8wTNsSZlnAklayn9
uca3jB0YhZhtQEMfk1yZdm/xtMlqQhHZ/UgGWj4VIvdIsQbMSfhLzX54kTIQI3aORiCEV0zau13g
RsdT5L9aEVMLf8kANCvLulYNc0MpD9r9VMWkScqB+mDrkZU8i3BX9zVS6WjIl/RcOtxPpRZoNqLD
/0yfrZ2P5DtyxFS6f5QLELcPyJhBxWwERQhLrz8V+whzvvZ/PCZcv7pde592CqNw2x0Fc01LUykF
Ny1iP6PZ65tDV5861YS7YgJNXq3+tI/Z6th5EVGUymOHnanUDbtjTxkzu7BGDB9smUu+R/ptaq6X
7Azw8my4a0dBkSawuIorQFNdo+nrUaibTGEy6XsD8M8/jPqN2hnfRLCmLXRLMyoI2AuZK95ZzRAG
2DTZlLYmHpTBNdSSwbk6bzSDQ5bJ1JPR3/TvJyBqQ+Q2VP1ahshKlqhp6dFB3KNnLG2ZXnpiUCJu
t4WqPmHFmaacx0RVBkP9LSGnZ+Pk+SvXE5qjXcZ7Zv5uQF0W+pFYBBj38Xi7yVsDJMJtW6Cab8PB
3ITL0SrNkvkkbIy3huyT7/NCabYFFlrrah3uj9NwZIgkr+StNDf+DvhFj/CWla+V/ThwxksSQ6Pc
jVQepOKQlXY5tYecl+5SWJFmI/6FQDWuOOFc0FUNpbL/gok9+Hp3VjOgd1VfktXRPBYelLf97zNc
LhB1cX1bkFlAw9ocUfZYj4kBZUTp6I3vD6nEoKnPWwFXUlUF0h9pWMGW8FuzDx7QQzoOexKAien9
ar41Wqdo2pvw0tvukspVLEvtnjO/HD8jZIgMX+yq3uMHjmJmRLdtlF42qgYH//6H1d5z9E7CrHQA
cbxncYycyCI94qIO+EpRUaBkV/9TxSLMvHEje0WpqARIrXY+UlPSS8Eb3pZ86WxnPn6Wjb2vikeI
2A9Zfe3N7vAl4gfqFw3YzroRO3EprW8atzgXKB7+I3rksROLUUUm/rwm1rv9w9jTdY7ntZ3Uyr0H
wdP1X2OhEsV3HfLakBr/wrFuYA4vFC4JLfB3xmvGhzxDS4qaYhcGNEM4OpXJPhGHsNf5xtXBc3d7
SiMH1VNYzQ/Bme/LXLujYyoCyTg0Nylp261ZMxUxkl0472cuB45SmYhosBkqujk7Nxqoly1gpDk3
gNEfVTY4HkuDzDxpjuGXRkvSPvcwrJUpJjPjbVUjZ8XncwcMs+Ydj1VXMgSNznYoB1gX4Al/ODKh
F6tdwiTB73P5aisC3R64cvgm8WytJgvSWrPXU4Qt5tKRdkhRPsU/dYjM+Wi/7J1dbeDuQEUSpYW0
kJuphD7T5j/zR0EIUove6AQ13pCSXS1FN3iCx2h7G7/X5x9Kfd1DjYJbFl5IFuLrqfFTHjC9wpD7
fGnAaT7PgstkG8iEJrWvgdDyK1+EbaoF9WHXCrfy6zHc5IZ4zm4PM4+TwDfhP7TVeD9H+Z9A4oVn
FCQg05Z6WRwnCfnLX/5K99Pi4H32uYixnoi7aISW6v2fhoRjZmdDU4RHSVD5dhscvEyyDE4qrxGO
0TtIn8EPm/b4RpcvKjNjAtp4mj/1FrTrVezW8gtdCal/LcacayWI80whM7dq/MrPszll+u84fEMD
4CueVdN1saaTVw9lYtQHQfREVOXMxJcW/9IUSXjS8ZET+YxB0WjZYjMsrzQ+trTYyvCp8eh16ix3
75AUhmcQEUf54Ep8E5yXR7thVfWMb3sil2quXwjf9ykvUY8WaS6EuhHzJr/+cpmk9Q84vp/b+qcB
1ibc+9KAjbanLHwY9VySZ2n11yevCgBmj3SoPQ/cZ07iyHxBnbVS59/jtCaTETzcfOhoISN1pga3
44vl52rCUJL1PxOtimSCZiGWcWuBQ64edgsNlV9S+X3SuMCkJ6539ZbO34DgBg0evJXxqtiXMmU4
FVIIIb/fo/MzW/WPwIKPCNgcADbwLIBSM694U1kbXYlnRpkNvY1i79wsp5G1rrpAtQsf/u2TI9Qd
PMyLrHje6g188EsJy4a0gnwdOEWeDYz8lrRiLPhkFtYBOGbpEwx27XbmW7BNNW08mJQxp7Wj370d
EKtsEKSvPn4E+9Dnd9SbtFksrWLwmRoZYvDD3naP7IJ6cCVZec1ar6AtOPrik7r/iF92XoLVr3iL
g8vkJOU2NXOdmYCTqtBcMktUhigscMd9SxrVzUeG7ZAzufi/XSUbYZ/OZ2C8cbsI8/KAe9uF63LH
xOn1XU69PL76NauYi186pjOlq9DUJOhqC/VqsN91wZPb9tPcEOty5cMWHAxsX0GFmo4jNUY7n20R
amE1Muxm1v02Kb+/yl9urdQk/XVJHrlphd443sQFTdy/UJGYNzkT+BuTgoxrm3xE8od5etvzy0KX
CU91bO9NxNK1iDf/oM26YfCEu755ulbnmqP67SWfiFPme2q6N2f0+jqNj2Xnn+eMEBjG+gAc6F/g
03uqcb/CXOW7F2sO3wzMgjNruYAMJxhNy1fsoi1FImZyUF3J64Rfa3j7RkunFtPuQmNJHB71WboA
UlrySrBLaboL3kOYfHMnaSqpW3dVZvs359opsvqxbUAfp+c1sE+RSOxGaD5NPTdqNwjCElLoqb8Q
0nBSv+AlqCMxKlBUCnnHUgKiZpYY6K0wegojGQilWwseDAnMEDvuyi6Qkek98gXJ07doHSGdD3Pp
Z2WgDme8vlaqGoXPe7Lp5rt4YecGL67mJBvrMB64iaj2L2BGomiisU0PGtDtZXfzVo01351l7tZ8
zxWbrfbHvOggi/c6vUNt7sQ3ZKiDX3u4EisjxaQKhfkEVz3R6kUxq/Z7dBUfle8xF5uvkt8T5tpz
LCOYoqQLdhFe8G5Aysju5WgZXQc/IyJ/xjw4VVA/LlaIq1l7sk74TRHN89cCBE1qZxv+zY5mLhhP
3XXzgfdiOVgXBkVlGPSELjIO6/ifYQ2yS1oS8/LPgh2UpxSMaKCSANFLuNl8n1VeVmafdDJ5Et63
RyWNXARHYa48Jgi/IrfM85rk4LUAB2TeHIbcuVeJZkAIp33haI7xzYvS4j0X7+0vuvdjasasZqzV
QZEFtekNoh/4rGK2ofYW+iHIuMWm8n4NlLhT6HwJm1/i5BAeb1kJQwZVgClAXLaZ6XoYxn1kswIL
5kLyb6o/8sU8drqHKxNyFzsX/pNQkjkg0HORQPEhO9WtRkOPR2SAHxMwHZo4WFuSSWh3KjauGiZg
c0aJqKex6Y/0kQ6bz3dQ16dY5rix4f5/6cDKGHFPJPgO4FnnkdXLRM49cPomEVhK4aK1lKASDURp
XFVwaDcXV9xiRSckz+EPNGIbzadvvZLAyaLQNHn/9uquS2AgX/OXJVl9o50flmxYu8QrTUaaf3vg
4yJ1iz7Rqgmo37CC6+MGtNvHzUALJPw+bXLJ3oC7MrkSGeKPL9Fso6K+15X29Ye1TJ8NFwVD6E8/
0s+py8i6DHfBguzPO12NAjOob+keW0vPsvCt1GjxnZFzz/hWlXKsoY4xBkZNdJEDEnVBLpzWfjDj
FXr4OgNkTLe83lKdfMLFAZCjJWtJGHLZTOpCj66dKHhh0b5QvsYXrlHn5KbmD0Dte3TxdQ/ZoEDQ
yrrTqwlij8yHKra/8Eu9G+dqY0Tsgu+SoyMrO3X7JVL6tK9xrxP+5lFdxxyc97L7g1OUuUmDzT5d
1cMzoPmq0QoO3CDKoPb76SiuPQEvoK1yIZ6ktmApJj46OCx2EvX+zWD5s+ZL6rmbW+0sW/WVr7wa
5fGTuySgpmWV/DVpMZ3/+wbijdsTi4rr6Eaj2YCkcCE+o7/e1Hv3lRw18fLxfyCTTPvKzpdrA4Sr
0WVqQ+B9KxfRq62eC7OWlV1SJXueapPyNT1Ap268D03oX6pwzKnBcHAhNph5aKYv9dKGQ4Kd/nOM
ioDcx9hxKuRVTivID4bL5mf2xLvWjtd2tX9MxZ/ZwmTa+hboWzzhhOJMwULLkJVeUY+9U8G064D9
KvXNUViLU6LPe7jNpKaNXhtGsNcwo4R8LA7fLrRpV1eGniB8Bfdje4Zqj0AVIkpCaC4PI8peNX4S
LGBxnVy+GQRGhHq3Denr0XTdQ6DirVQHOLen3hEGUunuf8lRw6iTFxvPB3NohSbr7dwB6g/9201a
3WxUntZctZWGveFn4KyeIW4eb3Yz27Y8d1V1y0ItmNmG0FQpQWiZp7v+i6vREhbjnpgkKM6AzdLV
FrrLS63YNcZG/l6bck/U3sTkhYfL3s1HBJgUXqJlo+b5AL3BU32an69bDQXpRWxGXziSAx7jqKF1
pmUgUk+X+u0Y1AARqHFC2sh7m7h/S2OMZWorCqO3/NtdAfyCLjuSvH5vVcf2Oo6h3DJK3mhpG9rs
VoEgS5j6mnOO+4g3Kdvk0T/435B8BAKLGVF5CDogC3tbgkFxsskjDVtYfLcj22CwboqjVwtFjhyV
cXl6Dz1agXIKdG1BjVybo2j9cWDgjfyCVw0oqXx14yYmMMRTc51tRmbNC6jrrPzQLIX8gKBLDqSB
Yag9DoBJcRozt3xam6AbQqrODe+nU6CjMGgCqYircEZiEPHEx7ibEEo7CfE57rL4zwuBWry5KKje
qfdS1miI1j6uFJDbZzbuRj28ZJFHPLqe5wqaG2WdIR7qUNEY5K477B/YFpXPGFoqt3y6GDGeBVkJ
wcoWrDy67ep5QavKur+uFpUglUm0ldsjFDbwvlcdLclBOSRbGQ+0gjierQjMaoNKdNsYyoRMyE7A
lLVTsSKJqaTD+33IjwgFenI37T9O4WMi0UVZdYSgc2QZKQbMEQeMgrT8H3cIX+3P4inRK2qUC40R
kX+k9fMWq0hCuPUiNTo9A9d2+W14wRVyEJKPcsiUHH2+rC1FJx58BHlBToY7kbSQTLlPAySeBqw4
bdSFifDE/Lx2CCsOEqYFF99i7yvwor8lJN/2c/KRrHCREucfShibJyo/FsPC/3lszNSrAhDDRZBB
zDNMIFDqL4PvXpQq84kFHUFDBV89rfJ6A1J0ECSC5FbJ6jFBV69ekN9EtbAzN9mPUy3AbR6eyzk7
H/vJMcfo2nzFLQjfNuBXVSF0r0XcGK1cKELCOtIgnmKFsk6Tv8uLrco6L72RYtcepcqZNEnBazDV
j/hQ4jBIGnSK+jyIFbVlnLahS6xtyfPl/d/8OwKblLzU6HUPeC6VM+NlqkD8FNSQbAhMAmO5XjTQ
Ojw1U676BGn/aSwscFbwQMeLQJYQniPw2wQSReO3XlH7OoIzUE9seRd2ykNVRObiNqw7V7Oz5Adu
6Q2dhxF8yvkDaBBuehqFNHKif4JHMvBR7urDrt17CvIoqz+8CmOiShQMWoEA+C4Jhx2lwuxY++Bj
zNhWSNTchZdpEKNKiHiXql+3UXX+ao+LLewHFnzIq7iO7J1Z65ZhHNqaYQ9oDz7pBLPYvN856D74
D+Y7NR15Iqiln7aKeaUtD+JdLYAVFeUFA6a386wMMumtCWM+Ogowzi0I1vbb0gMY1c90ye2M9viK
GN1tcu/0JMcnjAbl8TOWUz6tJ4NUe7fSJ4vV/xHyxmB3ujnaIHWVzEcQqqJPJbyLFBw/nqQeCYNg
k0b4tgq5NMHrbpdf8FDQ2qE5y9hnsykbIDK7lWu8NMdqMG5E1U1i8SlmQxhZi4UGE2ae3Y8T9aaQ
TSGTc6DYzxpKkaeWBpYWmvXv03pABPlyTmaDXV+97BqnG3BOXhnO+ICb0b8nDqUELbiP4O66hACY
doON3Uxxbu9o7N7msMckJM49z2ut2ZhVPAA1dLHOx/LSAbW0C2nVDSxg389SgaoZzG1NaLGWX8gT
bhDvP6+JwP97G7E6PVBXr3LXOYsbDIRPIUeeGbp7iuRCa9LmNmX/b6Uzif4g5Q8IfggyIKBOWmMf
pSJOcNSmbsCsnUZQSnb1iOwR88VraFY2+LrLbrdljxurNxazWg5AhLSS31U9TdfZ3jIzt+jNBT9k
MumAyef7j6eb6bTU8tMp7G8Ei2OtW7WuR7e+PnRLkKUbdjCKsvKycoJSHSQ1+wyj2DJKkQAHzbdW
RRw+LRjugYtsfTjEyVTrfGz/qqG+zym6K7FE5eWDo44e+zwlZxx9Oo/8pXgOOyCJ6351q5yYqY8R
vuRz/bwttxn5UeA02MctvH3GMHfLIZKeaIPX0gFJJj7XIsKJlkaRDGMkCylz3fqBAzk81gTQAVBd
BjwEi1u9j5pDGWn3wrRImHNFg0MO+cWz3XIntRMMEAFiRul1tRDOglLwkWmxmp+OrcsXvzB23sb6
BKmwdq2msrdEwfr1BbYZxmwN5v5IEKjGW7xX1lvvabA9urtM9ItaqTu2DVcJ5x8COWnCeOFS22Oz
LGtwIdlV0Do9lJO370zD+XXJC1wvd7Ru3vOG+x9zlOnOOIWYbk5lNDjdQEjA7+pirwBjJ/PejpZT
RTkNbA/AMpEV5JI6B0dFUUBLDivhnOtVRYiwJQBgan+TxIbQyBcAPVuYyLWLtDhFNlf9p99BFVIO
mVxlNzrdjy9w2JA2xXRPAmXeVChNmNfVoDfK9IKtSpjj5C6AGUHT2aBB+YqMKY2f+rVAXR8cIAen
Dv71cePu16y3dmY+V40/OvgTHHkRc4SCLRwlsHh0BF52tvJNAitT9qAkZH3d17fglbpxg/DH2Tda
37si528mh6VpMGVZ58uwLU05y5UjcD8iCBdXQy2TV1Ci3dObnfEWA3M5apZ0YyeOsQUoNukwAtKg
Q5QJ54RRmOvF9hyer4ytT3gYvO4okayYYCvyl2FCZJ8dMfbHFuv0DoV4Y2hJMxpKMLyA3fJHorNs
iXK76JM4BReIwRx2dA6LLOwC6c13+PBH2vE7f2NlERmFaSBk2977Zamj4IhQmgP8+XpaX3iUV+xB
lW7CQJb04KGOwgHM0C4jo0WtLhJ9DqeaFEeQ2FG5dJN4N3o/2XT4CQOujtY5aZVGNlJzobhbmPlc
YpLYzxnrbAbu76SSNahNX4smJIOkvKb2maQ40RrGHDyzYOFv1wJk27WVuBwHPeEfuGsT1nCURlc0
f60xYnKZHqfSCxO/PmInuEuywtVn499J1KaJdmP7KLUXnDq1hxwvK9HmTi0jILYdx5Z2Kn08cavk
mYKAaRZ4TWzJMKezxZQo684T1yTtXncbLUasYBdbOryezH00YcG0m+J85LMJZ6CTphfw/QfUCrA9
ZV7zOuXoZZklbMUJE3NAr7FB+mQ/FSfSFyVWj5R29CeVJkNRjiPwt/x9pFtaTWhwE8ZStFIXJ65j
Lh9m1iB5ylVn9qCKLAxYDMjp++d/rEGKRwO+Gg1uBoHcnHm2x1EY3etzZbakXQ01HGFoOavWeeVr
ySXYqeWLRd33MCityAfS+NwpQosEf5HxrVR2XVHBXOBzQ0QRGVnt8S3/nYG3lB8zI1D0QDE=
`protect end_protected

