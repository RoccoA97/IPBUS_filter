

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
YWwSN+9l5ahBqN8tuQHA+pe+2Q7Fh9//dR3H5K2w3KRc2pla5S5ifvTi8Ak4V+dzPFwrZE+Uv4ZM
WqK4mWAaDw==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WcjiphsvP4YifX33L+r4vrauIXRkGno8B+olsJNjoqAxagaZzNDAFnvGiJsIWLTLoEkntxsgRnIo
WVce53gFCvnJJkmdaYhg6W308/4ThcXkZ2dT7Q+TUTpvKAEe2vDwO0foHspYl4iLWX2KqDyY9jge
moxvN6KH420mg96l6zY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wvng0RPku5m5MHpJv9WwJDWJ8F5PUKDSPU7V99zR5erdP7PcyDhypTKxqOMHkizg+gEusr/QYxdH
b3OK1yRKUZ44xzg4dZxpsvitjqx51I8wGaS5oiuyKX8hGtgTVrbfoHo6u9pcLQZn9XK2J/iSrjf5
dyOg2xTIXw233HzwIrCKg5RT8dfxa+iICMhoGVZIGJ68DJPwrJbT6Swg5gWMje7MS+Ppwgv0Jxqb
7HSKZuEIyqOKVjWI9mOWG9o9+LBatVHO9cQqYlFkeCwc3YeZbVHELaty1PZ3GYbJhCtr7obXWCNH
f42iQcUXnPWhD7j92uOOj9mnGCfQwEtmFpOg0A==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mnRNLVCxq+sgQJhai+B5fZRsJzZ93rdvyaCrmwTY5fIgoqSgRC5N+TQCYgevu6oU/nSzurf6krRP
lHQ0Ztrjgg2Tj4+uhFcaWXWp3gef6Qsz8XcVJ4aB4xMaBhgkUeweDC7vzOKD05WXxyBd0/qZdLtt
lS8j7xW/2WXeJFqpGaMZ30TpyNYKEPbTG0s7zfxCOI79Vadm9yVGLdGkntvGV8guzxeaRo2Qkmsm
e1+jXsDbdOr2euBE7JiOnNqartejTWUhtjRbkQnS4YCtUcNrW9+ObOoPjivEDKhArV2d5T5dFhZd
vZIU/RR6j3BExhd071LKzolsdnCqR62C9tEZ5A==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
E6549NUXinEnqZcngO+xA/zs1xe2Bus1VEuxweH9iD+10PgNtRJtsG9EF7ZdZas4DjOhgJh7DHf8
ndbSlKTeJx/4QdIH6iyjSx9xrJbjCC8TeQlSsBzTcSKNDMh3HuElLUknuM+x5+UC+hkdrw0waGjh
tjj70YkP+K8Te1Nhfp5PHo+OirttOLZY7Bnhq7x3KDxVSyWnLuCBlLcRqRosb6oaQVAF5dnEKVG3
DDqNFX/V0KONWbfs5QSo5gM8f237iV+nwxPmst+L5casdH0vfnMagphcYI2Gs12f9zJ/qipttgTQ
46Pj/rGC5IRv5Z5f3c9wnJBWRVPQ0uHojBicwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ogp/UkagRFxN6D0Tvatf3PJ+RNRc6aGWLVAuekDtCdp1urxgWDpgdUpLAqv4gVFTloxR/WYTIPAy
tqnoQwfvxF8+1H1sANWUqIMweNpcUZzEYS0M2VRPa5yH9GDRSd+LmMbbrq6RbwvXiR0tPlJ+qF//
xXzjGxQQlbn5MtTPwO8=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WS3NnUM3tGvHLrK1+gyTpPfI4oWwTOYDJPYfQBcc9ol/GaO7Z5AyMRqRkk+WEY00WrbCfviFYMzU
pGl2IHT4VRRzqqLR91kr2OFbN6OGXGirK/a2SoQqoRH7NbdhMzwc2r2DD8mzssXGs2HnjNYorDiE
Vs1axIRZ0Xwgll0Xql9UnW3+H+bZdCSjNWd63t2LxcoNPpatkn50Aa0uZrOTFNGicGTTryERIIjE
tD/W23CkHq3rM2LwJimtfOkZfT6H17TZIlmdf4GzYYEZqzxs/jkYFtiD89KMP+/WhCVPGWSzHT/R
ZumbUYGnUPG9wSLIU2c4b/c9CXNngT5yj0uIjA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
vz/1jllTRUd82K20Hbmgxg/SxjQpatmy9fPYhywRrcQMTJ3GatMdPyHM7nMzNBWX0XdLUeCR/heh
bCer7IDaJ1uVvUNCYe8zWKnNRiFZ1ifOO/Em3YDVespiRcYoQcMKsMyjCOzJxerNuAY1kYiIFqkp
BCLsnsKYv1y6mXdGsWRZCWWanA6wEMAS62u/D77cLf0c94GUK1GaBnxsp/bvjwfWBuhlDxWTD5GL
MsR3tDL2PmIt/+4ACsCukG8cCRMJyGaXecRoMQU9oIS0hBP0OyJhOhRT9RzYQE4yHhIwnWmeZUZR
YNDhzGQ0hDSyN9nv6krq6Qvrh+Tn+vA+haUbW7p8HCLjumCp8Nrb9SnP3VXGZ0163CqMdvC+WOla
KYgvMTctst5P4yOKHpOxk7eeXUkJXkFVvf2r1TvwdcJR5drZ91rt2qO6X+NZ6QRif2BaGr3ivZKe
t6E8yMWoY+V+lqc7/tKGjzyn3sBw6fAu6/ttgDAOBmK8Dxe2d6Ojzv1FZYsRV91ol9TF36m7P6Rn
E/BOG9JGZDLKslJwmYyRCdcpLXaw1/Wo6GcpDan0ZKE/2Cdfj4IYgzA7/AXJwc/UVjrn4az/2vHy
KENASNiZ1/vnaZbInn+HFdM0gDgcetIaRtyTVF8YemxpFy/JFAzrZJJo3ENaM3j4aEHYL4btF4ad
vy4Jfb6bef36aJjExX2WYwwY5YHvD3MtrxsuJyfsj54Hjy+T8Bau9lwi0dYnfspC1vFatmidW5Yt
nx99joOBrpGZ/dpdtqBlTuMUc99Pr0xiNgyDX+8yeEOZfLaGTDnXzxIka7CsXUq30lyAAvHwwjp7
Nq6k9tKNUx8nnNxMcbOcnfPlWHslThfJ6LHeXpgbp1v0HvybfSOwsGCMfBTuhlYrCnT+kCmBnyul
h/a/Jnrt1dTaeBlA0h7h+1Yx1b8rLo4QxYgEPB3zA/NA/M9VEye5C5APWQ31N+7hCPvxC/pFsLS7
x4o6DU2RgkegcBKrLdj+rVnw7jjd45CnbB4eJOwBDEEfBEn1kXvpSGyfRFarVjjMK4liL6qvJBgT
HsRQv0Z6NebsJ+GeQGKvlP8iEJsCxJ6M7JS69He1aeRZHVexYwryItxvLty21Y0kCzSQc3kXCx3O
USaac3TW1Qm/3/EJtozBpJ5jaK0XdbdOruWbxQk3ahFgLRDjWU3CQ4iTX5ULYhO9Y1HbQ7TIGEgV
CWcZr23GWFpLtm40FJ/SjIn4ATABPomL+DlVbQ8RhUsvlkVFio0sXbG498b3/J5kYd79e119vsCq
ArUk5tEP+sb3uctPxzccvJwJb8vlr3SsX87qIIpcnW4iP4xSQa4XV8cmPoH4o9bkJQQ3tUIXczW5
kN/qEoW6ZTECQuT9jE3vrWcSsGhyuvOIHGeEaNR4YvXQyY60G3J+CGi9TaJ6rRtIXCPNhPjBgE+E
dtK6eWEsCC6vAeiX+gnxthd1GfOer1ofVBhpHgfE0t6RME7HzvRKAiMouI3P3Bstd/D8Y/0r7VKI
49BVFXu2rVU9vwALWI1OTEr06uJfUSRekFYL3gaQZU2hP7/f1IG8/UTi/lrdq4KUzURJkRMkqqrM
e5+GzW1yUqWx7iFReypWyijCkwKVTvgYbeb3T/YpLvzyMqRNRwRfKARQSdFdXTjooLwp7hrCAtD5
56o7nc0RFHWOc5acdYvXhVZrGOtK4BCxUrmtlZtxi8HlL/oAVoWVjsBoDmCsztmMIL/deE/764l/
u9pLtspwhZSS7Q7biibwrn2vzBPhK/a7c+cjU3zWJejP+mN+LP6AoVZHGhaBceGYXexk3jnY/DUX
NwZkCnPlR8ZvJojf/D8GSaVJQxvkrR3Vbwnz13029rWqTpRero5jWC0dg1d16F/7qG870K2N3kGb
6wQ9xYgkvd++X3pzktSI/o6ohLci2xnUmM2UIhCHifYqAlGAs+6TplMCfQnMTnkHYGEJ+DcmE7RH
NWH1xLdqwDvdJ+by0pTsIyGNgbyhhmTMeUTBTW9MX0FBjGOiQ2XNOKebs5PihaFTz+eiZGRLlSF3
zFAID5R3fXY1M296wFsldbK4+9131pO/p3FLAejXXepdMZEBMpxvjkZhZg9mCZ6EPaI9w51e21G+
dJn/6TDhmYu6HniBNt0omUbCdICCapGlGy2ga/agIho0fubkCBuIRxt+qyZsqJ2937mPpMN1c13F
2qyFpwoxu14sNLelGnLAzESdN6h0InZO+68HfDMaCaO5uUyz1EQmUM1IEniztyC8QzASNA+OSu+l
Zjx5tqW6Qpx+s9ULFjLkdrUrxuAFXwlpDakG8YKQ2j948FiER2JSFgxXyb+RpVLlZAvMTrQZZYm/
p62Ltj45rhHu5Coo4w5KoX8C6u3R14SnK1SE8jj/voZQFznh7vpgfxAUPzLxGtfG8/374TtX8FRJ
xSNRi5jfkU0EheyDgvBXZSJkwTbXeCYLUuX33RPYvz3UpQY68HnvRQy8QmTp5V/nyELbI8pFyO9f
OrRezJodec1CcNi6+3o7FK/9cM0USNmxC0U0tg2KwgU7SC7LeRFFLgT48un/BJkgZZUvmWeQ52Pv
CKbrVWIf7hMaga27td3S0yhaDd1lBU3/es1ihpv1YM1TKp9CfJsVPrF4MSNmZg7KrSFwFZYTy14n
x+zS0LGCu4zCxXiip7qjt43Qmki4xCFtVgSJlUVyUaJhMvlkCpY8XW/uERdUUqFfsEZaWzANEp9/
hWTzicn7g9q0b/NC4oXt2iCGA7wqGFesNJGUCBFhS3SKjLgpPKuUpbv8vQ2F1MvFVdyTbzblOcTt
veTGz7izkHaWRCg1HR/4yaks4Ljf1nkG/0qgaRQc5Mn0mFAKSx4l8hHW+0+omlvgIDhMbZrbgjhT
uzHpBg2p8WicrtQptXwMcyhcK3PnwJhTeFd3hII5+a3tx1ULxQVNKlo4hGz8qTNxKBOylapYXcQe
Lx4FKfEPYXemtPC7cgUk++yBLK2e6/MbTX4Px3dxBv5QDwcrKUzj0cAQAT3jxq3S4FV/IPzrlQmu
AvRqyEs9+HFktDQQmMAjSmIrGer+uo1LrTCuioMpuHci3duHxJkxyhlx9rg0BLNon+97GpwRSyiZ
QeSKhAN0f1OsRPMrWbhN6NVtbmHWF82PGTGkcYvDeA8tRJildCNmgbo3Kl0uy2Qt4NQ1M57meQQo
EIzOOZ+lJcMmfjhrUgITUrMSyBg27oBWf3UMTAuy12hQrq/e5EyT7Fk7dP5WkzMlXvox08DXWKMW
Nq63OheUnJ8/+i+g16AqjKxxx+EGM2oIL7w+npn/TuqQIRb7MkUTFQ58+rDO+dO6V5l8p/t8lc+B
BdjcI1RacwaS3w+g6vWe6iNO/Zzd2HbO67ric4r/F8ehMot7GHx0NVG3IYP2I8qaYXuBo8VaR8dX
+y7LOu2W06xpIp62E6Nfqfa5c67VTc/AUFzzc0N0kAh6oPES3wlr5BRlWR5drPgaTWO/dt+3nG6C
jwTqSz369sc0h/0KsQRtThIXHF9/X3i3rGnk1g0syxPK7n1eKzrtfL5efazUW30upfMO2L/mdIKJ
xZy8gvPEq/Pk5UiW1DOLnbNeRYcexvb+Co/d1RCN7gGSSp/Mxcsk7i66tOgGvg7BZ9MDQU+nE72O
M1a28T0NgqfP0e+7GLySwMzZgNJzY84G21//qCCYuratn5ng+W2ddlOOyTrUo1M6BTPDiY8fzQce
rziTtQd/U4xJVdcJRJme9ODMyzUq/CK4u9VFPFBbL4AnPM6H8UgZs+T5nF1T3ruPu8wbUtrgSfuu
wNe0hsWa7ZVrF9Ce+7fb8KbMi0kbTFcGBtEuEN7o1SkvDcScrpG0YFg+NGRY9J/dLChmgaRTu5dw
YqZis/G6ckbml1dl9l3SpZaengBK84ARhb39IHgSRSS5J5+n0reU8UP7g3mV8+MPyI9f6JjPXVmP
qd5vbwKA5kUmIGHZil0lmhUHi52BtsHQh9lS2qukUOxLUFYLNqtBjIrQj9DO3IsY4ArARtzt8wJk
G5zjTKc8pGykAwxo37vacTu5E1HPdW9h9KErb5V0V0NjA5vZAhxKUECBNxi8wPkDg0vIuc1gBkIn
IYuXb4mgjmziiyd/YYp33uBOqRWgs8jhku1qb/Qep2Qho7KvgCt80OSJwk0/TxLzHZC0OrIjojM1
LJkmIMDmVeOc8au6IOoP4JEENWFkqH/vJiVo+w24zFFRpTmGMM2xBEoMYQsONCGEDKEoft/YDeyT
Noi8CPCpubFsJweWr9b5+jpDx0GjOqqbTADqKyVAD4F1dqfBYPTe8tRkp+2qBORZd91f8zz7PaN/
8J9dGOyVeMNlRTrrlpDattnqpCQdY2TjvyDfiFRqXoJGnmLM1hXWT7LnHpLuyVnSBhX3xTEx5iXM
vtbJGM/3x7qnL2rxO/2vTsXbOYIKqK7aUtiY8wcM556taPIiwmTDnp4q4o09bjAZ40AG4hKnGrSj
bZDDODovShCTr5ncWyY3kjpANLxnATZ9cjfY5SYD1ZF84XBuS+dSDMGSgSy8mjphoSmjL6Hh48wx
xtHaiN6ZQbJ02p7yQb/brqJ2cYq2wnWR1aphpjDFP2sDAKFWxgN4i65V1XNqRD+CN/GG5jbWNOi9
eBfQlYxMHdDIro1n8odPGaC6HQQ0Ki7mn2WrnUSE/FAYSTYdBRWnb/Jzh99FV8T6WyUjPiiEJk8n
UsagUPjl6Vb0byqRPGfNy24QQqT+hL97bGDYTiIJm+yggnbso4XtVNa+5e3K7v6HqreqUz9CsxlQ
h30gDQuzPRTsyVptR+bUkApnsUIUyPDU1XBKeqevpYohYFaoQdmXIYvs7VtNAe6bxhEpujs8Vlij
SEB8nNzTKH00sH2ApTdPmtov8RMdgymeDuZPubcnw1ceYEZwo8myRS1TxU9zRvq5hgDbVr1lx7G/
MOuvotRD8cobvG35JJDbKF677bqJTgTymdlPGwXJTSwjGWzcUzhW5QCZ12BpiuKe09BYeuVXRe8l
/qn9zDGVkCsZVPpyiEakmDr4fskyYqZT05ZDoKzWqLu2YMIj0nTEr0Rmw3XwSdN/jm5dlNKIwhqw
qPwH57KAn5uqKnKEzayrKc0ZFVdDxuc0TxQLSLhL3wWpXoTNL9omTHAPdCON/Mz4lMQni04qhYO0
kmQLiIvUKduNQ7wXeR87hxAzaio6HY4xKlN6FzvNGagW3yZyvqsNsIZdnA2jPlvtvu6GWwJkfa5I
igPuWgp8NFAaMak1XwsdhdI4sTH6SmkBofIu4indxTac/QJe/VvM/rBLKnYPeWSnRQStoeE+ebqs
ajZD2QllwXdSz3CUpVif//NxwfYBgKAzYu3boynOe5u4T5pHRo4u9JX1MkT0e5cErzuWGN73LC+D
Ft36apXmg7BXHjGS16kwl4R0XLZ+V/Y6Dus3I/SofnaueAnQyWxVUDs2s2EgPnsgIm9C0zxFZUqo
zWS5kKqMGbyYCzkk5uE4ptIyMVq5tfX+tZaGyz1eEOpKJsEuvP6VobVJP+Qd5cyuZ7laAOzPA3wK
3buqfUwISNBIg8XuMHs6s31mWmfO+byX7o+GuXnzGXx6lWO9eswIsO2er9KwD8JG1sFoYhHL5h5N
LZnjt2RXqpA0pW52Z6yzfWOHtsfrwtU0Bq8rjSpEu6lFZd4WucsYo7elMc4zqN71soOcAQ63qzGi
BIfBAQVHHq27kHay5Tk0PaYpXBPqCy1jA5o4qwy9FKhwEchFdVusZuDnh7gdzwt1FBYpMkdtF3t8
4S4dBc/9wmN0n1MDhd5SHTYJPePbrm5S6kQWtvOIQrUcQvUrUV+I5C0sbEbANlUBfw1L82NjJHWv
Fm9KMQCUtWirOFGEkJysrBURocje86eRLRFt+jD6T5omC6Gd3O1AZj0fa9NrIjSb9onhAjyjxQ+7
cBIrMJqfuz8tcyezYxduRJ1zVASvhLEoJ6BAj1dFaSS5Z3fi9xKE599kZEF+uRGHxcduzh6od53f
7j3DD5VWWc8LcW8nMtlhQaUsjLWMTSQACkaVhB93f8fztJInaD0I6M359pTHfGEaSVmV2a5bG5m5
T3UKHCUnYHBjEszc8iYLQLzk6vjvxcMqwEZeW+hlph9SpBJ4jvGCy9nqLCjj2rNTyZtkoN7tTEMk
LJqxcogmCvlQThx/eLe9/9Pf2AH0AJjaIEePRIhPMF2+9ypRhVR8q0KrnaCV6M0FZ7NZzrUiUv5+
r1G0IxGGplZzUW8ZWBee/W+c4TpdUKSt1cJUtEaL7Texf9ZNfpQx5qbbzdwScyvXSgvatqdzyLot
Abz3RzZ4GZ5am6jykPXMRfkQ2P9Uak1LEE/zQYpl7r1AP2cfNIsLDYc7XAvzMX7XXGB1Ky/k/mgD
XEftJnCGEOlfEkqsKJSINsn1IYlMsxsdJd7eSD6gFPSWqVXumcL+bZqJEiQbD+BZdtWbqENusRJF
3uoB/WBhYxrdOI42Tcb+m5EnvDosJrW/GLFvE9fEGix6qhmP+BvBc+8H4auWwZr4/rITdZxrU5YL
KWkMD92i6iIZ8FH+/3/0Ol3tM4Kh1dNpIRSFfPsR4EF5PSI/6vH/73Ta3T+28zADWtr9/yMnJLTg
ByBepuGrKo1Bf5G2iIJspHhpC/xcV6iC7HgEgKepJI8VhWa0aNvp5cyFA1DlSyJLRoR3AVpb7Ud6
Ir25boSZKwCaAaMeINaPeN22y+tCkkzcMXTpM5xwZdlpXKlCA50w8Ke3GCIHIqCawyomX5yVMvcA
QGYf0PWEO6msdpefkdjOZhDSy2iy8Sr5vIk+rJy0GujP/W3dJZqns8pn18T3VflQ6Gx8IDis9D9L
yV2l2/s/dOq6rosVH3Qo1VYgGoYpND3yeeZ/bvt61+7mP+zC1BVgpZDLubpxZ7Z8V+KYKxLOJHis
XCEcRCW5DUSBhQ/qyB6w76CRudR3aDGuhDnrUEg/0jZfcOt2VAZD05aqe55OLYzsO/pnMzVAz6NE
7Dhzpr6GpKdiIApsSbTjU3MhOnWdmnGWIfEbkOaDfdBBxFgqPsud2czI2jYAz9W4gQXwfvABsx5E
MvIjUXIHTKmnYP6X2iO0RuNPXT0fYHE2KW4sVYspgX/0lsjJvCXKruAlrAsBkSb9L55S+FiWuY/N
4WTA2dC+RjqQM4VmiGXVcLV5z7AxjUItQJAdxkyhxZz8teMHtFymEz4TAqA1QQvcOiMH9X+hZU1q
hvZQeXwh1rtbcNTl7Xb62jqekBETcc/5OjhY/2Dm2Tho6rbGTf13GpHDg92Ezn8Socn2o95wVuSG
hEAcITDfHM5pBLqQ5lhMofzg7xa+xsVsWY2nQceTzBtconhnZYG7bOPsiX9ZjtGupOKBNTCxjW+P
Zdof5z0d95JiwiwiR+z8iKd+Nz8hRnzmySToi50ZRY42MWRMiOVQf7NrGItiLiNA9rYD2YlvZgTU
rw75OFXFJM2X4WAhB8GzTPyoni/WnQJxKyv7IY3aCX0/I60w2uTilJuO5zr4DAZcPGe/6OfUC1Wu
qfdDMMVjAJlgBSoYIw2kx0F13GA2U8ERNlRCfQoe4rl8+UTkxTXXC7husKg/20dfPpcIXQ+92+sL
sI5p/Z4Du7oRf/wN2Vmarb2GzRYw6lKmJ1wJqq89IP8wy0cEP4ZPHGvukzd0Eph7k2XsTsZX9Oym
TUgOW5EvvUCTNdVo433PoGQdhZJ78JefMbhQx8QzCOdbN0BvS2jL2z9FoCsR0+DBypicpze5F3nh
oZXRRVyY6l//PceCm8c+nfEOod6bNF6lKA9jwH3UP1OYiPIEkUMNHRLNsIBTEYluHgGP/+5L5I6w
EIgJhXUesm59yPV/tT33RC1MAe18xgcVTFjW8vdj81nMNbbYGr0k0dgitSV8O6pWG2MKmB2tB4ER
ebHfYL3Dls6On84msAyQVAn05+kzvQ8PLuJNR0EVyBk8HEuWbyQ/uJ6rWKJ18e+gE6y5mmj4pxN2
vUClQQQzXlT8r8sljLChteDr3eooS5eFnIBuresi40DA8BdKioVVI6H2XJU4jmfiehg/cvwcT8vA
2ZXCjrRTf70+ZqZAjpxRWTOUaEVi3saUFjIi7g3I5Z4iwHKWiVUB0a3daz7zYROTnMrhHYlIYnm9
oI62AibyhXRTh/6es4vkGZxdfSmjUeHdiPNr6LN3wzoMwKF7VeSgzr1WT/5O8YUO5kXy1SQCyy3U
FBhtvtIMfnAcopJyPti5p7u0ZAM4jElcN1sK85LyQMghBzXF4IWk+HkHzAhJJDDcrsYpy/QQiVeV
nKO6kSK7J6XOGquGsqNNI+NyDO09Ulk3gSCLhwh7YZMiU15nqEoFERFHUH5to2yS1Rnup9K34LDL
QjAsEbSkl0wa1iyrn65nNmBT1wslExeYSSPafBulb9A7w23o6axTFoBrJ6t9SBe3yBuAjkB+6rBl
6tpJi87nABm2/YH/F0UZYmLdWOXCZ+LRhWinoqswLnujKFLXnLI+H56IhC8SXXKDH1ExS9mdogSK
1hM26r41WbhOSzdgfNwXxS/R8AVYuA1+n5wOCAZD/3fuDfu0XUmDY66lMCSpUoR+R+ejKJ1EywLL
5Z7fJY/LgYnAsO+NUHo1XrKZ744v6u9eRCuJODmsrzp4XwAiL7aMmx/vOdSUYjGRwZO7b9RNwgch
kqopJ0mGFIO2XozAewmlpyClQffTULjkGWKO/SD8I71aVy7G3tUt2JxAGHNocjKUzSuEAneb8OFA
hh0DClf4NQDZ8uEvZMCI9XgIIznRk3G0509C5FrEqszZEPYs/U1oiTZFFuMeJNNkuu3RacuIsCq7
ebGqfUKYj9sG+wwUcWVUb6RzZL9Pr9BpVVL27ywe0BuoeALXBKNWKPZyktHKk1r3GriiJcJeyOTI
IloC35epHmAsTQl8LXsG9TDoVMcmPKHNr/GxrX/QPpQ7M1Pu2ZbuiAb5ODld606FmDscQ1gNlwz3
pvjTjYmbeO785+peXKuUQny+iP0DNalJcQVgitiNCzShlFIE5xPYRuiq7ApSiHuTWgGe5oxcXp/A
gDK9gbOJybQXnyiyFsurQo64jtOLF7EOTrRA0+oP0fQbEMC3u37dqDOpzSrKe6ZkB1437FLYiCH1
a0OffY/waNU1NnCnKYwuKjj9k1LB/qmrr1GnbupaH7+xXI1sbGJI5h4lgCMlgZ4MBUlD021Vtyz5
y9PRF8DiNnIvUZ5Yriy5j+6bllNHmmSouu+GgnOAlx69N/OHABP2VwHcxWiqS9i2TFL8uZvRtsc7
Clxsl7J6a0hYF/l2Wq1jrXcfpUoeWv5SyKc5iOhZNnFunoHOkc9lLfznNw7sfrRa5jNncYF77O+q
OkxYVnG9pQXkmr6a0uqk1SmDDkOpeGuGW2U8Q6ougdON7nXltjRp1XRSAS80mv2eOLDGcA4fHdsV
VIgNpJHFX975zuHavb0RbebnipNdkQErauP2QK85yDgmMUB7o4iNZbpuELQ9tqmjxttdOmQZkdrT
8bN2lJ2u6/HPkEWHdSecQWyU+02X3Wg5IHy59Ye4fX+qHbXyMtZx08meUYfAnbIVODJm7eW459K4
F3VajMCUB7YvVVyCLOTJhO+w0uq9VHPJjp8Nm1wGMv6DyH42pirpUZzoZcltuvkoywHizYxQ6gVp
KSBBhfaGZ+kNN6GREcy95f8802v6OaJ3TP5406WyDLPVwwIQXb+9sEjF7ID9hqyRnZl7HQStnDnk
wiJOqoNu8P4+/AkDC1+cyCwZGK2ORCAc3cv6g17EXgkKcucnFAGFkzzD+9H8ckVwYWh4TW3iGjRT
08AkF/hjOcAVBi7QEj+q0ehIW7ELzYNx1aXv8nxNpTbwrvdraNJEaG3eInTgFDxKf3sagJ29qwMW
smKrf/Uy6nrM8C4tXtyIBQXISQ4nC/v2xyqPivADClZaXvE+CNzJ4kVrbr8O3Gz7s13i3PAjZdft
qZ3bqqfUt6PaPeW7o0GBPj/Y/LhwHuPBGItNGz/R3hrK1SqxraEpYCeoJddBp1J5kTDLvMKrmgK1
wUk/OhYIT0vaUHbeKyIPM+Ftz8Ivcqg3d385hNVCQAepG7xIJ6wBIR+xqSUtA7kf1o7qh+p7pd3Y
W7ykD/B5nX9zbdU/xpL8E60un/wc4QKshBT0iuuj8Yuu3AqFLirv2J61opnFpQzOnU6ZPhkarbaH
LvbXE+2i3vk5sxjobGwNZXaal+L7bDLqnREbETwMJIaCDI3nD2a7kSn2nmMifSivwb02YSPSmslc
F5Rb3knvOtM2A7FY9vlYHfPv25dctQJIMwa4n9X91rZ4zjkXBXL40CxM3KN/sgMxVWA+l8vmW7wz
u7VoJogl8HAd0aFMwD1Ip9Fc6ZKh8jHpyHGPD6jdwElLtQZAbea1i2dzUE8zy8vhZl5jnMuJlKMg
/SosuAEm1A0AT+KW+bO3sOtslTA7dtLf7z61yaDH7KcipX/STbAb6z/OZlza+nyH1UxRixesQNUX
q2hY88CPyZtTq71zVaiVP1FVJYfJ6YcRFsF32RlgiXuWGuE40IYZAiaOTnlcgwmOLSdHVJSJ2rcH
aHLecPi2Ux4n+waEIrUQiGkuuJDkooH5QBv06XlITcF+XFGB8fIB0AFcGyDq+kqY5gSjQjvXhhIs
4o1CZRWYQkgnoh04FURgfNKk2bp6MlUNPwiw41nsRO83tonDzU9P4Vv4n0ds1m/ry+nXB8BmIXPO
mjIv3MhJ/rQRN22bHYs4CERV6HkSFSfIGc5tkZ8vdd6J/HHmraR1fN88Pi/OcMfo+sWYY1Mlj6rp
ycfhYFi60mbnbPej/JTvSGgGGm11+hAlU+hwyiJ1s3FBPqPp+vlUrAP7ye9W4Bw9Glul/U0qIDA8
YRkGwgrUm5bv7I1CG/FWzDjP7QydtRkVBLf+tHyskQk4Wnfh0rnwivy+4Ze7mqylug34JUAcXRzg
5dyswmR6G+ZMXEBT8lKRglNpB9VUF/GF9OAKhx49rRlKhyy3MDnIM7lx7jtnqMAHoewAL7IdFb54
ZJaBJ4nuQJCXd1hXxx+LY8HN6i8VsWh+ysvtRV9q8kupWyZMTM4dXxWQ9E7zKh3Zie9BKZiqa7xL
SP1mV6aLvIxL9WSp+iub541NNJITw9prpdEKGWN0nzTfJFEQMiyRHYrVCPfq/U97IR4z+oZqnnLZ
pXjpu6II72ysByObqymml2XfxTw4WcMJSsbKluPfVbKEf3UmgMGNi3K61U40KhFQEhjeHqohE4B9
T4q/kgW3Pl9fAS8Kjaix27XJ2BjTS20/n2MO3vKUaT0VAAv+x/8sItJ1fO9W+rz+pQ32I0koy7Je
L3KlooQ5oY+GSQeJBJ79oEfbRhRCWDv1ivZC8CILA+tY5rLaguq2JoVt/CbFinOKGwOI4v3avszy
38deIEq/rEi4+EhF/WIkrIBZQc8A8PYCqH+uJZUXHZ8oytOgFQIT6sQlDaN0y1s4Izn99haZ6bu7
RJbl4rTY85eeOhoKOfDTyMw8XaRUIOw/mNhmEQvta4qdH7vlTJMNWqALwi/uzm5av4GxBI2G6o+j
JKbmTpp0NPhB6RvS5ekrH9Soez6msMa1890bmeU9G/bAlmujwTx/H9AwYxhBOM5kT2SExykyngxu
ude3irsoh5XaIYNR0ggVj9m3hF1CLCKz/Z5xENTkI0hKeZnfLK9XITjgkP4MGVlLzMLstugUWjAZ
0VteH2jKMIloIq+Gbntigzu/7PZI/7kefy+GCnXjJ2CgrP1eDmIwJKwJHisgNTHt7tYBOhLZPymY
LwpKwEJ6UzReYF2ENJjVLt0DIvlk38fAp2I4J7qF7E4Bsn26xPY/j4NQNXP+2pZQ+deHGeXiOUr1
qpJ3wfhW1xlvri743cyfnEsMQJuF71RBxPnkyfb48JJuNt/9FUNo7KJQB9t7sfWpyQoQs0l0gQY+
RiLJT1mfUMjT2cIeqge93uystPGW4MwbAdBdSTnSjUuor5+9PV7yohfn565XM9Vw56cdSVJe8no0
oZGFoL7wiy34GZ5CgusmOKEJFx0zCSv8TDzd17BtvDt9n1isw5wSg+hmk1o3ecHYYTf7RRF+QU5B
20PbxUz6Tcm4vari4M5MxuzVsQoO/kWS2yvDPapVcQ3QXTfgb0DQ7nsxPRQGg5IcpGPdArNfaoZf
tvnm7exTX9Go5C5H68Ss+TM6ZCvH7x3TF/ks934IYgatm+IF+ePGMQSIMHPvnVwvZIN8gQ+Stddi
tZMYy6xY4B/eGo5gH6aZX0bXeEaUcHLHX2EZ9R6VTnNyYU6jVwbx/W+/jJQU8ym6ZehoUIecqY4K
BkxWvR5swsvdlHLTmh9JjDaZT0hqYdVUGZ4Ra6ZiVHkMC6nsggwQZE71WaXxfn53FH7QHHniyGuE
1OYfTF3K/zWUUshUbZ9xPpCTgDEGJnDJRjiTDXWq9U6EAQKgVjOObFC/ZatQcdx+M3udYHkjdEl1
zmcbl/Daqjm6I61s76+dTqP/hTi+0m7lP191l/+/rNB/xxHkR0kpWyOcg2Q3P+DpyurRcsR2Pt+9
qM7XecvYiHCS6YBRUSKyPzjpw/gmkU9TX2W7E1xHAi9TuIJAaYTInN/J4qaQXS4jsQ3X9hfHOtf0
RsKLjI/Hcre8rDPiw1395GL0UgwduWkKHA6bPslwLWKicbivEO7NzRFASQcNR2Y8EBeWxG7xIV9l
1fFiP6I9K80+IrnNzNwEPwBehJHh52oKULUUpqBsA05cRskR9vvM/jltLxYuk7c8rWJO/usf6nPG
EjoDPk1Hz3huWbuCMMLlvlvonW5e1/WJBLI2ccKSzDGUnf+pAQABX/HwM8YII+0hXGv0+BCrqWf4
Nb/gFy3rdZekDJkhJau2txxRMBYIHiXnnxP8sShvhW8HuW5rcGzLM7EfkIKvlXaO24CwtzRdDrLP
FQmuN+SguVgjEUC/1PCqvz8PzEmb/op4XRYg3Uq2hzRghL8YAhe35wFMbzRj3D4zaAxS0rTZrzVn
/saC3ctAJXNww1MYH2bn1Srn5J8orCXcIA7dhsypsyuXFp/sH0B+PQtOBio63Y8/Zi5c/KKOmGG/
D1hQoczm8ZvBLBIV+GooyGaObNKOLp1B8jt4HWCxZqkc2/zFa0TEVzMvXYA/nW4EXmI8rfSRb8yx
rZjPgkTRXEiR038TY4nWpteEgBuKMeD/v5dcJW4fOAzcSXTy5NpNF8+wB/mRz85sXfakpUAdQMsd
npeeY4fH/bIdAvRy5UfPDJskuJ80SbsKgh6opFh6uDBXk8pAOvm/knVLzeH7pLmdsYU9XoymF/tY
cpwmmNbRy4lZin93oQ4FkZN9XEBdEb6q7/8cLsYO7WLRlvk3/5ML325toJWG/pFHJnCLkuddRAfd
c3MsZucxfcjBaPI15fy9dJrQzbpvaJgELCffPi39zTsoJuQ5fNQg7nR7orspms689YYy+fFy3f3Z
Gtg9RWiYG/AKHTIRX/9wxH7LchpL6sRjTXyMOmD9tJsQGEW7jk9/hb4IYho3ONq64C1tZw/4ZKpn
V4hV7Z1PLzCdCglUHK+uOqJ2KUwXRt58UJA9XYpCpLtiRuon00GahUUowhm3rQxwvuWYxC43eUZ4
qmzNkYI9p1P3+xme6BcfsqVJQk+l1Qzw/4K9BNmztdykH855mBSqmCe25Kk2FeI/RvwM1+I82dN+
8vFc7CAPsdIWrfdF899dh9l2r7eUnWRMG/hY0UjYUlXAAaF9pozFxLqrJlHt2/LQIdw1L9U5+qke
ZLfYCqv91wYUulIJIqwEDAS0I2VEmHISzAgX7RWJBHgVoHQw3byl8CsICez5gLNKXxztMbdXSoV6
HU1R04ExVJakjnx8VHQnMMK+4GlLHE9D+c0VIqiRWbk3tFdMYeO9G8gqN0Hwrcw3aY5fPJlQFzLX
ekOgZki7FGERUFB4950xGipQSOt/NuGd0KSnJB9Ep5yEF3cyikvpdDnraAOCvZBgk+0u9bNOgXVE
aGVGM8vY56vpRZHsFnLWLfhKMPWuc6sfbY4eMxJbUDk1PCBQcaD445a5ege401VtUCX3FQQfDD6I
wrxnFYVBaSm0StLUV9+O1CwZKirJDxk+xJzH+rhVmatZdxQtmu1cBY2teDBZSXNH7kXg6UyIZr6f
QZ9NJcmevBpw4uIiO5kYFtg0zRC22aW+q4P5FYpL8PqzPNhRTouXQg4lAH7yWWp9/JFcKgAa51r+
yBQb3mwbws7Zjznp8I8VcTfj0bD0fNBUZLre+C6ZU6YyBloo6OjGAh9gSvJvO2OHNrWdZ8bsCKJf
I0vNA1Bb4vpbuXbzY9eaXlj1naOnxzN4IxlkmtVj4xyQOwSINc7kfYyqPHVv0Ow0PJHdKM4EdZbA
ECFhiJ3YaTBQNPk4DwUnp732yW+tWk2hcHWLleiW8PHaPbzK0KYKMgszUnuMzCn5cqCNmtFba3Dv
xhdkjlj3aLLhX1ORPaoeMyNg/rpjANcMwXq38jDsPvLeG+WQlQuJQTqNvwCKY0Fu44hbL8euN9Ww
+cQqpqhKZT+0uOvCQ868S2WEBXSWQtgYiUCP8XDG2z0de+gWTiQ7L8wvMyvHKXvDPKzJchQ8489e
4aS4aQhBX8cW0Sy+gFAySSmFWs8yr1yNHmVz8lpvsSxig88Aqm0Cq3rlMFVjoGBNutIVRogzOEvh
/e06ts73bw3stNpNcrJDDKeic//IX+PtcA+cHUKyOBSnXfy6CgXBIq/7Z70K1Vy++aDp4uAE1VTX
w/6Wf1ShfoBwVpZnH+67Z0jnYnuscTt4nXNCEQ6MsILalwwHwkHajvfoNX4XU6jIamCjutCEtJFq
qDvQqlXOXLyn90cAWLRAvazwdTjYOB1qq6YQzPbEys4NvdaF7oizPokrnbaLuvhu89VaMtyhxAwu
Ni/UuMCOQKmnWqm7ejAVSYx3Iu7J7huBnox4AAV/3tVQFdmbjkdQsQ58j6OY/cttY7a1dUkUpd9j
cqaHUijZnSXqWihFQNjicOhqyKxfKx9zyGa8MlFTIpaWDV2zDHteIoru0Jss/1Cnb9niQc0hQNW7
4nqnk4bAleL+MmUdd+cod5x1Mvd4G1oVDKqDvWRbDZ/8TlZmNExUezdYlihhzTLsnetRpZYRZWV9
Etwm/NT0cJ/pEde6h5MgonauCkc7EWcw7ZAfpU1gdTfR7weVgXe0Rgv9H1uxzIoDmh80vai4hUSE
UYoOlr2gVbJpuQejNOiUCIML3VkLOFWnULMfyUieRd83zqEfsaP9jhW6GfrDbmEK2ZR3uAkNDgGH
jbE554BpNrK8lk0msuq346ly9JOyzQuL+ZybHBUnaIrhtLX8MUL/n2IXbM86d3hswtfc8KBGyU25
GJT8u5IjVspKXtHSIhoMBiFKOyj1n4wk/Bk1qYEez1IOML3zZQKNhI5yyq4LFPu1CKZa9CBM8QKn
BYrjWb9ni/q0KEfRmg2mXTAa8Tug05lm+bRgR+sLT1nNi7+a+LILYrnIcF3UxeVJvyHtb45H6b7f
NSQml8XoZbHsvoAGxfgakDYJJJNgN74KCYdRYK2aXJq9Fg3XcS6Ah4v3PPNow12cCtQJP04REFyC
xohofeZyEslytIZPfdjBP7OPK6YIdSD09MjOSYbZp6FUhpIY/yI/q0vEJIPWTL0SGWh5hGVTUZc+
3kuqfS2/0l6Qf1L+jvB9AcDZFbMywSowlUuUobsjV7IVwJWI0Va8WuNWlYtOeID9WhgGAoOnOl9z
2PN0+lyWF49UrFDEutoQp/6lLQNNhl51gXuMdNGwj5HZFCh6Js+HmdQre2tjuxIyNU7j4EwdS0c/
IX6N9tox94sUQDewbMlUvV71p28oCL01DwULF7eqiDHorcW50RPMcQcBq4nm2sR89A5pYc9z76l0
Ls03DNyLE7L5XE3fiikxz5mDZK+NkSTNJHbBuVpo8nRP85rp565RzwTuVI/bAiNRse/gcZb5LOOt
al8i7U7tiFqS1cN3rdmwxyf5j44WERdjTOqlH2HWtCH7EuPLLj+CZ6SZ3BoaFL0EHF3nYN1mQsm5
lo1cTdJvHO0AKywBJaASPtUxZQU08PH6lgpDhJmI8A1Oy7ADOUxe+cyuTBAqu360kdgy3fu1Q8ER
WIRBBsOR8noSPNeFkrLT/hg/Z1ofHHew8YZhGsMkFT+yKt/c0vPZo8jB5oYsl097ZAdpukZZI1Ez
dbpSYaqeG0F7MBsFNFgygx1RhC9ApSpE3AUTCc1xkTFySFqmJq7Ky9PXNh9u72ZQrN4e2hMLOuLM
zqscM0TpCklmJtAiHmhLVMRRyVxK+VKknGXlO4DKCUaZYWVhR0uHi8iT3UqrhU+KP0L+uddIJmPa
qaiGn/mpLLWZeKTRYRzrH4LtoqNpvBsXNWfh/zmA3F+5Z5996Sr3Gq1aQMmaiPhjpbbYqaokRSJv
7n5giHQ9ycS9MKr1G3KSedwPT9TbbEVYIJECetcjtGSgi2nnkWo6J2aLkiEeoOsk5CrRDh2KHUmG
hyg0Lw0aIvCySFeNHY1DtihQqRTzVprSI+fCnEqV1/NUN0mhOQ6ko6a/NMnlAo05huRddx5sG+FF
c0eKa8xn/KyYwj5/1d9t8dONK2GId39JVwthWHg9ciZErrC1ckb1ChLTEEmgJ4q32BtWAVxszYum
pFaWagQsou7vpRiv/CjFoFPzTzSWDzF3P9PzCnfhttHpx0JRpEsXLnsHpiO3a4M9SGP64c9fDNft
Hwn+3YKaR17Mq+lrRfSZoUZE9a6dRcdGYXn4ZKYY1s9CEUR0nQJV+M8ORe8SxbuQjEHyPMaex7Hj
WWK+6Hgh70YXBWYT63mUxZaG2CjeSlHab8nnPHdOW49Xz18hQ3RyR27gV5lZZU6qqKlspsk5fcTD
BpSS/dxTzmy7fKpTTTQuKouwQvAJxwI9wQoNLB5w5hzmCg2XD1SbqOmu80EJxx4qvivaCND3d2W/
oymhmCG3dAa2zqL2/Dfs5ig5RPbgV+dTftqSFzJz//Sp9AW8Rg8GytpCbwl1nrRelAhffFbwN6+w
cYPyB1LyBKJSIzI50CgeAzbZUKcXo8eGOugqdCGFijmRHRhC+ZX+l07Xyo52snxeWtP/aLcqDIBI
eDyxQPWdvas0Tch5Yhf27wxHidi84dl1zNDiEkPYSNcWErxHXX+GCm2qgJP4VDkE2j4hCAJH8uPR
GKd6fDZzFi5bkvyvt+w/oy1Q8dd6orfW3tCkLnDC5p7KSEifug+T/6hnruWNv1MQPkxnSC0pm2x6
9/csUd5xqBQwdW3bty5BsOSSVz+DiZzz4Y3ZWiZx+3FEXwNQbdieHQQMH6OSc8KooAs0WmCqMNl4
KyXL3xe7SNiZZdHgzZRt5wtxb6HM04qZeYEMFpHuIHKFFzOxyJS7/9IVFBqOU4sBcCQhw1JWFola
6Xgp40ixf1SYXzPHT+uXnamH4PI+auijzGiRCPdvPwa/qsUfm1Lrv6ekxGksJYod+7s+izuUaP/T
Si0ezBXt14aoknovNwy3xP/6unQJPFZ/bgvNXsYmNkyrcikAdVMQ+ytct1Wx2H8zcxeIk+hHdDdw
PCoU67935RxLeQtP2nFLCTPSZ1NDtzqVkvAGMZ2B0yxj0sSG05hgnT8+i30sXRaCDhSo307IyqpK
6fRZAPHEU8f6bU5fPMg1OwzmDoHLQWx9bnSj0T4EL9HJPWVBxrzkSBeNpsniWVWlq2hJ0hLcI0bK
y4juabVvPFSqpSei4bzveomHI/SvrEfwghEJzcmhJEMNQroCWnzbUOHvQydDqRoDo+J+p93WFXol
YNPxkgSOJn6Q7dhzcev7U/TEHSeldBEmYE1PLFwQ6PkJGdr00yw/Lz3fBA2kKDlAZkrNqAslqrdh
G4DtzDajkvCSDv4971Ds9C7ynUK7K8jvxlRlSimMPlhcKpX83XmWscygwFxZ6da8+zqqAAcQcdtf
CuLqFtCD3qROyX80PPVDCf8+xPaht3Zk6XRLV+0wW7goqgYmklqz+TWoXO1AGqHtBVAj+FMZvsJA
tn3H4Ukgur5KfNruJhS+IsHh1cRCn+gIozkvUKPfflGo1VLGS+LCaVIVCUPv5fa3bs2BpPhfe2zJ
SE/URk4w+N/aHlaQtvm2EvghdfRrDkLM/jzZRD8u77e/mIcrYt2By51VDLu+my9KC7RF2LkeuiYO
J2ftog6kjMoSUd7aVosQKGYw8IrLJeb04Mjq6c6rqf4CVacU+6zmhdZwdKZ2GvQhlH3Rx4ckT85h
4sw8fQsYIuhzfWjjqSJGeqxdmicDC/mGssp6Bny7Trg+vMg0Z3P7MdRxvRUebJYi8nhTSceO2V3Q
ADWFgQdFzLZHgle5OWDUmCeQBDHtFfRwJzkRmxqhbb/c+Tk1JiAexem1k29eQF9BWLSL/bLvLiFe
jH5g7PaUIslGvL+XoHWUc/0lI9k0K9tt6Xq+qt9vpUpeWkBUMTRfZ8JO56QykwupzPruJdpVhIpE
QlgfTv7vgXnQie1UfXgIYEV8/wn5GE6baYcYZtWrfxpyMA0kuTwJBnBr1txlNqSAhAsCLI7aHA+u
iilqWifz7dDAJyWra08wU50M7xitipyiQu1n17PwVBg3GY6TQ6NlENql8oCLe35XZRJ2bE9Pq8V3
KxQ677bc30SaRM/U9tDGkkTGB6w0Kk9TIWDkOtCgp8rYpY5e33sVrs8bo9OD5h3Ba4Velxq8o4o1
WKJyKXofudNnK51TeJ66qTlTQLNFLHKYZLNviGXKBlbxECD/of4t9JBv/sw+U3h/byVlCg/HMuRE
jZXBKF5+fhcBMXPQZT45dukhjlpaTe+5DeMM3uMmGSBTlb0lzM2hflcWnoGP6UE+yyh5YadWFeLv
loL61wk6ldu27/LY57L1ie1OHM8K+pA1+VIV3N5hogwn5ADIZI1gndpqWWFJCRfAfrGDz89voBbZ
JBzU4gY52cvsGLk7xc3wGL3rXWxL5MLCu22iBXYWbuRBNbAJ4XaSbiNr/gjNbeUWJlDDTKWNmUJz
cRp0X8AKKIoio3MrTrBiDzTR/cBB4yQwwJocKbp5yHrJ4gNuqZFKquJLXKb+JYAwI2ICzhXWbVFX
ForhhvF33UTQ9wm4IFVrGi7W++p6trzoLbsbsqrMnmzvsT1yH/rO57giyEAY3fbmNoNT6qM7NG0d
5OGPUkYPCcvOwioS0nelGhaRPM3Rzqkte27wUBn4tzeXMHh1cbahFYzlvhOC658MM+MVecUaBb/0
89HEU+lqT4hQxQJ7sp3L990/a0zEwz7CC3oEdCeyhU+1mvCDK/FunqFCZ14q5qRoy9LnsQKboMIu
vYvIJSd1xDgLjj/GVw5LDtofWaWHc37k+kHOvmvlYCN0fO+DI5sjiNo7qaFTAEr18vjLrnPxEkDJ
tCxxOIZMsZBIp/weBo/o6aND92AL+1XRrUuM54p0leM2/0+kGbCLd5vDukwkNGD0hUHrdQC/40fo
nC2F0g1Ph9i1z/YjJSuRWUo19qYNhK1BEEtrhKzx/NppvCZ8gWuaacWcQ58w/5ZhHUbEK6JfTDRf
vdL26APnXLDRRtAp8P6s5q2tF9y4cUm5cEPzWh+3gbY16vod0WkLkdPhLOuvx2i8q1TRr+97JOxX
2AuWcGkn83Z5kkGyeyLjSbYTyJiAcuHKEKLKEpCOhm0RmRYOPnUfHXcfSy2W3MickLh+/2/A0j0t
a3Y+crmW4HYEQdnNbaHR159witVaHEps3jD10kbUgLA5yrORKlsqwMgtSqKyR+TTN5jniseCAChP
m/HkVKwRGXEafnELf6wJieX3vPBK6UlXOP/8aJ0zbC+ec5qDVtuktfcFyYkgO8cgBYmseYtk5RJr
8+E2ewEB1MFPnWkB4wM0d7FpKXcCPaMeMbsqwzfma3buKJNIZr2HHv5ewgk5jBJW9jeSckei5Jl1
UOA59Zy0i48CpKZu5OkW2c1vcuL32WHyNQPVLYi6KP1Il3IGZWeH0dOu0KyXlHSZ+HZynw0z0eh3
IIkyHoLNF9wmiAtqNkT+oapqhlUKB2mr7XpotEfzNKC4sFrzG26aOPUwJD5pfeayCPzHL39ZZkEY
6A63Wr4HKIjnWU2N8CJlM2ujYmISxZGZY8S0+VBVYZLl1B3sc/Qb98cBGIagfRMkHuYEovxY3t9M
f3/58o2CUTXOQ1+pAFMN3ageLRiz2SxQr5z9pzMl1BmM4TadUu7dKGmXxLIF17d6ibMFzwnFmnjo
mNngOi26QskClwkm0enOGRyRjg6DNVqzQ5mqVKS995H180txWfSm+WNPwBAf9INCmGmGC0PwvojS
V6MizEXxPiWWZQGB6zCHIj19/XOLT+ZSzF1+kRIKBZxInVpf4bYqvg97yYAydeHUAxmIVhpwN+O6
uEoDNBQL2+viUmq6n4rINAWPFr49XVZwf7WfUa2DRPisgXFP801upx/HRQVbSh/wWuSEeZsepl9f
kkJnYRXoUPb6Je+3BceOv11lc9V13nOOEF0U5XX7NZrT4zTjVJZ8eLmu1xHzFZ6v+si8k/zHucCe
aETJXuLRmcoCCye5N6JzBiPob7enHr2lsKrraIle2v4tnkPOVzsXhVe2E3mr4WD7ZVl+hTaFwPQM
uYg0c1TcZqy+zwpGp88PZbycE7zEBvEGAZV5sJg/JvevWgKYCLbxcyVdTlUPpiOV8K3I5olpSULJ
LCJhO8I98Yy4MBXun19YzngqB4nYnYHBIKeT37M6c2PxrfP3YBSKXD2E5bdakiXinhrsjJXeGWwl
jBbMvFyD4As0DuNpzYYJvvUxjDi2xoLpa3iPQ69k36rfLNwoLdSFfexOVRTc+0UQHYUXNcmJmY97
DTJ217JlECoIGIQqzAr98W/EoiHLFd81awXfFt4vcVQw9iR4yegE0J4PMZFVmI58EHOMrn/lqVlg
GDUL801aNZwXOX7anaUe7wJNXlo6s7qmosDbSiTMJlWAnH7BxuekA/VsSwxWg57ddkaYkOwWJn2M
qs3pom+8vXzijTpCFg9EfrpecWHyO6G1VQpLmqh4VoASOejN5X7nPsgxztxIQkKtoICYYHgewNYJ
43TGYDbE8oZ3ixLAGJicd6sD0W8B8nnqBM00W2VvwE7f1SK8ZvSS9o8GREjwumXxzSc6NKDxYNTl
Vaxgt2EjY7YZgu1bJxsPcpOuj2ld0H8STZ1jdN3b4Qa7t39MHZa5PuhG+XsQenjTpGURZrutXYAU
SsK5oNLMnbtFpR1EqHGqjFbMDvu4ur27TYM1sSeL/axGpupW71qr5BVJM0NEdbIaSqcjW15B9sQb
iLeQAoX4we9of8xG+RqcBI7QqR+iS24mirydjdhTYkIf0s1Jy97MQSl/8qKCJbYvY8fA5xgJBZ42
/5h9n6wsg2f5KAx87YgsJixJYEIdKpYjAN1ndPtFCPbufk+1GydZ2jg4h23FygAiPgqpJKJhDrep
UT942/S6w7CKYs8L5vvZIYZshd6YI6eIzCWxiA+FSSM9hYOUq12Gn5XNfy9fNs6V7KOFLBZd2r6w
oNi684AK0pYPP/738qQs2Y6oq63Ms54dFWuWn8k7nahvpFs8k6cxLREiiQe+w+P5AbyerUmT0+mK
+6GGtrTJVQOPA2X/ZgovB9q/8J6WuGJQdDc1qMIjsUYTLiykar8u6nbSrEc/rl7pJykgp/xSE+OM
D9w0Oro4GKkQNEYuFcHbhCu7M4iF/eUUFZjjJ9MSonOqT3U7W3QN+/rtSzYiCdrFWJRZd8h2dffM
NQ2Y/tTbXxmk0PSn10WAc3P/iSjsHSLoFwW+rO6iR/gbd/ZZbpyAkp1WsaNxXxK1YGU5PHhMLTNw
mBcbGvKquzlteWQ8TQL+sewWzAmjhe0QncuKspjZyuZ7fW3A2O0FCLHlUthvsU49CsQByvocx1wd
DR37gLbB2UBPgGWat0DA0rHAPSxerhj+4OCSJinAzR21erclGRW18YmvyhQI1Zgb98HqxMTzi2c5
5mM5UT/aoBoOzdCXbqdn6KGNamygZ9vgOtQFeZ4sCsd2JqOnqUrsXAOj+ZmmbcKhwE43JEvypcwJ
+NS1z3zhVfWmiwSbDDCQydGwO5y+Z4VvHzwBDUtiE5RGNHccH7yQpF9Lr0k5AZ58l45EHS9f+tp/
G77ox1cxgxI6gVd5Ovm90zGj0iHaoMqoHvU5sPRUj01nTCpy7AbBWKBh2Qns71xlwdK3/yqH07FZ
MsKuY0SHdNTpFKuATRb8kwhZo9G/PZXlTyZGWkT4jkjBO0c24h2b0XmPOQnvW2QZsuXQRx5klJqn
yaEt05yta8nq4fhVFbHQjptmjaL4XtZVQ4yIh1RlC5equD8R7d5Gk1OkYq0ucrycRPLcujHX4euE
lYOXBQm9tXImT8rinVcRkXSYnb/7krZiyUozO3oj+wQbGHgevQtp4fdUltIt49tTF+rWgvCJM037
V2Z8MZC9b60vqo3QRp9Z3rcYnbhQVMAtswv3PRARmbdFgURuTQ7kjoUhzjYeLqyxO8rnwvT0hSjv
bLa6LWlxINVo2ykbDad+8WlKq8q6kMJNKLvhu+Z1ApEjJj/9txTQn0Kpb/PSP/LFerFYvV1CTX15
T7FjDpC9obOjSNMMfljpwB+xu2656pXusxGUhsJho7uV7NmdXcZl2iFcKNky5hk1TJu6ovfc7dxe
1dR94eVradpUJ8UZ39Y8CU/ScuF/sq97Lv8YaFh/5a+KhbYnUP+DffM9ktdvbkEYOf2tGJ2A3OTZ
0Zol+6JK8lbOl87nWGvmGXiMaBnA4Is8dZWz/wGuNXAh0KyAaeULUqCuvKDiGmrVYxBe/Eo5zPmt
ZOckVXqa6SCTLPOGZnQm7DpLay5cqwdFOMuhEA8FtmnlU+sduPuZe5S8kgebHppqAO4OywvJzW8s
eskYQSasSczRwvvkU19qQ7CgI0BrByuyWheyCT8t77Ezf4va45gZ8h3mIXi3gWu6OIAvzdeawOTi
8RgqwyMRLShkuidAsLoUW1iFvV+TajQhywzAkNY+osF43JtE057ZUOp/CZUwAsBDY+iVuanaHiJv
etNARNPQyu75qRQPcannyiYCekD3KQDYT4JwEwQb40B5mrxQMuSlN7foHpnnuXVZMJdRCMN8UiK3
wv7y5C3acX+L0VUjDhQnUQYgHD68Pk1t7eubb3vLDdgoL1ZMEq3+bLTTgra74L27FKRQfH6Bm/Jw
GLBy9aHAlqhPcz7v95WhwwwaLKUWpwylIxqU/edsevshqsNby36O6VYAhqmBIt91bzQ0Xra07dAB
k0HHdjY1Nu3Y8cqj638VFaKE6FLFP8ZIf4BqdHjNK55uDPzugErQVDNRk2DgwlmsEYa7FkLcYeue
fgyJzoz7XGuaRAmnH7YfrFVe8yA/GvhPThk5+sac5ib8M4xl4In7oV/aW5HyQ8S6gIrPRmxM1dco
c2VzM12A5T+a3Yk9QTYWeF8RYHtrtvSuuOBp1zMTW8ygl2bacI6oWPDLw4MKhJcYYz4yhuMOZinQ
2AbhxOUtc2IUk2nSByduVzPwj/4OfTnSSa5IJvR5B4YE/zvZyJSoxPImCVToZ7Gt5Jq0WjL8um3b
KY551eRojVQ6QewSD/o7pLRnDG5/HuvNX4IaKbMHIl5553KFJkF4APnjvADbPJNILKc2vhB47WqO
32z+KjRQtS0CX9qSGoPWUnhUYHPrZZHhCPUipVpFref70hFL+jRCxOAL1YvtvWJXZcAWaMv+CHEk
b1zJpED58kgKnXCQ5FqgODzhFwduELtPqXZD27lQe+e/g4NLkzmW3M7+bJ0voRwP7pn/2cald7xI
Y6pxU3mOm6gbBQIeoZLdNYjr9OJwFtDuVpXlRIURmmfdczSWLCZVVSpR3hli/qhITl10VUf44sXi
yDeidv/Dwy0PIX4zycvQ5Q1ullCIDTGdb2e/DF2FZZwYVFjOvNUL7ugFgQzNy2X+T/YuU6Yz98fO
wtFXcahGNqn/dGISjiiO0KJkz6I1Vaj9dZe/Q+FOVyxiylFwDd/Snn9aSNa6hI7eWawOOKnhJsQI
sVRLGNKkH5OWLyQ0wTTBixWnoW9Se2c+UCr7e92svRdAImNRraYdkC8zKdvZPe/7Dt4aXUk8G6hB
KKn2zTRnB4OypZ12CSeGbTJpuLS/RxexnuyW0HOoRuQSLg2KzhWDEFt1cYVRwqF3U6PNpnw/sQpr
GvHyCnVWv7JC6lw/MFVWpC4IwZEOPpJnxScUSNBe5m70ED2WLDaAUlX5kVwvQFXycAh9hcVzZZXg
/DXov0sZ2eMcQ1t/EwK0JdEcSNBrj+v6vSQFb1jeGq9Vpz8EscY1snlLdvk95c0M2uU2ZY++vFQ7
XnZ70EZkVX5apJPMeyqy5y9HEtaGDxLRxq95HV4Y6Rzl3tqWpJ0BmYKQ4AAXdnM7+DaY7t9+DDRm
LIUe3bO0QQnqS88j790so8LWo/+5xSESBPthojj0SJjspZGg7CFw81p/UXvtPF+pcW05cdl8GtyO
cEcWzT8EBp86ZBuVeqHZkv8zpHtcrthzbBXxMFyTfY3U1HUrcqNUNMd3zzAyF9BeW1gw+ahAn9WD
cEDxxIXOQLksoPNIWkTHyHcgXU+xboWDjBl2mIS7gCIDCPXZAFOsoT9q1N9jfJPFuZVzeZ2MFO9A
xrsgtu3jN/odgXGiCqv/2EcPu82X1nDtUzYxFX4n1BBl6lFiijKR1mtNlk31+duQjTZNnqjqxZZB
6DKEOOB76c5rRjFb3JcUWwb9aYVeqsbbRMMVa4O/5Afat7fu34P0q0NXQIrL4xiSrEP5jAP6MckC
BF41BDiR5ZWhhIkh1H6Y9kCQSNHj7XRklH34pwiuBs3hRURRorC5RqmLO2D5/a5gBbdxXy2WKV0O
drb9Y5alyjI8XZ5eTr5i+yQsG6IoXaXUsXLVFtR0/q8riMr44l64oLDyG8jtAPRmd2wUVKCeHDeZ
cf8qyloatxFDzu/jTiAdClt3XawLHwaK5tu9iLTJl6KrhAjUv8FIUM35O1kd3+ElsGuFkG19ONi2
XSTezU9pYTqYbE8jjbjf88fCrOTEI3MlS+ADGQCA8aIlZEsrI59xkG0v/lmp8CPJNnMHflQ019di
qq0ol3WOBZxa/BCJ+v36vLcbKOmNUI6zoZX2sHiTsEj+ABPJfjizugnf3pNDXe/9XURcXFQV+ogk
sCwYXoJH2/CxoT/11fydTpMF9Ck8pw1iNnRdMWGEaJVHsjEP0Wk9d1qxs9aOvEetOGwkLc6jYbVp
vwvFEX0oAnECwVW2uXAVmH2/lovwG9jVRs7OsFEWu721nsAcu2Js3CEnSEdySmx55GhZbUlmwH9h
J07MFZb47ZuQPVawm+KaGD8Ds4djGmgnSf4L6xU8xsMUCZn1N4BLFNiYTybsoS6HbzpoEziVNrZj
+ZNq/UUkwVfnqBFzcVHTAYvVKXVlyMAL85S32cf+NI83UzqzWupFX6g43HycUO+RwvB6ubKzrOX8
6eqMGE519N+V+OPKL3CWD1gyn4/i3jDN6Slnedccff22wlcml3peYXi1JBnc5p2XVUI/P5lTqw7j
YWlwM0EXUqZxPiqz9EBWsDBtEe0KUwcu6jWmIqIKG9ILohCWHJD/UincP0ioR1lhctb//XsY1SK7
pAl603rbUT1YR6iy9DujBae3jSLeM46Ky5Btb/XHi4E6avVX1et0cmj/0Ao2POMM4mqo8nXWq4/x
bGIqWRp8LwWC0PlFU0O0C5FD4PRH/XooSturCSBc/M2/AwTKwi2zv+BGMvaPYPno5lEscKr/HIpI
LfdL6gW0Fk3UtkTxVkn2Z0aqDlmUhk3pYhesPc6Z+LHEpgMNJGYgtI62uKd43JceGJjYzLDwpzKU
trEjvpj2c34VkMXF9VyU+R+uOY7vg4K5fgG2up65pbMFZuBUZsCc+Upv+honXUH8O/TD9OOEHBVE
D1qneGsDKiz8n8W5RKAKOQSq7FL1eTe+3lL9Omz6PqmyRDYeC1LDnoRPJQUBq02mXvCRyZD46h6h
FfTL6ov8BbThPv78V4GoBihktHlFqmvsEKHl8g1tKPjm4IIRpvQbHtB0dwMpcVVhBTYHz7OMUUf8
pBE+cgFGodfiPqHMdH7Cd9ES+dy2HNTGmIkFX3g24OV41hKYr8ro2arF8BRHbY5ezdLvMDbJt5Mn
9MXVgJRyQ+/35SwfIkAouK16VRqxC9t7RGIdHIAwF7gFLoFNB60iJfpp7NGeZVzt3ZcSjy62SGoY
WU4G3jQcQCiegHcFq2hVDG/uC22U58CmVUs0s4ISq7lZT7+dl8mUXGn6lt5pAtCVgQdUB3jAtmf0
g2dzs+zB1JvewT+zihyWC3wDrT40Jm/T+zljNnm1VVk1y7nsIPmqm43ChxjWzZTAb88XksqtXtPq
KBYEKyx9G1Db6vIOJd+ZmM+hYRbQblbh4z6gGaKhS1LsEN31RgEkwZ7YEivmi+1ZvWt8noiM7E4Q
lRO0dBE0C5Uol/L5HAWBuEe3glSe8e1rxEe1ufTIwhPwblBDmlAIyFmYjdVZeiZQ+MOFTnbDB77X
uLVTWCGt/bVU5HcrpUlpT45fMrjCc72/04PmnHPLZzL9wfUF4BOX3YEP3jWjL/KMtCqH4qk7izAY
R8r7hsWhEm7+zvQZ9VAsTxK5VyiIw4hayOwOfJebr5AFHb2Gc4M5+fR/V67EoCLqviOWzhVBd4pK
nC+6gCiH7eCkAENge/70x/ArximgiM/hgKcQxTE/C6dx3EJlIo6ifJqq5JPWYTUXEVehSqGvooDs
h5ws7VkTGWVTNBncqlzeBgcaTiIu5Z3X8JeyWpOTg69LCqmxxw2RiP1a9MpyacTMcghVzk0rYt3m
MVW/xrQz0TTgky6BeifSFCR6Alndt3tN+0ax/7ZJNxcqhBV7dabgSDIQB9GPBVmPfqNXJj8k7Xj/
53Oh+M3YLKzUwe5gS1M/BRFBUwqblZ37HMO7DQUUmpCaFku6NHtmXf//kMJoA/K8sl3ms1BlnZjo
FuywlQBxQkHyjILCtAKRN68Re76WeVlD4aXQTJc1XzfVld45+vHoZk5OS0IDmO+Cd8x+1MmXHXBN
iobN1QipWUt4zuSIHtsVBPHFnP3xwjyoWXzdQ2qsw0NoP4kZKmkAZYCxIe14ib1xCdZw/qpK2t9I
pI1WSscwIvGPqxoJXttdNKs0d8nhwa5dtGtdklps7dEK7vq7AyjhSSu+JXB9a0+UIISfniIUdS1B
lO4B8x0gI6M99d6+dzLrKAnwNC1u7Keui8SmTptMQPDXgBGOWDOBPdZAVlKCGPF70FzS4JjDN0Ef
AvpmZRl74gMH4h4AKiMJkAsMzDI/jPEq++vxdQv+pH80U3x+tNU1i+tXp+1vqWtV+jVoy8t6inE5
iuAv56eIYf093g0NGSP9LnL7VIdMhotnjX2XhmdMaNfD26mHmTrtI0HIFVc/pAH4IbatOoeIe817
LWbkWjwggw1SqlvNgi/OGba1VZje/plBlPLUAVbUQFFs2tzSVwAx6g5r28bZeHXPY5oj442cdfDv
QDcET9iXbciqLhEtK5Iax20MJxVC52qJ1vLZEQBdUTcI0WcBI44F1jAt8XtSXK8LpS7yBAxDSRqz
Yn6BPCvu7Ms/Qqz0rrrio2uQeJKZT+L3SZqP2U5/mGMHxQ2RfAW1HjcFEyIJFRG/MoWvAqUUsxLW
JImjJOPRIBSAO/ebpzmLz+vn/gl1Wl3uTqOSAbAsIsmCbSy70ja/FX351/KXOlhkh+e8C9Z8iwc2
BBmu9D/RSJSWpG3gQACgat79sth3PqcIoIQTi12Rwo1/7K0zr0W9bCuAZYm7pmzYocbxzqFjQQEf
dsfCCL+O8nYPeYyQ1FaTiN3ijOX1wZb76wOyHH4YqdcCpvZ4QI31RbgJLX2jGd/od++xhUKH2xbp
YTHYaS48u7kS97zt6D0mYaX+d0byQwNesAV3yNVZ/+3rKkRbuvQz1UlqBTPF29nEU6/IxOk0SauK
brkyOeTZGXr3VPsChbQgBdrLfZOP5xAe4uxhZFbVctNxq33K0t2nGfWDCIu7K5bWjFU9HWHpz6Fj
mn82zJV6b7liUqM/t+E5JbxcolAPIIypSkEiwwvhLulUzHpmI4rQkVUPxu/U0pkR+bO0lTfciAFL
BIwcj77c75W69lqgeR/MunEVJEPj6orOnvAiYvk0LCxccfxOZC7orcyXmX09ck4kuQO5YhN9Or3k
8kXLwjEDxyo9egkJwwvkZiGDSMkaJwBS7IPNNcRBuqqD1HGd9mra3VRV/kkNBPgo2v0x7/lq3FR+
KtscxKUno9GV1Whh3q4PPBmIxWYuhgemqLMOAWSaVhwRYELypajjYzYvLkaPykafT67a8F2OS8Vo
UhXu+HSOOdXdjvsUmLHoLEgRfQw91Cb5kqhMR8bdmtBj+Vrbj22Uk9AgitQ5QX/dfGNAqqz83REw
bjs19ryZb/EkF4QVYL4H2z9wWLRWkYXMgKGn8end7DJgbtjG9fp5Dz8Db7+D39pRL65lBnx4fQDc
1lUEZzKrUU0jMCeII1q2jIQ2Wq5TY7LE92RbcE07AF0otasLqlQpScXZibwAb1LLKK6wOB84WOsC
+PxWzAydgVxMJAnfHMTunGcmpxVnbJBLX3WaiQVtz9fdOEqQxCUDn/pasanm6rlBNzI4mCIHLMrA
Rwho2mzrnBMtdK16r8PqfA88nNxhcIGHYwX1Fi3TdocFvg2JoKnlcRgy+O+nro26PzWukUwaryLK
qFAofTgn6oPZe2JeZRFqg3RlzeADUJdDbL092pbjEoMIvTnTVtd5j1HnWk0Yf9NTt80ND894mSal
N3/2ivJ/rELcbft8jUeQg9MSRnQbofOYF3F09yQ5bR/yqZIBov9dX8C5aQzBiDK7DHzBGEJ0i3Ug
1jaA40AAI+EQx2YqHCqH3WrbxqOXQmQ4H4xMM547mebiH9s9T0VzjAH5r7HiH5XpR19Zkt8FIk0J
SyqdS8MsARsQDUqGwLVWBNKCHLl0f7M8LnW2gYitXKStkNIQNcFNO2DNc6gkameeH11dGAdrexHU
K2ZdOMzzyz6GBEZyjForOEwAglnQXGz1G2CuG+qBby8Uc1FyH98FQKlI+Og8ijLtmyAts0rPZprD
YHDYE1vXca6Xjb1nDdSzvXzdHBbu6+rCqEcbNOcoQGID/sBZxy3K9TrLGLKsO+sZ93bZLz44j8g9
gMciQlF2ycmK6Z8waQmZjKsLDl/7BSaIs6gNiFzZkBnlXed+7d9lMnnrBf55QR2dkiiE3kGoo+Sd
QqTZLjJUui5KeNi9xq2jVA/SAOk2dGr2sF1bpYDPqqAhjCoFpvbgKNGuywH/lL9KjFrqiwJo/t4M
K1PSd6267h/asQ5LMnVUTT51Oxu7PJ95U58xsh6mqGhwj4PkBNxkxzzRDMxkopkXz8H99y/WQIva
061DuyJ9NUAdqPHJzIxd39JIkfszm8LbH9XDFtbSDzGe9iNgP6UmlzlB7XuEDbw6Qfbdp83kYRUK
gZ9T33fxksAMuCvQvJrJfz2UP+D0kzq/xptjLQeIysAvLHoYx0KbNOwhGo9mgHY8Kr0aew+otIKn
U+0aQr5D77AtxpodYar2p/U8lJEWUBZ2XvH0V/2AyrTEB0jgLx2C0HmeRfsDqPQbNlCxY1e2LTcz
A1NrTXozpkOxG/CU6XoqM2RxHP6bj1gb6kW3S7T4UWcd6+w0Bfc2Vs3SocQ34G8V5ZcIoEDUeT5B
n766mJyUMJsJ6LwD1/MkwQM/27ogPn5VCAFxal4rxTCAsG0AMNOkzEhr/1EWWHt6jlYwXbweu67+
mP8TyhV+Db2DqXx6AKx2L7J9//AlVqclq4PyXYviIKe+BGAjoDMBzcjqNP8j4RQd8KcbeRpAtaiJ
afJe55zv7UlgQT7onJZ55/fJGVoM8Vlk7aSt3ypE+HiSmfDAKBS8sOncU/7/25EAJgGfSdoyMMhT
GWEalFUtnp2l3uaT9sj9Jwcrky+M3NqBJJwA27FUV3Qe9kN/to2CZDX/puiyd+phi/4unVJErvyt
MNPq6RVUMpnzTKTUTtzdZc/OZq8LKwsBibxZ+KtNYlK7Ymdh08QNcsSDPRV+jqtLR6Q5Ur64rm9G
9ZM4mKnJdSj+2jdRch6cawpkyX8U8pdLQf+t6t302SjIVqIWbbKEnneVRIm9TvE92z0p9db0ugTe
5jbBVGm91ZN1yxJODKJPdOQzzDHANQ0x0POBi6/kLs9YtCgmyd+pZfY9NRISRkbyjbRxpEga0U8j
UBR/UHi9Itm3tf/8MkjpJHAwhHQ8IEExvre3sqkHyaA8T8zpuINPESbQh25gKxC+gLCUoNXAGmu2
w7/jkB3wAH/3cQdeO0mhU9iXTBWQ9BsBzobblnB1nPQ4hwAuukLs1VdDd9jeteO9ltt7fhx1MN4q
sMN912qnzq+h5j4ECy9cDw9fhmjfUMLEAewC0dnbO0+PuOM5MBbVbIW+49Q2jCcCFFj6Ua4tLv/W
aaJFcB+Al+qdW/Xl0Tg7M+4AntPL4v/ZC7IWdrabVE8BSgRdsvtv1/6IHtlJ1NSEuHj/yOgCcIjF
nRg0GZh1Kn3hCFbWNmW29xN2DdO9ZTS9Ja/ZS4pfDRe63HUegon7BeOW+w7oaMHVbB3Y0rretIJU
TQkxG1MpticCKLdLa9AuZsv83u2WK/SQSU6DOX4B6VbvsRIP4/VfNnPeo+FvjsGeQgHRvDl3vOll
AEKoTPeIuAk4b7S71Yq72SvhVJq/i1cZBctmGyfY5TepIX8L+MM+/FkshSDGhLuwqugzIU2b0T2q
2gROuhULw31qSxmFYHqhZzO9wT1mT7TTTSENPS1E5u2Ijt3Bvu6AS/YIK5nDrP+peDx6h3jiPs8y
ARes2yyramOERo65iBND2Mxf6xd894jAt4Yd8r6Zo8+pD6QJ0P2gYrv1/esa2sXhLIzKUbXyTi4u
cg9tOhdv0+Sei30frfFSMjujV+tsWEX22eLnMvZr8bO5kcUXW0QrzlB1/v+hrtHY64W2xg2kC3Y8
jqZDYXO9hh+pTZfqaNSO7qobGuQhac2IPOP712lrPW7bwQ6bCgn4fzGTd/88/AJIX0W4V4crobaj
xxbnwq11VVVlzWcEDA2ZHmeYftwf4lbKqRNIZ6Cwn6sATJsWp4Y6qEUrLTs7ev21tvC4moSmYIB6
4iq7Ri1ctAkC0lDUCinr7zWi7Ez43WIW0TOJjsI9wfx5LU05Ufe7kBo/m7DNUBVP7UjJ/4ZXtPvd
Be+0T4X2ggIOh/4Ot0wsVaUFu0dPpvNpNwsR9805VyBS7AQtELlcTMPaCt6KlcjpeoVHVk6yy/F2
qzmGWv3LhQjCzGy3kLbnzkXQHFWeQ3PKem7aqgslxq61HRlfU7OS1ooOYr/sW2iavFk141pZLkfQ
ce57YOe0TAESxXavwInCMRQMaXUyAXKRwkhOgbd5XRnCxCmk7hhZqQCcbny0L+sIL5tkMNcx52EG
HUeYo8x+Mm9bBPwv7P+Te4YsAb5nxMQjPFxwVI163I97W16LChO1arXxBiNjFejQ18iKOCPQfCJ3
Lx3gvpfkmsH14rw9oRvA9hL8p0nx9MC5HvqtKJOlahRGabGKhuMFGQGRYXkgh4LXIKkWtjK0nmae
zyw8i8UnpzJnsYd9vsHQ2nqZB5/d0jageTs3UD2ul4RA/RPsVDbKbBn9PIUuq8BIrSboksyR+8WZ
5Uc+IrB69oc7R0lmujdOYuUdSI8qXKPCk2U79lEr8iIF0tk8b4d0Dd2wJaTGaTxfkwNscRlRFOby
ZFbkIiP+SXQLyQaqSxMabrewy+bmaqeRhouB+WLnB6LArlLVoFfZBIxvmcQ1TNxFXCh0YFDgtczR
opGvKK9UFNBkJlo54+Gzef7+7AIPW1SZT/ZpHgkB5oVyoZ779HsAD7QO27WxhAvNtBHsA/OEksDB
gMimr4ueGIUmS4lxg2XhzEUuyxmvb+UetNwEkEDBcgunNUxbHxHawrTOwienGYq1WNUKOvDwp9Zu
TNIdI2TsLmn+wtlcBtgnnqj2iBzeH2w6JxG7IklGMoPOuNvsclf1lZg4AnzNBJdpe/+GDdJ+nPp+
n7knaf98JEj+uIZCbTcIAm53rwD9YQ8tAaPWA4JMjcgMgkvIJRsPVNb3niBzHG4NNrXHiUzgvk7I
COG/MtDMjcpX3POhrCC08cqYdBxNqavdcTxIP5PQmSJ6DSNp44OYgk9g+Z9Oap2W29rBbePr9ETt
1VWuep3VCA0rnJHGfn/EZyB6MXnhZQwaChzYMuua9N/PVQX6GywSN6/eOY1rft0atHvXaJ01tooT
GRYPR4cjyJClQpK+yJpO+n7OfhQyVHSeNT9NtuKCZkcJ0koN36MJi+PoU+18Y6YFAIh9ddTyXB3X
nJWMHy4zhwk2MdHTLemL4vWkd1vulDxgr5M3677f9pZGvfkZV30cGKKNMjN5UjLassuuwop1fFbp
vTks4hK1+qR9QoT3/u4CTR53VQcNoLRLzvOeNKygXzZmmji1mhi16kfJlcQ15Cc1yTvOt8QDwh4b
x9eYLQvpXkL5s4zCjbYl5hzA1cpZaF5HptymkIEDydWCHoW2wPNPDtVfP23t7sDKXTw0/VuQdpW0
sisBV5oI2JfthHEJQcAuy3awupFxG/ML4jN0ynF6rkuMApUbhf6RVGymDC44myoK579lly9KIDyG
taQAI6a2sx/c/Ml9gnUmcwRaRiQEH82TKcMRkYV2HIznLHMcFEVfdTmSti60L3zXx3AIulVoa0KA
b6OXwDxhYdMNE8apshDNyqiKygevwp0yG7jJJYe24cK5Hivc8HH5FebxdWywcgxy4VC6BbmhoXZz
gECJCKGVxmJ+X+5DBy9f516C37SScuqqlbyPGojl6u/qkrywicikOrirc3iU+JdI/aQDyln85edp
BCNt0VXDqlArlj/hIhXA4EK14QanjKbZql8xmBOTvQamEQ8rB1Gnq9aVUTcA1rAiHW5V3Z4GnAj9
SaJdy7LC5mTd4uG2ZEb9eovw4RR0bj7qVhvljLSAtsocTAfdMr2UbIZbHoRH+ahewuE02TrQ5hJN
RoJzTpmV6WUngL/R8adkrXP/wFib4S07edxMo1TH33rHZiyxVQQJFBZexb/UH9LcoqtCxkv9Inth
XlzCEmITrnNkU+KawQf2As3cYmaBvky61JLj3p8ofnjeHY+YHuc6/J5RgvKfbrVzDC0NKO7mAR9D
r3da9Sym709jaARCT+3HP7dGuQUePhiLK0zhvdozz7xI+UpaNSYM9765tnk50X2l+i222L3vQoUJ
mujIU0CUTqnz7lG3f0yss8HO+nke6r6pjIuBp5S4Ic4V9AxkIvW5y+OwOSxZ2deHG3UHZjjXUHOo
GaTq9Eh/9JO0CBzpl20eOaceUJlBzuFwBNDjGkCtJoOdMo4Y2WMGnBpnfXw7OQSf9TqP9tgzK9ds
GjdJmgpl14ilb/D5H0GCB2M/NnSOjbQCjqNdvuWi0pPsTwKXH/rR3ekOAWlBjlXa70CbkLJJNKZ7
AOHUzlD114+VFyAz2k6rOAk+c+1Gj5YNPaZQEL7uWo3pMbN7fmyAyseejpQEn26NTq3JsBUMqoRe
GwGErFXFd8RUSuiw/m+ghTEQlZXrElRRWUI2rWoVyaL7Nk1ufzSdP1vsYM+eblK+jZZQxeTaAnVO
jDA9ptVHj/RWGWYDow3mWafh1sk8n7zrSPw0LzrjCFadRdxYi/gipnak6QjzC5/M+0LXY/HvJORX
5p1Q315wVTSf5PplepOBqMJ/7xZvtK09NVd7XvTmmieIQumSZyVcomon0Vq7lDgN9gQzj023YOZ7
jeb0X/BoUKgUAhrjz0tMn55s6TzoFWX/YFDGOsU2T+rgD5CVceqkIWA5mMqU97JRCiYw78LrC3Cv
zk5Q9xNC8GuUgRUPrd1cZnjEcbUBmfRTd3lVrU9RaoGJVtWpYaV2uX6+iq/d80JnUSkoeAvqW6Z8
NAT/bBa3dtB+rPFoJ8yio/+qTOhGMhbyql5dkPg9ahlhENXxdEAGlIiHw1oCkCoqMttr1ik/Inpg
YyuNPQld5WeyELigerx0sSRZXSTHZKNB5m1uCbLMXsPHdgv4vJoshBicmunozDA2N+FKrNNnbbmA
6OercoxZP2BAnX2J9CG5ZhHrrp5Lqn8iMUte063ogoh/IyApt8NoUwVoH3qXEECCgaz66dn0laPo
EPwRV/1nNaQbqGZMUy4HkoF88oPOxvPF+CjjAEFCfbc7yM/CQazZ04YgaKXvgWpvE2KFbIymJ06t
rQ1e9cUCXkXpPKpLfo1JbfIFQbnNxlJKQoxMfGL7h7nvlL3PeYMIhnbqvYEZWmMPiQLjjDOn9Jbu
htXj8IeZSI2dg6v/Eap5Nwg2tuPKhhuC1h4uRYuu5EuKAYCXkVsO+xR5aEPq8Qq9WsPxP2x0jAHQ
3+MgvKeQZ1pVbppQ1H1fuGSd1BrGiRx+wpWVkcTdN2dzRcSMEel78pJYO8yQpDN7nMj+GjCYJU1c
kfT/Kgsk+1oIe/a2lYArVOYNLypdR6CjwE9aHt9s2jGSFTwwWevLN115JXMrx47uUSDSF4BqvuDi
9JIVfQaw7z3fJN3u8Pz7aYmfGg85eKB1jlrVz5jQudPdOAQUiISEy2rC9DA9qWKuN3ZXzDHU7xsm
h4qhOeWd8Y/lqfHu4o5Cr3XvLo+GKmfThxjbV16Bo9jrIVGfoAIs/aUeVI32B4ZeJGh5us699Ay+
IWs0my0pjK4eg2LfiiJj4S0cj+DBTB1C6BX75z1O63K5xXGMKGVhAh0ZyegQgF+BlcESb4IvQ7+b
t4vTv4Zm3mueJcZ5XyZEJtcTa8yYK0b/RWAkiy2R3eWVUDnfmYVn7ogkxD13ph5Vbhn2ba4zrrtd
pxK4S/1tUNpD4zSclTJg2sIEEI6Vy+Px/FN1z0ANpbQyqjxqgItcImnwBBb0Z1MsFQeWLiIU5YuH
NjNIRKJBZ0tV8kg7xpDTA2LjIXR+Mj7Bxg7FCmiNlPuH6F3MQTyeecSvfOSpvwAMIoaEyQs3RvnK
EluZ1EBB+f+vMz1Z3j5C9WJYBk37OrXb0g8vmyZjtc7+Nak2S/odoLupz5TdaW10OHLBZtqSIuSC
LABvPM3DqJEwTanmz15TZS4raz1xE9eVt3HFS6bQadDKbhlwCgtzp0I4e5cbl7L8KWFY0y9qnyhO
EOGDdhEbPZpSe5CuZsbAWsm+4POFpFZcthmQ6wn4bXASmwCJ/orQCy9f+6HgaEGm3BJ2K6gIiECe
VcNNTPTrVPTlA12GhEodmnOsck9fLg5q/uRxV9EqmLV+aNB6WrtmRb8Z9rfYUG0X+0W09YKhesS+
VeX7wQHxmoW8tyYGXP7GBZPVHo52bzE0j6QResU00MEQUz9p1wcfkXSeuIH4x2OqiJ31jfs+xw+1
6ulRqBRThx0wvVJSC90SONbCrla9F1jhliIN65GkLWyZyiI0e8HqkhzKyA8pPCAuLgoaWxA3976N
0pxzSlfc/os3BTP6Xs0n5xtH+VvYXaK5xdalPzKj4PHl6AqiAKvo0GlEe8rj/CuTUKzAnv6bYV8M
uOCEuhnWuCZVr+uEIkn1cDQewjpoXpp/oi0+46ezsDKtIyTlcUO3CU9a9YlOJKYa7jhLaCFhLLBp
5GnFuFSLgs2u6mpn1qsDXckjP+onuItVoP3rgE32/fYqjAYMnixugTh/8XFRzQZmTHYWbUh/jvrX
55RsrlCJW1OvkrSU2B0a3dhIq8YQiVfv5134io4WuNfVxBntsKAUAs6UPX7NyIcbvKpmGXhYILD8
WI/6XCN4XyInFXskWwhA0SDVQ66KsJUY7sUKSCSmXuKf0NeJkos177t8r04xkD/6IyuzKJBzfpZE
GhQ4TZZxxfjY+1LZg4XCb5HI3OWqDPOQdU4tvmV5d9vSxB/B3DTjXoyKpRjiV7WLm32FewFAoqwh
ZLUdAmeTxT9bJoMK8PiIzu2ZWadCas6rw+Lo730t8mUwxaeNfsm1gTimC1FTyRTKF0JKkhFbQHLg
3QInc5wJ9q3X4+NJx3o3YILlzHfWfVjs32zd6JlPlsmxXxOVYxFkHm4QNxVeTfspnUXlSpOZBmwz
j4TVnvCUiX2KPH7Q8U++SL1QLiVtXFnYIDml/iAx8LNGK9WF7oVDLFbnhT/2TknfP2ur6P2cSp94
5cR75k1Ueo+qvTjq5ZbJk1zEZOZPP7F5pO1Ee6Y0fnlWbtD+blSlU2KyN3nmnzQemrq34r/tfGkj
IrDnFFlL3pMA3cOGGNN7kEPHVjpszLqX2IzDaL9z0JEcT1kXBNyjIBlQQMfe5kNB2JUL+MT7lmAu
yIHlE0b7jGzMO30PBAgYFCton4p8PefQmxqpQDR+ytxSPdowZG1JsvUzbPmJG6D+RmOiSckoYF8Y
+aL+nzv9Krw3wX2VZPLZzx5thTzN7nqfnLjcTdE3eb+lQXVZ6VpOmddifJDeFWI8GQcreHPDsI4+
6CNUDgLtqnZlr6axyOvKgDa6p2cggvQDW/N4atnvwyQ7T+zcIbjr8VnRjaBEmZYvjdQpOiQ4MYpW
+JsOMM0VrMOrDuwPl4J96QOMEL4cNGAF81ir+uBrq2OUHIreQuATjepTdt8Pax/roX2SmhFtQDs2
nKbTidEXqxkVNeq8UcbIZtWeRcjTE34Olm/iSnuek39uOfgaTFLbDY+0hKPwY6N7OZYXaBKyeJo+
wNTzB/AG0vvkUegFQJYPHjnm6Eymfzh+pwXGSB7YYjfYC67KNfp/USh7ox4o3ViTn7q6hnJbRP4M
tORIRcxgQg+WXhdMRsmdLI0Mc/gd09k+AFIBrQAYsz+9apf7bBhB1+gKaCaXKrpm5kQbCJjU5QIt
U9WoiIt5E+V90XB2F4N3eV35RtDb1NY/eKHfff3gDFFi9qiDaGIxb8NG354LcFMW0jKwxTusZPt7
7ZZboOHtAa7K9/IPyzI339P3FI58qtEicPdsBAspJI6mEr4rQu/d1Zf3D2XsH++dWyYDuD3X3K20
ToO+u2AidxuM6chqw5Bu8gccYlRmcTlWizkliQ5s5VUrw8cj5TU1WruLMwjUp4sEs8Qdi31uRtTN
dDgWPFQO2nSD0h8+nW4RxO0D0Kk75tPYzCplJ+8npUuOV6hgCqGaLL3Qpj4uYayvS10wurazmggS
h84iRxh+xn1G0rIaAicp/UUSiPImOQwhKlLFQ/mV3lmOrxnvjV15N5JLUkfeHI4vcRMG57vy2uLa
QvF4OXCCUzYBCrcctbf+J/W+n/2EGZv92utFgWQXkfapO4M8UA14x3dUBHSJ7hU0tgxYWhEciG4x
Dt7vK/bmfE4ErdVNTfcXxr8S2kXw/6OL3TWMOg38M0pVBfRYUjBVPtOLUj+knXNA1VWOaoeBn3yQ
nDfVAYrqtg3ZpUpJ+CDFQmBo0dR+lbZfnQ8b7XSKTR9npztRWIKnGZBpDr5gwcEmyKCW6O6syknQ
//zWnzLyfB7FVXqWCe9urd/yFAcuVPNA1zmV9VP4uYG4wln8oKV76klE8rOYD9DS/eXWeZFSbaRw
3xe2rG73tsf5m3AsyvVgwnOJXpUDula/7NCU5vXYZLz54RISis5qXd8oP2ZVjNodBKK+7FSCsK2I
UT0ZH88QOM4e2HIlDBo+wShvnlgPw/Ulscdl5B/Sj7rIGmCLfZXxFemCbivimHFIbi9iWNKs4iYR
JdRAUINWyFeEFs2lghEXY7LgeBgjK5lxyLJPxCU5par01asG4LJBA75bVL18aPOFRF3iI9V89uCw
O5/MKmXWOlCPtLvAK14yUiKGWp2zCNahL+n5OdaeGFqE8SoMik5SBK7ThEL95NcmynbzTpkfV1e5
4m8l5/TxfVHDrFBn/a9F3SeKIVmKSiBLTdb5zpbTU2Xdua4he3mXHzmFi6iSU4YadleaW7Q4qJkY
NBdsiJfeHM9q9tpQ86m2mFkNdnw9jzSPtATFHYvSS8ZQ6wMr50shfLsU4yPzqqr6vYOnaij67ZRY
5eWO0SZ/k0JjIiLS/O3SO0isuGMS0keCzts+a5C3ZrKM6Gf7StVszw3U6qlem+KSmuv2/8Y7/r4l
U3ekWMsDr/LVi0WsZLCGw7I0oQCTb2fb9PCBe/UTiXlcOtJ6onbFTick35G6IfwE+GxiyTxbzuSv
lel09h75FWQZFawy+zZwCh3/POUsBa2nTwwpv5iYEelUpDDy8X6ivFPZKUx828whfQYik1vfzgcJ
7c2/0DvHhQ5FNrLtMms3rl5RFvFGsSLHEvCGHOLTEVA+1fPGMm3cjrsIUz9O1ZA73l6n4fHdXHzZ
sPFka1DefL+wQ2rnsG38s52oSoZntMnsNtOOzflNlK/rmSxXMMy8Y3ROKFWwS7QhqFkqUK0bQPYh
/GhW1f1vWpTodtBtHScZhnpIZEM74Nl66OeH/Cvs/rv3/oYrjJczsC7bobt1EKBJ7Bcg1SFawlJ9
B36NFTHUasqapxQp/KDXdiofCSaeLUlgyqP83oTdBfrH4/4QTu/+MnbhUXPYiqiwkegLeDxNfE8G
pRvZi1ko6qSyG+R9EdCOmhYD9WAfFXe+qKK2jy1mCzgih86T9SxCmsHMSoQeDl66C5cnXrOanZGE
WctOdcuw45/vO+l/osQD01RbHAr1S2bDofqhQJsEYgo2YNpBUQVOk/8RAKlrILxN9OHsgj385cgd
jKrltsDfoVppDFBWJPjimwJM9KPtZMZtCU9NdrCpOO1l544EW5LR0i58hhwRKWdHp89EuAEzl3pD
uKR/IfztRLavY/vCZ8y0h1I1Ckhp9tyHMvcQrG8f9vHO/4+kMElZCpKuhH0fisHxU1+X4nY1POB/
VEaU9Oe8VQ5CZTNR+U+iALBVwyHY9KJeaA2d2C3iN9V23YvMcbSb43nfhLUv4V8q90F0lVOz+g7E
qTF6lBHspIin7A1J9vYBg2GR1dYYwsVrYOldZ27NT4c53im2CRzaTBrdCKdh2mMBE9YcYB4vrNM/
ye1zKINOwSiyY4VB8PVzaPqhmmlOD3Fn0lfr6870rquzAjUAAsRl6YZJcyBVYanw9KyZmymxoRa5
NV3m09YHEPhX6x0sHga+w1kG1KHg21h44xbLXd+PIJCFyx1EKJMXLU3Qw6jSLkuSew/rPP20UTF4
k2k0LjuGrtx92NDjysoP66vyHCY9b6LLywOSkydmoGZxJvwXnTeh6b2R7zDs+c9wQNhvHL11SFSl
R5dLlm+c4Gcb7ISvggVMlAC3rBTZVyyGtZIjNGRPhh/xdzW714Zq5HhbiIzP2+JKiLlnwWCtC3zD
OOBFdU1tkBijj8gPOwUMcr0QGyPNa/P2kFx8kbcl1UeaAFUf3FS7Y3z98cepjCAB4vljz2uAKFhQ
lQ3TpRlE0W46EFrNquJErWt9226+uTJvwFbPoa5eQ9GBEgIKO8dOMV1xe7Ggu033xmcNWKcwd4E1
nOj0Rci8QB/TcCZ7SvdhA29aZakeeBhKoohkHMSmJbM77ISWi3+wpKi3OTjT+GpGuaHvaTCnV7L1
iHBjhZ2gXjWUd6tQ+3e9mTvDp2vVsH7ziU/g42n3R9Z1oqMUoNFxI3MbCVQ5tsByQnoEzCFlUU8w
Y8IbFt5IJbGx8jo3mhEYQox0+YuD7YAUiwV/uCDaeP8kAHrehcnalvOZb+bkpbGjpkSRzELfa4ml
kgLJhjBRyyJXuaTmzweZMiUDSXJ7EQU+vhtIyKy49+jjaqM8JibnPECW2UaDtHuYLpWvrEB3kgau
BBJa05KBCGrUtpfRDyS8vWVteFy7MzvHs91rxcDEQTCqEUwRg8Kfqh+8DUtTrE5NpzWRI9CQiSj6
QgQ7EmNnIGDHwLbNmfphMeWr5pl0ceQ7mV9QIwZrXkfMaaAg2ub0DITkB+nANq1RLtNqJpl6WadV
xLv3ku88yPZbKUSaGGsGjizcyKFy+qCMYevcLG8hP+sYzcpLwvK8EQBDJv2aJG8lfP9KcUThQTaq
QBiLMYtVZb7iuKGgSGrUkxmXigm3brOoKL7ycQx62sc3wsgZihg//1ztso68n7iBuolTjPgxK52d
GdY1uybwdC6ZZtRfnKN7labVIaCFHPoB1QxwmOovf6COEjFvSs+6Ffu66+CbYnGn/gQnto5JDz31
6WKUfwf5NHxoH+o0q2aTRXxJIQVvFJZnGIYajIs87rbqQGeZY4G5VkZy3yOPcHCj9WWlfhFC/+Kc
KY7t6tGaiRtHvr6xBz0Gvkx/t58LXGdq9Eayie1j4XEwaAfMALIDJPld33c6JVXY/QrTgT713I7L
cJba9TZE0sVK63gOnE0ngRxWnFf+yMNuWpsVJPr4vGjGag9HsFujwApRFaLYh23VFLZAHhHsQx4K
QaPQxRwnH+MghxJkUgLFGY95lZpQ/F/Je5a8Axqk4GsbyfniyY5thex2TIYwRl+GrHYmxtyRc6aI
XazbXsjdRW6PNk0IMP7KShsG5ZjRdqyjAO7pRoe+7m3ak0NytNV2DriAfrCVvhBNGu/Dbdlm17Gw
ugW/+TLBUbLLy9H0S/P7dHvSffl50kXLLgzNCK1kq5n1ZPLs0j3R4VplfOnLve46tF3X7r6B8UWD
jggWZSZ3nmd0Bmw/cgd8qNlDmnPG3aqxNMBFIMivlKYRx4f/pqQH0aAwdp5aQ/9erOqKCWUyVxyg
5wx9P3fTnxLd/WS2wqI9HDsnr/I+D0vxZ/4KIXD7Jo9CqsoJ1Q0O5PWoQrBS6nnwn0O6zTIo+XX1
Z1TYKSdBXPPp9uaCaiL9f8aitfBAOH20qijtyibtFVr3clpqJa/Y+JLiBbU8GLGjvQmFQwORzDNj
KpZzTkiJXNZ1+hMVIWmOj5UTJf76tRLA7XLEZUUn4gdflpreUI/hVVrxOnKhB+vyZLwcUZcTV3x5
EcCSZL6Hax0fgSYUS2QiisLp1Y9NSb71M/TRXBhMoD18NRXoXc1uTGBvWfb2tD26Zz0WIRLK4K4z
uZla1D6KPrsHmJgmOdl7kaC9rNZDeGXQAI9gUblisq4EqYhAM9Oxtt23wl/VQYZvSgrlmD874ZdY
af+ZdZQGTmtsanK86b+PLmE7MCdKMTYglZmhKzW2ji6zmVO2ILCncOakPHJB4p9obczZF6tkUXLy
EO6Uuo1Z0vikv0Vz1WLYMxHK4rSn+YGS0DvPHNacvN3seASMaamkmjdQgAev5E3Gj3kIMX6RyrQB
V/QWfNRMUMBY2V4yXtekJC9sYRjy2RiE3R2o7zTqZCo3LOvJRVyX32V90GfirNBgsXqoP4/8Z8Nd
sHhoU0VJTbPoOmeBI1dd5cXncoHbqlcFx1dMxcH8l04MKHuDTcxyHKXNm+UKIfaKG1YXrsE+x8rC
rJrt/VDPpVeRjziLNJJ0sN577qFHhMoewRo7RX2TAMw1Qg1R0p4xktEt0yMU8C1Gwc/iw6UZEaYD
x4GDc8BcEZF9g/TUOjyxg0uUmJ84DSFr5PUHQ53nHbHqotZ7rL8qkuJS9P/gtX3u6i20Xz4A1YGY
W92RIF6hxwa0ED29Od+/QudOd1jWWVcoNSTZChrHf6GSfIs2mj9Yyw0FnqwVaL8RgO2os6cakxPk
jrtukM3wydUBUFfA07+ihUPewpBcKB31GF7kY7nf9u4PHs/8sHd2KodyJT2B9SWLMoVm7/5zY+h6
IdQ2Vgysub6OV45pVHlwjhKfm5a1CdOWE04ExmaQgvE/S/r4qYhAu9S5FqufMBPDpYaVfcrK5rDj
JaVl/VUJcMkX59gxormcdxW1uhmvT+XgUobCIR8B9tqou1t2J3bFriq7DA5/pIoR7PrKIrks+yNt
buucU53ys85mOskVlTfNINnm0sc/d7o0IexlQwg9XZr/X4seF34rFk/55JA2Tt0T3/DAmwo28Wxf
+vZ1KGSxAiViNu/5+9mkW3yMAnX0lhrRVXLXP0GeK4Cz7RXI23xq6eNxW1gaHaC6iLKq/Z6+FlM6
AXepohaaHlfmrvCivoZkn34hOGH0lqKNGfgSSjKuFMZs+5QD4hehID7DluxmSQosCsA8dlVvbHeO
Kw/TcbF0IEGl/awaWe7Z+RvkHYWtuZFwOuQ/sboezr7UW9QGfBLtmIkRoZQnF9+DJZW8Bi1JHqHA
y+Ri3XvVYh7EXvZenNM1yf/6W5dBnhv7weKwnKAA8w3QSk3skEm2HugvhWSD0s7tNcLPxWQ/nzD6
HpJ1VDhNkKk3VHDo+NmH02yIxYna8dYcAHpguFcVlk6271/oE3pJ6PfaNKK3KjOXFwCADnjy0/K+
W6emX19cOuEBeEBEf5JWGwH49zav8QFDo1qd9fkj26y0+MVWekzF4OBHukt3kVSyOYo5Q+Azs52j
tCGgaEV2SuIX6iw+3GwVM7jlvs03rKxb28o6WDgKIzzBkbEhuxnTuR55KU0fOixdo/dIWjHEgvRb
9uzBmsNIJR3ZJ2yxCLoAugP2KVpbtgAI96UYGBTeOuBpxs0rG4/w2p5nLSH82+3/CgSXg7B6yNL9
Ytl10jiugTqErXQYD52DOCubwuXghTV/RpmxDDZAxkQ22RJK5pBJXI+2EIWIhDru/TTU63i6wf0S
r4Gagn3JSQVS8Jp8fs57xDd/YWDJvJnp2qoG+S3C0I36FirOvfinRLobyy8qLolVsMbn6SjQmhl4
VOghG64zSf9c3uQ7vQ57ArpsrdEv2Ppo0horxT2SFhWPINP3w8F26SlJ8zVl9Y4PtzWQz/Xw2oUN
w/Et0PDsF4Mc23PE//VOLv3oSg68D0KcVpRkTZEWMkNhS62XlxfN5jrXrufWHHS0NJKJ0XToxqJM
cXkKg6nxcT/62nJGUkznFKVHCL5DNYd79baJjptSLcnO/GCm9jmspcpMviQ6lnK9aJaQFMRgeojY
Oxq14ukMyJTMnp+ngP0NIuGuXfqNp8enfhglHrVWVcDFLDiQ2Vwn5UPCSgFxD4/2OKY+Epz75gVQ
So4UNCyx0Q/LXYcUiDRaIczUpIDBxPQrmqw2ah+v7SnuFzABjHV32wTRGk/0JA+xE1I9QUELG4qW
jZLXSCohlSD/zybfG/TCEvHW68eiHB8mA6g7WmyPtulISMOtWKSG5aOIvrrjSjdr1c574NCU19LO
3+1VmNqiXECRWKds8KhQ5mh/VVPUkmGCB2WI5NyyTs5EiZ2yDN6LIHd17nb4GdiWGkWM1KycTPBH
eHE7mNTI0mfP6BSmhjUNNJOiCGWuycVdEi7pX+o5+tNvD+irKxVyFnR/+IJYLjHr0+GxKtOZ9rvY
1TI2aZYRjIMnI6xxb7Gh0ifcBgFu/GW+xo3A7AZTgJQ6ogjO8aXHqLFSISjcP0o8SENSkHNDIuh6
PG7O7MOw/mm0Mxue0tPxYphLvSyZ4sP0ULmlBehpqCc8Uw2chm6fPpDK5unrg42Kx4lY2/c6DmrE
UqwVKPC/KDj812AG0++d8nMP59bM6b5MWtB/5M3MkT8gxqZzNmG9xTb/H2BLkpMQU1Od97VdEvuT
gS2MQ58RQIlkF/gLlcONi3bu4G55pCT9nGIsLz9XgaRp3JVsGOCrp2Y4BRMmXytqEHqwWsmhNnD1
nz0eKNOhzGNLpvywRJN7s10lbPwD5HhHFoVqCDFM5o8uzhrG7UqdmzL9D3To7Q8oKtE9VAwzxabV
y/8CDSXLQHZFkXCsr63oxwDPaszj1GxU1+yGl2DoofeLNTR82VyJ1gzDtXruFUnk5GiMZty8SD7o
KN9ApUVK6bPgVu44I+uZAZG9hCfFleO0oiMl1A61YNCVxM6DHmEBP/RMA2Z15VxISDoz2c+wf0EC
80rehZ17TPKqb+08Zq2khJ2eQDAYn6VPgDfgWKPD8ewAjMv8ZIELYPzx3vjxWIuUvGv3rf7EoiBn
gM9Oexz4ZG7FbLlN16wwnkfciDfRPfWZdXWygApZsDFExGnFXq3GrxctR1Itt+1fBV4+1i6G2y3y
A0RUoy667Ai6a6cMNCOTxHCfayCEusxl9Tv9L+KZCKeCRVqns/kgZd3I4kC0t54e9sWhtb1CGuud
GTGMK313a/b6LZGJbl9FOacratPANiD8ByGW1PMuf1Wxr+UvqDkiZdbXHqJA3gQD5+A2uRYJB3//
/9N4VEEhLcMBaLE16NcUueLrzPlTlwkeXVkOBBDXJMTgaZYyBvk+U3h05Te8YiijwPlcKyzc0ePu
bLyuJBPYkOii5yzA1lmdh+rBJ7ouDUBQQeKEIx8aGmUeRuPNth/1KR4NeQ2yT1ny+TfH6zsTH/U6
Wa1H3r2jeFDQOyHEk6zsIBEZKxvI/AJqTUUf+3pMYdCkXN3lxUa7IfMdyXucqchExwjS/QOaa5b/
Qr2DM5xX6LwO8ejprKaosODUIeOv6rfktDxpQ6fKeQNGtfIY6S79KW37eY3EuxS4TvUy10fqRU4C
di19yI6Mn2HcnrpS78IFi0SEAXuKMpNZBHuqI6Jwu6JNWZzkx8c1yDCEllTL2WyX4T/cF1nyy7bn
rkCE6RuBXSHAiUxeBeHqYqHjFUgadjkyWfnaJc9yRQBNa1Y/zk0A8LvjzvLwUJCN07h7Ao6RQs4u
87Qkcbb/lrA4GbGz98LQRZd427YuBKO8w/TSqOPBtJHOjyeraPWvpdH9wioqiCg5P9H10u9gd7d/
cAG7DdL3ikTYa3FIAOuT3XozBvIp2nPcq2EH9lLzhRpeY3LNZC8qwnW0IOByYfH9Vi+NsbY2GMx8
Yxw6HaoVPiMMdnhsqk1IE4Yp/T3WptxyBLXYz6oHVDIcAJYRnYpaf32IT6/pFyTbm6bmlKGlyGP6
Kavp1Fgj4/3K+l/NOtFCOcILEwFM0SH7wXItJ65psKjRxXRyJmRu1+Hyfd5tY/AcUt8dAQOwcxUI
XfwgOWC0eBPd6ujGYH7aoza+29o0bZ5/3Ggcpk5fQ829u3yotxdOM4w5fCg9iht7fm3Um6lbIGLR
6Z/fFwjQU9YwIkuB7os6gVDqOPmRZw4pa/oluXMjEDyyIJFA3KnVgKupTj4zH0OARiWlgKFaw8/m
+VWB+Yt262O6WODZtGWJaqjQM02z1yuivHYQfbweNyYgeA46FRnAgjULjXpmyDfcCtAQgpMG7o7l
wbBVuoqTqtlvrrBX6fdjxuYOcC3mM0DjF6tdPOON2dkhvzFh7g2ehH4FQUZC9Nm8wly3Q3A//iG+
EPckkroogmIGXxhoMJZwIxazGkDRtnGY0Aj8uo+msSnBAV3umQcHmSKPJ8uGSaJfdZggCp3WiIj4
dQqckUu84pPWtUoB/OJD+V2RB6gR6lzy+kfMkhVk3SyN2z/dBRG1nS0aVE3X5qvKO6+GpnXra0HE
09/LnFp6va8SEdGAuosQ5w6uDR9eIVK8c364MlT7SYUWL4gqJtXOXvTCAu0JPRrX3FjUJNTUCMqj
vaiQJAMUd+US1exaMlPV90/cMY5SkZfoP1tb+xyi1edK3u4S9dGlmZnYjQkYP5yZQA4jikSc3vFE
GolEdgS1dKRR2jyPDfDQVpQ9TeoSEa+VBslikRfQscoR/tTYyITfezrEgZSSXjPDQ5zMSjINIXYL
vIc+OC/PG/LF9JNcJDsdDldw5Q2PDRdE1w++ugrUgbJ1D85sTaajdeFW07FIk1ijb7LXXPnt5eND
azF6XQ5beYmRq3x4gr1nPaPBpibTVoy1jTws9fxt+FMY4KDurBdlTilfaKYjSugIB5gp7WxGWyiP
dgnOEQTXeuhLkBI8MCyOvwU6hrgv1CWgowDjrV4NoBTR+hl4FfGVEqoqoOjkcvcmoHnucmyQfQFe
GtQQkproJ9LqObwjg05TtaT3c3lYcYxtiZrKWqG0qnglulZSW9SD6EHcvfXH57TnhshLs5jL7ZQG
QmC7hZoEXq7LVCBziChDdQZNF5tuxro+tOJlF35ZWUYDgY9Aonl6PqCLu5HKhLJGrQlUDvRm9Xk5
OpINmMnrEBSL7lHWFKcyEWEc+LK20CdyUNv9Sw8hPTsT5erkiVi0/qHAb2WVCAVTGa8M3F+puFl1
egE6tRypkiKGPjX1FZ9Z/GrD5qBiT27j47gwfsAxV0nfcgbbZ2LhHohjVF17CCXYEi4zf5h72sg/
ykOT9Uk6eQyz1P1EFSAe9IgzMWgcPSnqOCHyMuEEoO8lK73exX8vzOQCZV5WK7Pd/sXjmRjF8DFI
qjhnpkkxLNKqAfvZCz8OO6JbUx3ae8lW6BPRjKp1FkS+ruyrnMxDyBpe273nzxNbTzar3tuCE9BC
Xx5Zz3K0eS86YguGnFpvF4nLvXWEuM/IXm182DKvt1FeD1VyfjKG2mwjVapGBKYKhNuc6SDL+gNm
kTx2lw7LhUT/FBtntVVR/6Fk3dUCLzZaF87r3cdBy7b8/3g3lHUiOa95C/33yrxUe+JNi4/5EyTJ
FZtt/mqyJCcZkVPJ/JwQf2SnuHWz7IAfGOJ/IxG+hwIlu6zEldiJigDwWlee+RKjCaoII+sTLcc2
K/KKHWV2L/zEnFBdidhW2g5c0rgqLtqRgAM/mwieqvyhpLqNd5kpLpcpPPzio+ogOrIpVKG1GTWx
5Il6dJNiX4Cp4pLF8n7c3PRQ77vWXS7HYeAW8P/vc3QxBgBxfZq2lVsSu1ChEuhuwydDLPnVDFPr
cSwVEb8DEUL+DZL76A1K1DDSW9Us3i/ME/qG2OXkJJeXjpbPZZ1Z091BjkVP2ZaxPY4y76pMW2EV
atFsuGMKYt7B9cFrA8SZirvfDhd/NGILF7GyaSf/WnOhi60gKl7OJ7Mb8SnMk484wpQsGyNAAyfh
wT/1SLn9w3BH+5IyjKNzHy9djuq6u0ffGE4iLaRbPXiKPEmwia+g5wgmv0V+s1d89OJ/fc9AHeTH
9uMo2gJuz8ppt4Gtx+hoAw1rQbPFIpTUC9Iwej8vAnyIR/3k1EA1NGofFQ5yYb28npUfN0nzKWfb
GrCzdYEgECL5PLaiJ0EdqQGx/aKJ/OagkaytlO5w45MkteK6VF8DHlaBov62dZZ5xsrvqm5Eaq3p
cOXf7SnAKaxugeg9Jt3qFADjGkGS3CkEGnWT/GfIueMnGAnZMp59mjkibnupZz6UxvFAMJH+on9u
BHJE/F6kGdCVcFzGC+RyHRLKP5/n++PMasZHZzy09wWCejJn2rxT2JD3DJ2j93byK3jhg+GxffBi
TRRkYdLE3ILDsiZdaP7Glb4tQykstV6UfRRenJsjpN8ogv+XhjOwyHfrG83YRABPqx+UZY+Y1ZBy
+JbaxfeUo9mvWMRdtXe/bN9usTL2pUWvkuyowAJWTIBW4gYlnQvb8ISH3esiSg+qFgUN7dO0OINq
yFcJ0CMib5lVxfOWNn9wWN+/29+KraaYfApBGUzOFczwcJW/3sIfteYnLOKTRigSyP3mcLsCKYJe
tNxRHYXlxy+H0uiN8MBqV33iF/EiQm8sdnXROxQazSxjhG4M6IZDNqyvCpSemgZnEvW91uIW93gu
3gzQpSR0um+b1fQyS5l9/He641FcxujHgYE1jU7ceHp2hw6863brx6cDN3nWNWiXiBZ4bopFJkN5
gmVYJCNFk0QV/U5JWVlrbER1CTsTL5h0+XpYSj23oCzDW7lpU6xFg5WREukpj1xgGOnLqS/rM/06
IIEgby5prFJcHe/40KEc7+GpwkU4FKtQ/IcfchhiM21gC8AFdLXiTPBPvMPPoZhxmTpryOEZEwE+
cWJhB1BjYzzIC7qOJtZ9KZ6T5v3mBXOqpp4sxP5qu1jS2iUYMXcGoQwkv8bJoBLHUFQLLH8DJuLg
pFyMU85PmtbwUWXfSvKG1VnDvjY5CH59gLsrV5O/FBQYOkPx9a8/p2UmzcGT5/tlqnDZeLemWIui
8U3BSj3/gf9jLsWYEyuJieg387pATtg1MoRPpoBXXPCkutFOAxUkYxBrSU+b8xqfIljLLugbatLJ
fZKIIoJD2YeN1+PsBZiNecBvYC73gJZeyKBVE4iZRhK+z2jSKL7EZEE5OjaqvraoUFFlQJyapceV
6Rj0u5/OSdG+1BdvptQ1eC3/RPFhhJCeUznoHGBmHeDQTgI8wAkEbLSvQGsG0QGifLvdpaRkw4UV
ZVNJq4EL3xq5SoFim/GJR3xj6U8+byYK8yzt5CqtdqG1mmKp1OfgmnIejkAQOdmYey3O7YAVcv9L
N3760SjlZbCmHTaq8usA8EamHsaGXrEE8ri8FMBlrY2GztYb4nULqPJwB9Kq05VX1hkqHF6fonDW
Fg+QSVR+5KWPesW6a9E1C9WIHScsXDHomSItLnrxDRnXidH7J6KKx3iBJcjLMJu+maAN3jA5Jol2
v8xesFzLILGS+Nn2vJIBcn0N8aRptlfckA/WNrBnv5EaGfiWjZ34/D2adWSjB+lTywZL6CC98XPy
TsiZ6foXKO9adk+LDI9OzGHEmtu+grks8/I+dK+pxC5CJsyYiyQtSLRzl+bJAfJXd7Mk8sCN4OY9
wTvDzZ5L1wWSTCp5yl5TGfsr8mZqAswsWdtWsRNB38iu/MQkNhtq8EwQk25XDZdVeLehq4kUWXOR
6INZDv/WNvmLMd+c4Lc/oYJ3c1gwp3B9z9FMviy/z0fSqodH3po2XQR3EQKFniVMjPPg/DtNXFqO
u63QykhpKOZWMf9tt20BCO789yn7WXfpVHMhTeqUOuIILiCwuX/Xr7wGNlgQKwHecakWLlJkgLDG
kKfMBlC10IEFx2ztmFidwDxZ5AvjqIh/dFmkMgXTIgljBffuCmmu3SQJ8WNEZjBxkqOXTP5EZ7LG
hmKkY0u4d27jZfakuBefrop4a19J7U6pmXOouC3+sRJ92PJBFpzUlQzlWhGNyRfqaS9nlSWML/qZ
IXK2lXC0X1a2vnEix11Q8ONe1vnudRgvFjbmHFSJpk/ns/iK2PEBcc+DURZll66uRTlhKpp74Z3P
lAfek3JHjc0RCP7KwehoSLWIeybU6szizy5L+emBseG6J/2jRNDy2Wp+UgGKpac++4BrWWCvP64A
W6SmfSW2j5NvlOWOOOv8wLuRSyNKAwewhpUyJAWuj9HgJQLea/OpEIwTnmm61NCCEG5sJx/wCNWd
Z+jFT0Qlq9CL0r5X1AP7g7hJyGBSDOKAAUS0iS+sA+6nrXpiZtJOAbF+kCqawhDxZJKQdQkcgOAK
PQqQ8ynvAWg/jBm9vYwN5LfQYk0MtYf+wd+gR4KmWudaG7rxovnFDBzkt/KJb83YJ30jV55jv5aI
VnfUPKhXRNaR1kH9NkR3HCYucYwCk3cWAkbvkPPAo+3Imu49uAdJj3YanopXj6IxQ7lE4WWgCJXX
gTIDcq2Kl9O061QJ/YpK+8dmxSUcua/+Oq7VD/0fgfs2uGd+tLNPQ1IBkqijq6j9HLajf6akHTtq
OR6M5vbWLHRJrpnzYN1Kw21/WLucGWGhux2hbFShOLrgxCCEwVDe5UHTjGmUrFUXoH8JwFG7I0MA
kdPAY0nKABPGUQN6oakwdxTxQw0eM2PBpz8V2lJWOMHhCPbNralo2Mhyi6gx+THRbBHM19Q5N0hC
EYnGBhvuruAu23IhzN16oOYeXWdVKatbQCu9M859CRpAjViHHzKBqx19IJvvthpmbgwdraAw713O
H3Lcktk9q4sZ7VsnMMgK/8IPv7FT+Q2HHoIlFVUVBvXieDHAl+CO5mmDzJoCba359L3gWMFX2Vw2
0ivpg2IsxppWgxUgHlwTie0z3gIOJ47AnGrruOD6hGS/kW/nxJedY9UGKfP8E9Iiwo6vbX9jCefR
rkPsxhT4um4vSzL+gxc/SJsbFqOWPONRzMjISlpuGTo+3r+qQIsxYoPRehEDjuMzGYjvKVshKW1G
N+tC/ZKWzFobK4eVsxsWi6t7Evg7jh7Iv4l3qTQYtQ50HM1M+ZY3926XJaIwBx2uewt/sMhJhhAn
kPe1z9rZR9lx+E7sK0KymqspHd/AT40i0IpBtBKkWAAaw10ov4FY7fhcwxfuy0lPniQ1gnDWwssM
IfrIUKv8+TadBT/XUDJaV93vjg5T1lqo5Kn5w/APFM2RUiUnR/3e2lj9kOssObB9YK4yqVRuwUCA
ae1g6shH4Jw4iV4RGDFbPWqKyG0z1MLsdGHPSSc7rSTbBGkSVxuX/uPsykiWgUVjLlyxsFhQP7i6
1qXuP5Srcalsl94JrRoy08TnAPnr4vRyFtfJT19SGc+B2iURngNsPne3j/9sCBFZZ138zVHeYuV/
0kRqBvBy8KDosFu8CfEHJkq4wlJbxzjv56nD8mTrTSIZlTU0kfs7BSNYyDDk4l8/RgxNI5uZovvL
ZsXzsk7rPyoL6CrR2K2lSIyh5vEzZZuDt3vb4ypQx3xTvw6uwA121Mtmr1WDYs6QKxGSDU/nI5ki
u8+DwAdZkjEXtI7GpXWSYMLHUnhKU3CDw0wnpXrosB27IHPucLkux4yqp7+J3bdRgOrnXgKlZwJO
G26QR81saSo9EbYR6I2TrYpM90bpHLpLFqBNTz6stYumHsGdzujQ+Q0tWvc4AfH3+XhdmecJpPX8
x3/QhrcuTpqFCHvSC4lmV2T9cgskjhZ8xTw/rG7O1ibp3UARkPJ7o9Ah2Ne12vGSrnTiO4kBGoBV
j9HDmJLZXfhjUnNQf4DZ0UePh30RMY4GcNxrskMVUWEkexW0aWdCJTAYuhZMQHpCtzd+Q/mWu3i1
UiWuuU1EuX35hKdiQsFz2OvWvmspPeeGwrPTNE/4KEgnvV1+q4CthTWYeK7LjWTdHAz2/uu0ZZ5W
uLtrg6R0kd+P7e0lze2vsvJtEmwVJbKsIHVCMDr2mohypm9oDyR0lhEdWD02UEHd/d0bomih+8Tv
1jfDRGeNuK4NysN4Xngrp9m5SDd4xoLI1JoOEt8li0m/kxjHo9rOdGq4ahd1Gs4WOlBLee1CzzQ3
O0T2s6S6FEzb9KlTfpliGIuYNT40d+Un9afkFUmDWwAKtnix0wwPs3YV/SC6lv/eI2wifh2G+nuo
2vffuNPeN4T855OW3zcPH/8W6kBI1aPjryJKPGYjORAoKOS9tgTlWZuGNDdfty6iwo5tScfvUhJr
eks1TEI4y/ZHJrUNofJZUZOrWEBbZvpZ1q585cFsp0SpCOCxHP8/ZjiKWAkiSmHPPtmrnqSjCaKx
Fc0j+VJ9zEqFKDdbp9GT9tVseo8lA7d2qGaKCTLb+sWKO8bCZXbEHt4S6uSXj/T2sp/yEZTPmSYe
r0/m5woxrhTj+lORyfJAYHHrlBwvrAlQeRuj8pJRjI8E9HXw6kpPLgunL21WGneyPYYnsBz4rhQH
ghcHxFLY6t2lf99rKnlMVxKGBpCu/TyL6sUBXkU+4Q6VRmUwcdZKYaapZhKaspw4p/tEBo5RxgrT
0RHf9nKpBZ4p+r5DlHudiv4tvJwSyW0GFtPKUOu/HVAzeQEClQr0dAk1vtZhmgqkr8VJhJ6iQQcR
dloY6vZ+p8BljMvCpNgZ3DAx3ZJCkPrle40nJSjKocgV8CyaOlZM9PkqS53VOr/882Dv/q1JNlBq
4iL5dJ4nuC1YUrsujVHY7s6T1yX0hdtvOLUyIeqTSzyEtW/C59moyU5Y5cFuc2MCKxQZfdZdCJoo
1lZCEHW0Dv5VJZIdnec5qB4WywpwzUKd5qY+nDmmSGU9crgyAWIf0BJQkiPndScrFCLKGS/F+WCk
eH6k3xIbFNBQ3WCZrOoN/LFnYBXU6fd5AkT30IPMiOCiZw6+gSwE+AkemAnFFJUhnIIUsN4YCRqO
5NURyk7XMXDjnY9FMiTdmz1CHfpjZ1/lehxzwDjgoftiSlsSQ8/AIFsZAS9Sqz2924sp2us3dT1Z
ikaTadyuRNJz+tgv2qCYee289JRitVLGZ3tDXc8vTcyAOxouwzFGm+qm6HjWRG/UX8PiKF2Rq8JJ
r/MqBsBRbkOTT7kXE8UT9PajtTdjCj9J7the7P1skmzf30ILksXFogVh82Nz00UDtzY3Az7VLi01
43Gh5WM9UQthnAcb6l6d+Hs+aNQqmdNL/ggMvwiK93eByHkFnIQgL4JLdRRbklP9xBrY/K6Z4f7j
p/WB1Y+pyWeX///W4jTr/ScFH1+0AGyLFQ0GdYUxIPUU5ps029PSKHJgIGqUYmEV5GiiyXDtnian
YmnBdmnprcPKGO3wdR11/uC24b/OZXJYenDDoF3k3cN1lMh2kFBDNCCUb1i2mrzg1J2ClshY6+xX
69tJhrpTIpK4bcqpfqHolC9H/yFLtABXGBdmyxuVdATbYX2c/tCGplJlW5JWII08uGVl6clhs/c+
N5IP7zGIABRKgrZVAkWlBRku7yucnfjWD982NfKudx7h45tSOuEl5414PGy/lBq8wQZNsI9+K/Ey
hTP9pS7hs26ZmPQ0N1C/2tEUBZSw5S4bn49sxDatYwL7PpBTbNT7TX4vWuPjnEhWgBfejrI1oU+o
IgAIuL3PnWONAWsQ1MHSRc6q3pgfyvgdoTSx6Gwo+EUS2z1tubso4NIJ32k3nT3nel/6cXd1CzZS
NnNpfFL740Z9wJccEBOjf6S61X3zy3Zirq84DT6uXD153N0F6+54KhIn059wN/C+dV1blV03af1d
nqEIj+HlLSlY6aHpEHvyttuO5GgMMbx5RqcCni11/0TJZUSfKaeZcAfeocspjg9j4t5hSOuKpQtd
7qTkm2PZYdEmSE0vMjAaXOBpyobp3u/p4ykAQtB6b3oRF4vU49Zhj2yAKmLo+tPKzrYG3RKj4de1
rYxzfParQtuYGJ4bVRZHAyUXbiihuKYJf78P1YcnAg0qF6shcBiauALxNfYWVG6i6Az3iU5VYvUE
w7dZZEhGYCVDxEEjG5giq4mhTBuxzZfXjfOe2aLGRTFHSPkTlaPhqoS+qxmAN95RCkpqm8q1Rn0Y
xZKT3giKPuoAc2BfGHNZEn56Z0cz6qDFHhhuSN8Knna15JY9kSJu89d03xZYvncjCqBjUSPgFPDG
Y9hcS3vQn6RJjqkw1tKzK4shCGLqUwqUpIGap4fp5QFHVQsVu4GgATk3QLZz+EJZu8NB5D1pXxBT
T+LUlQkJtA4Zhd40Jwcwd0idT0MEVgOdYtlkkK70CJ3l45mK/jIjZh5Tm2trJLGvI+PxXJXjt3mM
/qQfHpvPkNV7dL45r95KRV1QfKJ4qvpWWQQC2IzKbnaUGuaomOnbnPQa/W3ppE9zW222kfQytLg5
fPjYfnlO1+ytN7EodJp0ynT8l81FJ+XplfoMbm1VXYx75SVdrCJJlzBv03UYuuBQlg8cl/2Unpms
cFwpayH9r10px6GKuCAq3bGAXjdM2Dbc8EmP9vfQZzw9J5XMUtg2wdn5ocmPTiC5n9wclIWGZrjT
YQI1xwWKd/ErY8qLmnQlDWYQbecMIUtC2//xcZfP4BndON9wtG/K726HeeH6PA6CCDdSgWRQL8Pu
vgvieVvZ/0XiUlZKafityvt6CVqCxwwVP+t84kMGVYQkG8z0GmHu/ipffQ5Y06TeQ9WYJVsGl6fH
pTpFkbMXfMrT4TJXPGV7ORDWjiWz33sOUuZ2+eWXGJeSlKWUrwhQZZRas2utGvc03L2asu6Ivu+i
+1+mnDhL62xr57IP+ggJyG5jn4Dhu3y4Xi/uRc961o9w1alayoHYlSziFNPst6MasVXF6Ej6w2GA
flimsXNvlp6HzUEkKdEEgzpjeweGzRXCo93Q37jxf3Du64ktgaXODuMnXn+Qaz+mSRfTTI7fkszR
CAAVfKEy7PbAklUsgEr3xwd59rCiZ6d3HIZn3L1uNEdLo7s/KGHnWwXLVkcvvXzEXrN1mJXX8DRn
9RICBMULHpBpoZ3X0mKkFNLHHRNWduBCnhthqtZ+oqeilmHMQcSSG2nuDIo5lUvc+dc0QQ8dYf1G
NwkezrYRaA1rboNJLTo5qgnsN0XV4ouzL8mz2La9VIcG0gCli9ngJIgdi+lG2PNPvhLIXHZ32ar+
o1f7heo+LgW+9+O4e5VIJ1mTPG+NntG73ax+e6arF1XFJiFiBQJtOeA4NGmGXcNfsz/H4CKMsd+p
ZrzwpgHhIj+HrSAej9Cxm7ERSbDOGYc1bU0GsMdfWU1QEc7zqeSMn7JqQxa4+NSJjdiUpY7+1fWD
0wnxWNmAuVyoD/falsTjxSaAdV+9hzNV5e2QYmst9H8pG5pgVIJp4jE1lo7LCxtMsioFWm10D63y
uS8Rk0CLt3bZK8vALEI9HPEPqrt79vWknRaFMe1VJg8mBCPPYkzrbg26Zv5iWZpPK9jxZH5CCSck
VYN6x52q1haAc+WkI2RhitaFuEKjcqTkYVxxX+Koby9S6RCvILU7XqZI3bniWVCHL59Sbp5G0qHh
W8dk1e+P8d0j9Fce10SXIN2kAnAr3pK2aqxgOmI59S+sDTyqHTXyKTyfD5o7vDZzFCFI7sH+aRfA
Vs/WyIaPreZhXO9Qb3+0Ztw0KcCEBfIOGCJV80s0yv+d1lQiXTSyFYf25abQchPS5EcFHnRz9ZgO
wlCYgz6u3pHPgsLjGLdrjEsgj053X4hb+FgUf8yettjwZVLcXzcy7wpXA4SkVCQj9AA/+hZM7lKW
1fRgi34TGDsOjsuQ2fkGauTnbElunE0aoN9emn/HTW3GJJxr//rVmbhCV+PGuR6VBIx4AweH6PJQ
rTeWv+F5tUSwGskkZ/OcHASnv57eEeoPvq7eni95bvCBhIFFQu6sE4WkkWDyQzKDquSlTeJnWKBS
toC2Fihlflg4YXlRZE/bOtHXJs2eN0/0+3eRcxs7m7BJQWqWcPvEakGrpA1zAJtK1GyJRw7XtFHS
RIu2lyCcAHJoLGyW3kxsIsds7Da5Q850b157OzQ6pDT6EWbyFZjMTxGIzn3dVRMnaxa6yECyVH+X
ZHUqq1gtwTXBdn5+7IU7UmJEPKJgAEQIMUZDOc7+4NGbdn8A6lJC3xzyLYLb7jocbjHZ05ZvjNyL
P1FG+Vm7E1BogzM3+e8KmTaIHkn5ZxABun08U7KI8ABbY1VRM90flxhHSx77JcoAzhaNUtdU/rJu
6SSs5zTEJXgcJPa5x6lxQheLB9dvLh8zfqoPRZ6ofOLN+UDqX+RDwSrSaVLZdTILCtyqfShrl7Oz
9XwdfBSZy7zTLkdMnGDHpN4OgJN6uGEDS81B6wBcbeUBf8I/xzFIZnEyWQprFaZ29qGHPX4u72FN
IGS+F4rpRhm2941F3dN4h7FzfrISeiNcuEKjQkH2IQltX9VIT0Hg9LtPf+1b+DrD7RjUH6jVEsRo
kcHL7HLAitsA7I+SS3+VtRVYpHzuZmMXJNlrhavgy1bsZgqhLk/gJvyQSRpVXtJXsVZAoAlP8Zuq
sTEhs+wPfbBKAVeyLQqenAOFIdm6PG0QZIpWQ5RUzis50Lh9+fcNPSssTwjA5o1Fzx8pHy7C+R7d
TjLNvotodTAil1zUhVxOsgFcyAyT98y7OVsn4jSqj0c9511RyIej22QlDh/4EU/kN2l3joBxmzgL
STtzk/TS40Gb76OTmJrTxK509I7lEuafjXb4BB2knS+5fSL+UJKSIrJPVPItRHKGr80h6838Lts0
245d5H3EwGrPPjGj47raNTUM7GK4HSKvHq9UzAJksxG63z0NgBaALP2N7DIG7FMmo8HCYJikmMub
92YnFumHCH3NXt1CBQC/43DCLJ2oUDyH1qLcfTvhaKqVzdnTJCjrsNrQ/bB24g4KnMEtc8t3c1NK
DAp/SimP/4EKdqgF/IDrQtRLcUnJzLWmbNR/lQA8c+KCDQNdTtAOKeRrxbe8vh/FRxUmg9JfETvJ
YxmnN8RjGZkcn0/NA0fY09BNdwj3VgWR1vv1yHoyG8BbmM8p+fK8peHz0Y87f31EL2zqZUM8iGXK
yFhoRGtsUXrWpMEqa+Z7XwJdNXV3jS2/8BuFaxRb/Ycqf/jpz12qxmhnKBOsRtB7qnL2ApTI3YZX
M5IIGUtSD28DtGojcB0G+rlivTF3f0cRIFdWRLTK6S4PK7YXQNY0ACF/i0ZWFUdNt+1HCMl6KdVX
MQYXB6nU605NXCtKA4ToB7K9ZH4tAIQeIZiPB4DqIJoHGgnWB2OyoGXQ2nHbTZbozA21M4dYbr3A
G1mjS135X1PVuz/Dc2E1X4bKZoqtFkQuCvVMGWZjZMP0UJ6YO98weC6EC3UO27iBe+wn2WkWvEES
GEMJboXhYCv7ouNTI1HlfoNCSzRdtP0zNk77Wt9+oB+gqsgI8tT1hBr6PGg1qbLdIf2Dxxes4HZn
NHVshTGdtVM13SFy5eK+UxAJ2Zme7TVqI0MkRD1NxCJ6s93pxWWjXVTu2kNKVI2tjAXOOFbYIeFg
k1+2YQWaliWv52HscjMeUyYUXIHLC4FZQDOSHZUo6MI98718B0Ba9blaAXDnfVMuyYJRyclTs/zE
XheLYpVqcTnOLiUWgTIjfh3TlABiylDXaIMGv9HCpIqmhoxj9UdQ8ghq9EWXWJ6XctyNbliDsDKn
wO5+zJm85oy+LzKTrtM1snBgMFUP6DDF8WJ8bP5pAqkjD/wyCmNcqhnqpsA2Y662rrG6550Kfhvx
6IojZhlyuuKE7r+CB2QadCk8mzG4oDEi1P6rp6cFMYdEsEXji2pmPLa6Avmu8UGmjyy2b87U3b5+
QrHT/SgBWtahBCHqw6LTrMMLKHnCE39N79kL6HWnQ32bniQcD2UyqNeILyx6pHD1/heY1fiX695T
/mqsng/K3LOzVVuRPws7tCmmSZsX3VGqXNmnjSdS3elR8B47Jq9+3vkBuPrtqKxImkVi2yQYrjDq
YlLrxLPpdXSSgWFE3YxFkoeVuwQRHLsbE9MjrS11ND351I/4S97UxZ8XWULsliJwkw7XXVRD670g
iaGmbTPH/ARDL9beP41uSQzkejqff7WAhE+YTnaBxJP+kLjxbk4QyceuqRFWt4BHKmDLAv4aef/r
pVLSjLDvIjl7PAqRO/spPs5itH+mmB7IPZ6q4DBbkVM00COjMgY8hAQqnfYC/ezhkG7Rll6qjFpS
VQo6so3Q3B6YwK5n1yNP0FRmn4C+wt/VMS8sZ6G+YUmyHSAidaqvA3k45KSc06HGTDYqbXXRc36N
4sw4SXOyM/7+3hK3NH/vbXE1XOlUwmxUXwmicD4sGwoVVLzSWsSIfubylBqXX2PzftDQFzGViMd1
JaiRd8d/zgWkGbmIc03WSp5MWFzdRYJBnCP4Tb0QQ0Qh3O2Xqy83ChYdbPHWmxrfj2IDPo8JCy3d
hD03jHaNj6cc40oJsV6dmDkKQVCaN81jkcYFr1lmIinSbur4xpUIMsU4FVZ78dPW7ZwzapAjpotE
3ohlPqeLq8Fu2McQd7lAh78PYptBmzaU4pDbS4bN/yScdsL8K2p7w8TWft3CWbb3LG9tZOaZgx9L
O+CX2+LEhML/7rsB4h1SZSYk9Wn/fyqD0bB9PtheGnzlYFuvHhyFjGem3LTZ3lAkwDIL6zHKcHnd
LG4pKEec+k+AXZX2a477jTinBbczkjaSot9oxd/Kjr0dATTNnAeRCMFpVNMXmROnFsG4RLz71tjN
sc6HtGsUinubgc8k0EVCzCiW9UIQqntRbjiKqycDEQkJHaAtlkjySI51+zU/sQPmooXVdjO9DYPE
SrB6TkgAWvk1NZ2e5lL5u8PGlAUi7v0fK52ZGeSL451MKSuCXwmfII570yXeRuiSRZJdEI0YOC8q
ME5Mbi1rBC+1JpQb8stF+YGRqpeN8wYWIkGOuZDhieuQ4Y638+tRGyXm8DgzR49kNBHz59m2kTZs
VlpDP5DvBa+IzkeQhbsiBgO6ucuyjpBtQG0V74tqnWDrP2Acneyx0m6NqYMYmhmWXUelynEIYyoY
oSysquH3B/gcAMMcXBcrfGQnZrROK86zUC+3LxfpR8Gv6xagTzKtY+fHrPYeX5SmNSjucrveNHkG
uGn28dXpF/PqCig4HuEta9aESzK2e3jbGQlGgNlo/PXCR6xQEfg7a98a+0wtFBHUlzOhVY26dcI9
7JE7nPNML1jZGS4oMCQYEj2DGerMyNdcRxcDIKdHc4xI3i6CAZDKOjDTcyFXerVmLDbhvNCW7fi7
MBUea4yi1umIzl0C+h3HsAA3ydsMAHLixcZ/DoOEjbxJI9F5EybbcB4DdY+lvdPQKgiogdtW6py8
FUbAU6TXpsuGPEd3kfySqbXiOmFqUfuqc78+x1BminznPOo+8+5p3732a/v/21VOJxBvSgSXmupT
n7Gh9/iimHDDvQaiEcFSbuFGaLV7PTeb5x1FCn+fiKGL6DeCbbtJwIDpd0xNTNCmJVlQ75Wcs9kE
U0wDTucZ0xh6AtYuSjSxnNySsXpUnZeZzu/9NLHhc05M00bO3opEcsqEmu2U8msXM/3QJBuJbdK3
m+mKZjux6H2CY0s0k5D0176Hc0pKUTOQ056c2jvd527F89BVxqA1OZ63owgjOyQpaGzPZrCoUvyh
BZwrkzdd+2ut4SFBsTkrwjHQ1E3Z8xL7N02gQ1b6nS7+Qga4SX1loaZ3EkkS7ItkWPlOToILc4fw
hHc+sLHOdecR0Z0xf7hDesxYmqtb1Gh1sgHeUEUcDYtBzFNMtatmLKuJ0ynpwFW5YVBcg3egSo21
EXIbNv8njxUy7R5ZcOKjjBqlTpeZxis2AvZKrG/ZWAOqyhLel2UmA2dv5AZrJLVwtU5MIpHDAlg6
CqpBEU6qUHsJjFYt8S3q7b7jgTyrGHFVx93VsdUTV30wMFGoqCyoAaEtxUi8DUC0jc4ipQ8/TEZR
xuZnWtQLL+Hpq77+Gw0/u3nFcuy0SsLTCZq20s9vIaos9UVnOjobkGo577Sz++YBXU5uxE4XS+ii
IQHCcC/jjhw3B6JJ1JLHvprZXIR4r+pYRIzGkJj61yc3nWi0qUpgT9Cvqq0ImZy2SknLVasmT9fR
zN24kY/InN4L5RWleLXaZ59iBT/ssr39XZAejjbtpYMZS2rHmP6mlgJcGD6szmDrbdH+BDMcgvv+
0GQ1a7OsQAgYV9h+QcFgufP2iWJxKb9TfxqQU1MRP5RCH/bpNiY+dlTSclKp0xSSIKvsjLWXqFdl
BuncRfkfs76vHAJArUlt0Vkr2lDZqCkF74xPR+AhT1tL0oBCVfGrF09SFL82MZGEZ5RKIwMfAHgX
eEhtgC/42qYOYQG3dSDZUMc4YOzDTp5Ruwv21F+ZyASkA3L5IUDe6VkpH5OZh9j6abnUy0bKPh6n
rNdkR3mngG5p+Uudufbbbfo0sz+O5gaUMwULn5OIYzSrQGdnbJToAtvj0G36UCzQipRr9P5C6CSx
0xe2aRMiTdh9vFWUnqlaxK7/7VTm9ETXctppBJVhcKWHBtfZ03+McgAuD8/4w2KYLd8ZNtHdyi8w
p/8OIEii5GCZuD1Lg0gdCblfu78fasR3tKQ0itHtFtpcBU8s7IIth1eplaXVWzBsXjfGoTjj+jNl
TLpakba92sz0HjVcy+ennjDS6S4j2JWjZXO1nrS5OtbBdOICgFrksXGsYUhyYxpsPA8d364oV72C
zei4oDLtw7Ih/o+t0qiAgLTvNEbnD3QLVRiepJReZzxOp5AXx43bLUF57LtqGsuoZCh8WrGHvFM0
YowScP+ntDxrCnvGFndZUcIxXkn8lG03QTxswygJbbE2rMlbBq/b7zErTWHS3ot1dHUYCACAEPBM
D1Co6ndYQE62KH+YfgFs+yFs34dNHd1ztmZbcMN3+LXkPvNEoVvNUG86rtG0ydP/Q7Ci0t2Eonjt
JdoBwADxFVkTWs42Kh+I/HcKJr2J2nLFffK+3LrV39TeRBPumucRBsYJe+u3Rsg+EZccfCUcoGsF
ig6ORIdlq15uabA0bazKuSsmODKPo/rRn/Hqz9INF+CHZDvPNcWswpUHTv9wfubCHxg48Jv9B0sE
oOSmLtdGsUo+nEFnQcCi7gQ9N1MiIEKc5RuTj72yaX9lxNzZDN/ZRmIbaFuEr3KSW11pRodapaR1
IIY2lOOsfugAz07ojhc6m1flrNN+oNEcCfFdNxL9jT5N+mhAaRlNAvB4GbXzpzqWXyiizQt3SH1O
0psU3fDn0x/uyyQBciyfWtAwTv/dT4BMTvlrUbNoa39tL/m9xwAnLDL3yqGyV0JLmK/ShAFZofJ2
D4hbGGKshBJw7LQxgbcxQAejZ1+j4CC4wXaesbKI0ibCm5IVTBOxwg+rOLLV8kwgBouW9IIUzIcW
Ghrenj1mcsBK3wHvvctL3x80UeYsEn2ZMCt7UAPVjbEroaj1DV+33T369/X1Ti9Ci3bQShsP2kup
+Swg8kbKr3CR95PypOk4IUaRvxUZzD8lxGIEsAP5dpOlLM2gUnlNlH/qOaCI1Xwq15mBBrLT+LkC
mRNpJi/TepVraVX8RE09obOnhEn1WeEmRnnUgNh7ZIx0KjIJTCJ9QL4Krbf+VzWD+Z12mGMrU1tz
c7JceCjU5xOmI9k8npz+eyv8ze+Qxt22xj1xwOSUCJ+LUT30brTh9TyNNIthQka+bMd/jJiQOQyZ
ScNS/NxS15uZKd1rRYrln9zUo/GDfi0/fyC89TuPkFJjG712aXifTntFOyk0QCO+NCsTzP0fIxXI
3uzH9CgCRl9ZQ6rxKOhaJKpwIl2fTa+h8wRsh53zyBZukaVefQnjB9z57Q6y+Iv2h9eDjpgCZv2k
+RgsgcbYyqiGbdaa3D/Z9COM5o2ZA8XFuc2gRXFTACmfkfvr0E88mSGdGJt0cOU6tOboB39cqDPw
maOCLdst6IOqyDnTo8EbDu+OYha4/P7ThcpAw5Y6EE/qOLGAurGUzfhoMmcjiyz/VMrk4Vp2OIEs
5pXAOwcEWfocTC/BOQZyDgxvzhG5VNgnevaQkhzXx2aEtKASKS62fGSzBz7dpDWtrGF+qcQo0NxI
dxzTt/pRnbsHi3t/IWdUECCj0sZ0qM2E8hJ6JTkyjX2ihY/7hZc9pk/QdBfDL54PIyzoSiMLpKB5
3eiZICaadhp3tWvcss8F71fiL96KsRpP2MvNX0x5WOr0XdTQGN2hm4t3sBVprMu0bRLc+HVLaw98
gjHrb3ue/e9Yl0eW3BktR7g8Q67GBir/Qkqwv3QCoA6uo5R8DdG/UT9/VkJCmgaz/haDhTI3xJV1
7YnKhfDxc708+apzijlG6hDoMGz4p5Vx+0fueZ5v8zM3BIg2QOTxZQxF6n51WwLeuE5fFRjLCMWc
gghdth8Zo8McFNZ2fuGzjV7vTOrG2vgZUiahy4GV6UP+Z0Wy52QIXbxYeiS0BHJiE0d6qeACb+by
kfe9hH/JDsYpv50RhRwr3aTlfK0+lW8eFhBx6mj6TCojD6lRvfO3brve09VRSOXHZSM5oYXvMuNS
VD9M+xKOERJ+lo/IVh8H40Zb66QZnIZ3ITufSXdwHQMFuyAEfWerOjyZpdy1P4fz1jzQt5nJqIP0
WbdaEPLsmq1ZJt7EASw3Uy3+KhVSuELbbpYzZwwhmbUyGU12MrXRb0LmY/0KOYRKjgLX6y1IXpS5
VOxerttxrQJA8HSTbun1MspwY2QuFhcFCV/YwxbeSTaptr93f1mRB0vHI9KUJZf0Pyvg7nZg8NgA
m7dbe1wuU1usiCwCnVlVuE6CUUtzAKtq4EBdWWssaqk7w1UVe6O3kEKnlbmgQJN+2b0AT3zwG356
2dy9S+y/cYVIs1BgVb92NAmfpCra3hSypzTw4RPd71jaOGgTHQRmDPUFtEFe+i0nOxQHpZfJ7ZwM
a5Q0HWzbGTDk4aL3xSFjyvVT/SHZImaRn/IzgHVtwuWzhElui1jDOkWgOwJb5xAi+RXIBO2T8ukr
6VYCZLcZmTOPfMrTlsoW1OT28EPXtpcb6sVJGuOUuHvA6grTMuYuua9zSemQT7GwomCAcnP7y0NM
vqq6mpf+OafvtYr74HhOQHK6frTImPOVoGjdjKPf9+jb2gNcdG+hFIa4zLYg4qOxD59iHGcIjQmX
IUPCvg+D2UEzhJlQ70EduExZqybWxf7xDNWFwZ/CqnpDXG5aj7H0nkC/vAbIs55EuJaBUP8mQABZ
5zai5a6xEY/Egdl0RfFvPfIeLR3wXtAVEtImWhX2v8U9gaAfq6Ftlcj3+b4xJxJBGwsSK0H8oGL8
FrdJVprLEcPLRScSvhYSj/lRUrjjOMznR07Pv5T4FaF9Fq3uR66K5Ak6waBqDLsVYRKFa5qgmiwB
J4AnfI8a81EK9VpB8tmFsQWUOBZcDwV4/AJ5pUjOqgK1Q8rTVuuBCL10nYqpcBafyKSEmgbiz4qI
q4cT3AWVmkmaSUr09Z7nwhqi5P11fhmy2FAnrRwL/b5DalvS9+XvLNGOeVOgEnZHmgnwYXk2lsGd
Lhw5lMu3l4clMM+ujH4gZIh0PB1wTdTNHZEVUCU3D+Prjxz4cHWsZ+U2Crfhp+vxV7RpNupDJ2WD
JdqA9Sa92+4sG/0A3b+qgFH084/+9ty2wBi/AOhATCj7sricYT/Ab2QronbXcrRjWZIgrE3DVbgC
pYtMaqN6aAqpdB3bORmebZmmMwWcSWE76JzoRmy5JvFvCNTQU/0FzyG8l9tSkJCY2OeXUBXPrqVM
aWe8pgTCiqvDCRcMz1WPsmRJkowdicizJMfcvgws35aFnvM2CFVrMkIn8bU0hOHv5f2+ILmyGV1S
l6ugbZUahOAXu5p78PnsDZhl9SoiWri22fM8kbgPoJwumkpFaB/Sdhz7Plr19N9yqAJHADF4S5SB
t9DnsIwgn6Cj9k0zQQn/M/7ESP8++YLK5Wfmj5HlRVGk0Gv8gZQkTKB281bsAVv4B1rG+K7bIBiX
9RbX9fZRVBwJ7dPzUQCYHiD4EChKkNUf8EgIYMWaSgqfEba513VBca6xkknXUsR7SkpT4mw5Yds9
P/XcGC1Z6KRCHTB46ysWBs+g42Hx78WU5iqjIlhs56lEGvG/bTeI1LIxmatIiAET5yF703Kwyebx
MWIESAcowzj3Jkg8M6/sRzuaiwRshPi7hBVcFY8iR7ByvUsi1kKiiPkfpJKEi+q3mbP5yiu9Ptuc
6o5lfUG7FS1dNdOihUIC1lNJvbpnIJgMZfrKSiSekizrs5QaQFDPWi4gNOCDBU/QGOZwILDbHNUZ
XSJkPBVU1FU1d1Wr258uVEGgx7uExm0C8a6DCV9jY2PTKrFj9XYFAg/5SKivd8zDVDcL1aFWR+Rc
aAoKTQY8dsf+N1DRnF3h+lLuvZ9NR4cqpcJZanuq1avOcHAunBjxRjKiV4/WsIoaj5/BQekmkqbf
LeNe3XlTVZBfiNkiBKFGbL8jiRjovndpu+jWv81CWpp0xAVvJ3CC0mYQvZlt2M8ZlhoDMkHP4ARR
LVZkZn1vEXiLXl9aOv3W2dFoncAqA7VV3zBgutBCuc8GBe8zj/Xi539tLhoTv9pxqPTST9NvfGJF
xvVF+dR3Y1ERofZJtWMTflambhP87nP3z5370rr0znKIbAhop/EQlCqEf5KlnSuYgNxksBjZugVD
WJfr1nsKdG0u9/V/e8fGY9hwGEJmsneNlRzo2g0b7jUWo43cmLfvA0t/Fx6rljmH5ZfFbjWA1K7m
GfAR8fhyhMXpzrpZ8Vsn7hHHjumcnUAGF+YCR9rMJ11MTgDOho0aw1O2bL753/O/ksx9s4i7paUu
Ws+gFjUZcTMYl6EtFV+VTIuAhf9OsUe3+lEd+FOCRDiJTjJ2QXjnNYAKZYhBuVrrrTE61TcFZHJi
/L7UXyFzYuPZbeCLPaE0nvIJ/scUBBsAie85MEL2Qop1FEy0TQZ6Ov4+b6CCHmwFyL3yVwZVurPe
aeYBa76q+JlHIsvJEJpK9dMnUkHfYtSIF4sPoaKgyUXvAQQoFwin9jTNXZ0fXEORvJJpMEimcJ+/
idHXZpsX3Bh5phr+CQZUAyE81LCH707Z5vHwoEQhEBPA5sThw3hczAZ9OeAQLgK7IayCkOQT2AUS
u0plqbsetuE22K8cZDqugm4H/CzXIc3qNg/n8XbVvKcXkVxDU7w2dJvgK94p9oO/fenZ0ctNK0Sv
8uXHZ89+3eDI6oLTqT7CujnP6kWLua/pcqKPCTR1b5wK8HBzSKpRQmXAGmwVuYZ8ITr75ZI/d7tX
H6YzcFIcc27vhsEbMESTa6kl2a9mvDAT2w2yXZ/kAqkEjXQAP6F7jCB2Jq0QiUHhfUH9iVSuuXbC
gB5i1kDd1wNBGwpCqtftCLQOaDwujdPfTWIcNxIxrIqLNFyFE6pnPECn8vDsUXitPzX724V1tjxM
GW9iUcWx53cXXnj5mzVxEyM7O6fH88LCStWWGfVIXBtmn9zsS/Y7hCdHNv4vJ5toalqnsnTZWrxt
EoZ6DNdPFd31zdnmjYTXswnDTm31s8TcfzeJ35bWdnKDqFBC50MGywtAm7nbfiV5hwc6UaDnTIwb
e12LnElBVxLTzKrUXzlkqna8Ph9R8C4aSfnHPcGbhLeSYsUkqUlhWlDRvmLZyNuh0iYb98ugBh8q
JnIdHC8BEACDAjsiEPuu274zKp2qnSoMnaPC5tVo5z9T8KSRysQgYsLkNj6hHcFJfJtxY4MQMjNH
pMCj+9YTDr6i7eKNfMzUwpmsy1okcl/oDje9Z3erUeZjcvaV64wNAvlQ9tnKjRh+r93ewdV0s0mF
8mvKNwz5QMxd8HPQ0HQ0Of79CMTarsD4Vax75gfjkYXXvNrcDeg39Gq7GafRQVm0cdZfxLH5EBeY
LYc0eXaMcY4mzK4x7M+bip1xsj+3UIiH9uhjD/QEL0nYZ2rI7L8Y7XSBaPuWlV1UuRh4qc9UFGQW
JdmsaO3uiiyqpcR5g+UcLvo4QXAP735R1Noy8Kb6+pamQQCeL3CT+blTjimuf9it1aj/DuNCfM/L
fFFQVt4qNqK5FfY/wT4BzXOQr/eEIeirbPDV+VNrZAozcm3BULnAGKlhTpAZNkzdHERmSquMjEnW
z7eQyJjSt/tGPv24cbGeesix0p6CdnRFBvDcFfqGFx4c9P2hAFveMAJncKCsLXKN/335zOPL6ndZ
t5ulY+jyF6JsxdT0aPGevocQZJpqz9Bi0o7WHkBZ8L6FzHLVvkN0lMTH5ZOsTQ9bUldtxkUpAvny
WVqTORt01HcSqKwb3P3wKT2MBUV5tuOKmVykzeU5N99l3CXi6xRMy/VCMytXU5OBGv2F3VB5USXh
cG+PuR4w5elcS3V3BsleuThaN25UBDGs5fiOnHWMgvufdCOEzqS8CNYqtTjV1bFmTdKU9hA/qd5q
OggNuMx+cnaTlCHLBAA0B1hBejIwP/1TGUwash9YB5PzNHyRmc0wuPDcjFapM8jW/oDBcg98vkph
uefxjU6zSItAXgyMenCcnQTaCEjNbcACQj0+zItlmbbA/sk3cnIS2UQddSxt/PxkE+sk2zfzYNJg
adK22B7lWV6VqCJMsTMSASoBFHtQka8NjwH6cVAuvgL+3QaH71h4HDufXNJzjgrbwwPuVU4umEy2
GTA2X1NR5NUAkP+bgzyfgEaBkcd2mm2t7vN8Q/lyDQoKiQVpr6Ch50oQqzdxEW+K8v18KxwkOjI1
U32+6GmaWHInyHH3zTbSsg1f9J/8ilZABcr+yt8B9I95Y/V3JcD3hFF19SsaeGS33G9EL/Em8GGw
i2Axl5fHywv9Kqp7tBYM+jplRI0BCUuffrnnM5zF0uxPiaOgkPk0sxHWbg38/jvVE2T91EkxoYJA
mkck9f5Pwinq2h/wkDQ0AF9PTjIC3LJo01qd6+PDoq9sm/5+jrkGmmbmp/EPVamLWsoVX/VRXlGH
dKyh6KmLLMUEFEfo5oewb+Bhxw3ATxClxYMDjc8BwvukX3qvHQroU+QOKcDpk4mP8lHN29m0SBq4
jHLUASmEk7IVF5Oa55vVQ8VyA6nI7Z0nvH1lTeCx50pKgKoKmyYeHxcPiKXzEEFZhhOrrO04iONC
vH5Vf+lIdiHh6s9m4Ni7rRmomhLq6vQbOSVPrpGQOl2m4ADmV8+YXRnkC/JFHjG0A/wLdwtiqQY3
LWp55gyeNzc1ss0TlVpGtWZbUPEg73ePrjhGESTabhqeaE8+ceTJSIlioHRRF0Pd9X/2Eg16sEds
ochaDrPP+qsizMcnosfHJtjzG2bCFtwUPT+Oc047lLOXQCI1s+rCFqoZ9Hv4fYAoMbxv+aPFAC6b
Ftl1eegouWbq58Y3J0xNorM3XGl97bX3tdeP0lwizgNHofsX0V3PTo19+ZCet8F6ZIZBP9ruPJ4s
grSNKPAeHwop9+FynoC2VcOjJx3725xCgxR4DIlv3SCkfXyvAlc6P3Rrs88H/T3/gVDxmfh2mFlj
nsEIzZy6RPQSKtdMyfIXKhPZuW6sOdlDYAJvfvLLvVm7KhqqT1qvPrUU6jKJMs0PDciVt8tEb9qd
nKZxyD/fI3DTUNBOGK79N0TBOVQBqk3ndgQA0xzCdJeka66bsgKFekw+HeC5IIdtYwT0hok51FgG
OSvOOxcz7M7lE64UVBvJFG+JakcEzBaDX1BH5Yl+10v59jOWSjHN17YgKovXkMmmyCNi7614I+Px
KNBhk3GypOKAxrhAgvEP7pvTtDngb4c8Xo37xyiYFe3e9Z/+oYLl2PmRXNMPibESUUym/HaXL66t
YorQ82acreMauXxOtgyCGsI01O644caDcCzuM5gSCIHz+s5OrriYWZb6WE7YqUcpAGDoeyU5V/FJ
BfiTr5Urwssizy9oxNe9XL8nyz9kWfT7KJPJONbQgVDyhweofMQa0mAzuG81HCnjsUvSyTtB0MVJ
8fxmC+NVV1oVB+qyoZ3u0qIhagUjbee/MpiTjQovEJU0BQlazAt6ao1ApubePkO3IGo/e3L8VuwT
b4nih5ZZSml5nD/IItemRB/gF1OLm/dGOcqbSROEvVAWou5/rHiBnoOZKRaDPdIPGUlb5uSC3Eqe
J9A7jd3nL5TmPOMKvPtqeXi1DpLfMJycGdoM65YTcn/g22qc/RG1KBx0f8ShBdjvpoLtE/DNge4s
I7jZpefAwpJP8oj3VQ68pb0efJuB1s2QwktHxCXUejeEARAHO02BZEItszZvZPDsIibER28gbAL5
dLWRh8bn1Hjk0u1tIVw97XfukRr5ITBx+yf4SeTm7I+a5H4WNf21Q1QvK0eK1gn6yrxiYOvzxX+J
Svr0OJxuVMsLKPDO5hHpwR+RnBEYrKnhexWs88r7Y2ir61qnuZJ33cFhbovelMf+kXKMjQ2vOw/d
grqdV72tnL6YfIunNW0eLWYUG/j0rOL4zRp4baill4m1pVGCs5qUR4bunRN/kDNpIpGuivPeXFmH
JQH93urE6cBF2Re3OPdrh5aq643KvcZ4eA/+p3jtMVC001gdYgo6h1EGDg+tqOO3ULuZpO6+kYha
sMBwGBYu8jRSkC9Ax4A27uXPQfv6b2mGqQjQNSzYAkMMOvW87udqKCCNj09tix9xBaCqzk6wANcs
QD7ZjBqo1s2s7AR5EGsEE9WWvcxCGxbi5A+6EhwCOjsJ/sDlcYpcAG8BcoYxcDm1A9RKx95rTapc
W2RLSYrkmYEDwI+PLWbwQZwJIzLjC8q3NaqYzsQEMFeyeTgl1qgDL5skVZ5YmCf/7jca9FwRDpQR
YTWVXOQutO69SEHwbYdwAn3Nn0kO/fUnBKWbcUrSt+Lscxw1BFe4wlIl+Vb+YU5aKDxxEGNksGlQ
HMishbyqCnbBCGsFS/7VAAZb0bhn+tJDFrNUx0j0ewoeLcIRCCwstV7ttaOpA4qg5b99UatfMxv+
754dC/gdSrezDvCACHu6MRArBhyKaQ8FzWNlPNlMpEwWSq9rGQVZxm5rmHxBSTGvt1ZaD6wc8gLG
9qb6DfB6hMZQkj8eukJh1SrGxgIaJlK382+FPDQCthPCDxWqYyp4V+Jj5N9i9aYP557cJJM+aYBG
1q4FTsL8LJsRjhLMzBrkoCld1WJ0PPCB//lX/od1M6+rqDaJrjh3DtQvojUkR4Vh48x4QgG3e0Ah
py9aUUVVED0wY7L0nYeo7mU1eTrmPxyFXjqM3YHPpjrMJU1NeUdwIFmnQ3f0weCDz2D76y7vywNx
K/foGwd8rJ/549mrWshciA7WqZ+Wz4UsYLgqXTmUG4egXawMZHVLM91nIPWGveuu8HZF4NjbYep4
Nj+AW0RWJ1LF5ODV3BrtT/+T5kRGav7IDz+8zHHmSweZ5PnhHMg9zhDvz8/rQ1woiL8WuaKJP2g/
wiGKjTLB69MObbKKj7vcSanqJaqqHMcEZA9bJANhXtAoMp/8+SmXvyMTV6NSb4S+pQ3BMki/96+d
oi/OcCqGLCxbLsnSHKust0AdIwQs4w+C1qiQICh32KEIdEEXXi6Pi9B1c4GqSSA46fACzrpwBbf/
DRpA1YVI8rRnJE1nD49jy992IBGiJG6II2tj4TEEybbkUsyoHAMrYVwqjbiZAdl1sDQXdlFqzNPr
ujlwmyyptS3U965blSCrbqqShbKJd676vQBP+vBfiFpDiDDJ6FOv+c9hp2s0XjhTjwtY8i9Bgz+J
Bo/pYqZn4TGanYbRLiBmMamOEVsLrDtuDmgMMBGIjp+36amPoN+7b1xPxopmpj2hY3Cv4uXxpJVf
stZRT81oWpMyAbvYzrBmOuiMmEFBRv/yv5flD5Y4h/Zcjc2Jq8sv6FLb3Mii40HWrHK888TI+z1n
Ol4I+8GFJxafsjsEhhHFw7/Ke3KDEqamhFXSwwiwdBNewhJ88/u9y235U6WRxoHmHFJaiuH2B4VH
g0AGHuLRgAx7AP6S2mCeUUBilDameNsY6ovTgZMQsJv864HUZbv9B0mS2qpW8o+Wq8Oj4J9VB1N1
GCXlNjSCIdH9cltx45jfv+hWa3Kvtu/Guy21UWHi1mwUxpuMYFtUcHUZIaJz0+ON9jFs36eXU2xt
WaXoeuhAyVHV+0qEcS0pYTH6qJ/3Iz5S3eu0p0W6qtgLRtwzV0fAjBRSwdxUM37Y0sdNBK/PcXLO
BkGAMvTzDR2ww1lfJRqTEsp+O3QFOihJeKdBwdjnWoCbhGy0FFftpvao0+zBQ+G/ymjXkRxA6IJy
75RtlaDL6wJrQ2Xfl/MaFdv6N1PECZxTTDYvO1GE5cW4Oh2Qwrhn8g7mIY2qB5lsgKCsfTGRvD7L
l3adE5wz8J/HaNPRbVd6V8YaSZPjT4meyjqhQQuX0JN77d+B+CvEBnl98tqjWTDkF+ChY8STEAvt
BpD2lsrxSswJjzOaNQy3L23MgRdWoF0B13i6WshsaMD2OcdfE9nlBbewhOTvnDFbto8XAH/furdg
Bpf/h0ZuPEGwKBXgYRYtASXClqCUff1V/JPVjHaqZHx4cJa2S1KwgapKlxvk5VVJskBNu7CNhfNd
Vw0gMS1bMRrAvSUgNYRwwfctBzBRLEvbxZs9ANTn65FQdgb5KAOsr63M/zBdjr9vH/bg5/cZrqc+
KBGMk5nauh+MrvGH3kMzwQYCiQWmAIRuzxAD5Xjxw9TQC1YUwVU0ywzsprM22HZgNSjAXrIUZI2x
cORzs8+j1i38jR6ebi5U3BJlFM+t80sIP+CG0qib4k0UmDzst8j5+FMdxehR0iUpHe7qDO+2P7Rv
E1Wn468CGAt506dJwYS0+ecqJLx5kRCE30ootsUtKyxikGc/ekeSiWapszfMhDVwZsCZwgjbNmsc
MoTz9BDKstJGwMlZI3hWiBHGvo+vvGEw6O8cYMMg8wQlkyxPxL9Z44VkFDcT4DfnzPY7JofvMMce
NbFLAHDfCTSsJT0to1teF0LhQAWvWDORCS1rKzONAkHcNmfLOjTjbdLi7B2pxxIBEkiI2PNmJzt4
EOzrgUsFOYmyl9KXWtbNkW6qDudfvS1RH9dYnKz3x4LX4IEewl82uvNLDRMtNCkhHNOdG4MQZMJ/
P/KrTysMq2LPL1JtuWU4wut3RNA4Va2b0rsvFWhIX+n216r640K5NVxPN0NAnr+FngKC1H3kq/ef
9+HqLNVRpeJo2qqIbwG6IfQcfwMANlPfQLuxm0ymSQ4GQyM+DMzfrhLx2eyVbEm3p+P/APkqdhaF
hXQN4OKsbjCUvGTGjmmYSXKfZtSBMp+ojsPXMYIEf35Ij8X+9YwNQTtntVEY2ch+nu0AucxNPBH9
lUkknEOTVzo2s8aojO9cydpN84Z+OYbUmE8/w3BrExUvnkK+NYuE0Lg5t1MpCwSaAWy1UcNqlmqI
GD04iU/jMvaIlscYIIfF/V+NJyqL8y3hw++3ApjFNil5xFNWB5rkuGdkrGP3VcvDoW1RJ8jnzk1A
vQg18ja4ca/ELrwgc9VTzXWvxWZm1/M1CmTG2dSR8GwjOlHRW5yZi/Y0pKDp5Mf+HSa0ZjkT1n+Y
S+p9A/oONS7jaNjJ8AeKN37rGo+VH4tFGoSQSDGUd0WXxziw/baWCk0vmtyRsQ2sa5e9/J+umd0h
cHwVl1becUDeOh4jRzGXBKEhyFFj8qNZuZHMqfXBzaHePFe/uPDIQqGMDbDD9IQIsrDE8LMlUypT
7jTJNQXkj8Oo7BntYX1Jxk1Z3zgCBczXKVbaMoqqKfb1H4pqJAk79E11xWtEAyihb8mBxXNtvtRA
a7lIpZSzQ8aOo3BjbzNUdviE+/I8AaTgHL6ApzecBZpFViRNgop9XTFedP8cxzb7dVNHNXrMfrAd
bnsWS96Zu9xBiIAm7IUVVRhycvyPzh8G3Wmw01Ly33oFZ1mkOgbx8ORPvqujDqK2H3A5LMZcaQ3+
J95p7KTQi8C+6w6mt9wvV9ZRKjit6vUIB94k6iGI7eH3sQpbuBmzkDGb5NKNzl/JOoBbi7ePPhxG
AOyvgAmnEv7Tm80XSghl7cfZWkfK7MGHiz/apTnMrjyq1flthcS3AGpIjJXU6sWOdO9RLp0a2gFK
6v4O01e83fAoIu2aXjnSFM4Gism1XSQYuEz1TH0e2BRxQznXyQVvSbSC+TQpqkcIq1KvNXG1S9cw
ktOTjRyx31IaTXoxvOlO1qbrPuJQFmaJpSQfKMUIByUWw6Py9Qcrmj0MkqlCBDDJN6vVonvnwzpF
u/M8wuMBjEI5Rci3F4MvMTeTjp78a06XLqNt6AkLpkjDPqd4jVkOpGKxFxhhEtX6AH4lc6KB7lVt
5nq89rAyV5QV2Ce8mnbkxqa+c+s1tq7K6QnSeAmqRBE3le2odlD5S4DPCtjf3aZmUzswAyaW4TF+
SxdNF1WeWyuF1C9dvgr3FeoRWGhKPQw3Ox+5NHNw1LgfO7hsbsLZZl7cSFHbOIkzo9pl6EDSYArs
Odr5aISMuseIjkAx0FEYxRPof+bUJP2oTXwhBekMtd8Pl4VrXwEKPImyZ94W08/j4de3a+yjnINY
KxEeD6TvIZ0+vcQpyPkGdRVea1a+GKflx0XjY3Gmmv4qC6GLhNZTwQS/n3REgK5nXVHIDIL4D+MC
wl/heu7N994uJb6NE+2htz9Qb73cqpShYrXYvdUpgm00n5h67DDG+tGLl76NaqW/wNZ/iqBxzPE6
kyMPK2J+nk7kBYbM/ouHyTL7oM73MFW5Jzv7EjEZL5IdnU/euZcOFJb0UJ+YKcv01H1qY/MjzOPU
8VOxgiEnJJQC7dS5nxEJJ/psmur5895iWwciaHQDgHo3AhdovwtTLzeUYr8uU95xOYKB/t4O3sBx
3dycfCTCGrFIyR184QC+yPApkUfBnO/rR2yHSdRm3oOFMJT+5qDi1D0ymnULv7Og1u24Bhx6FGEx
sPleOgQ8FX8+3WiYXXhF6emTLFwrTh8AyjztQF7ANMnCB067HG7iC8Lrdi+EzLnpmgqdl2kFUmyX
4gS8MO52dRSiMG7F1aDH8DD+bbWDw/afp0niuu+yubFyzh4t7UkXWE84W/eo0sJLBd4Bz1LSEH0q
Wew9pXVF7FyctTSX1Bu+CwHUdFgb3mVegRVKgLD2ZHupM9g6rvZXDKIU9AxEM50w2AovJRZH3Y0O
m6dtF2+DMph7X9dvKLWV0Sa4hQyoxfD3KY4ntKukB0YB4eqFUPFXWTE67VGVJydz0vQ/pUOeiDLk
nC/nP3hwPPx9QJz3N6F7osRMKjRrEtJvvvEoKJ5bcyXVBatKbbaC/leFUhyEaaUro0WnZaF0EhBZ
owfkFc1HlmTwnicKn+Ykj5r3e75vF77imCtamRY+PWS6i/x/4s1ha7DKov/iPizAWG6p+mYOAKQU
YaVNdxcXbthdv0WbmJSsBAsypnavZWrBGdkiF5/g5Ae9OTLTkGButBaN5YEenZsPdcriaxxBADg3
r9v8iceLv/JYIu7cWy3HhffHOtslDWXpcpco7WfgkMBo3i5xUx8Th+WVkGiGDex6Tn0dv3b1Qpzl
CX6aHdmXIv/x9tiZ6eo/6/L1SdgvXxO2Me+5bco7EvUnS9Ud25aCQDJtuT0V4Yt3GMY2saVZTfxU
YeBABjpmMXAvs0fXAoOxM/O4XQh8UEvMQXKKrIIya7sx45IMroplCAJeMD+xZbUASfA0qlYF2dUy
oZ1jpGmy5KnYMEUoT0EvNYA+lLZolnflTDpfgPW3m6YhXSLmF7i/9t7PjV8uB2QeDefp9xH50sY0
IzC5Ck0zX+8mfnNNopdaxHveKK0IXse9+veIzHywyxmLKkM6ENoOt48ATAPB/g61Zu0yYQM4Wy1L
J6VDkFycxoxV2VO2I8jOLSrm7ebctMEs+coWnCYYu3qtrpp/dQT0jmNdviCXB4Bu1OwJzdet3lmN
E//Q8+HIpOpykmoJsJOk0qgVSGYO1VZLYVHVKGdStVyBk6MgPVPEy6kVbJQ7ELzf5+1nDFgoqpIJ
L0prLP+Vr/q+ZesAPyDi+/Y7RheQFc3ilfrdJpTmJ+9C1SpBRhCP9qFig08o7JMVUt/6tBPA4Oiw
3i/Y4gDukiONE111rdHDld1wFdBcKXIyNn7npyNZpNz3cvnp9lSJnFkyk2cZq+uTjc47S+8BgXsG
JHUMp7PXYYQOQMWjB6wW1s2FwnmZ91d7Uch6VR+R6EiuND2Txdq++u3QNfOAxVwis94C03AqAuw5
LC1FLhD51NfEL4GN/2wBHiRcxl8/wlAiSrWRnOjoCwL8pzTeYuYMmAWisydBz5wB9ZYtKrptgWq+
dVbgIcOBM8r9aO7zTsk+azs2qjJsQctcrG/aDRwam9E6bDe5340pGLcQ1JEYmWuYYmx8G0Au4onS
/w3ns+PQJUBWw6aoE+GMjwz50fmqS02ss4mAunovyOSGcoJLpkqOO6q9IOG3wntKgAenaw1xdsUM
2mPjOiAOIhi30mPUi4bP4vTYWOybtoeAFuQ8mMMLqNTT3bcV6xYXiR4rBFsLF/V7icPfQWiIIQYw
kL1LeVCmfba+mV31hHi4Q6rLHB0bFreeyEgwIiLbQ8ORPXemzwAJAjql+JT9afOvPMMjaneL23jD
ypvV6zqWgrKf0XnARpFXSWAOXTE3Rm0Ch/5xOm981h8qbVcCOIx9Uqb7ze5ntSS9acOQPWqa3I4J
UBjHgOOdaggVkhuta9TcZnnogu6yI2t0/PaP+13zPTbDnwhax8e9IgdhvmUy1rb1jjUcmB6KFTN2
44POoTBHspwl2N99MuK2jomC1mOqu4wKhQTb2JaoHUKP1/+/dx/0q9qlnJCKw0iNAzlFeSoXIHn0
L54o9gzAoRT68PBJ1RBqdclkkzjahRCtDfpSHQ9LJ4HdiTXR8yWUnzl6PR89s4ziTdcDHjNv82Iw
O152QbUKWXeg918ZQuMYB+lxKZ/b0Mpjq/DN4040i6VEhw2GW25CXl4g/pFDjgZmlTVAS5k1h1MZ
X1KxR9bMJGlOmTGZqkgmJIcVz2THLjpRur3GyoX5k49kvjgBledk1+BTDHMWhrgCC0m5fg7Cv5Wy
+YefEbov2pHwyb/mwaz1onBCy01xzEs2zwTyGS7nnON+kR00sTzkMjfel2X4n1rvv02wUlvOPFbP
EKPRLDpyWamFKJ0xYsNBuIZrqAr6vKZp+rfVIU8YovInlVEZUnm2BIJ7mEuD3cBiVzFRVP2y+XEb
jYP8edvBTx7C+GGXZ64rCtuOqfp5eIajYBLtDXPbEhBYzaZAlNs/Xidu8Sm7nYWa1CF1bsbTeYXu
8aHAzDwBWQkGmn5aX6GHi3hVLJlL5ntLNTNErpNX4c3YWzEUA4qrhekbQSXD77n2qS+orciTJ1wn
5j/ent5yOTc7XClKlFMbpwhXyv9ME7OqMTtdBVZrT/lwo/ho5wB6C22hFGqbVXkhXDDXJ16pT2+K
b1zz3YJmcKvLM2eSB/RGuH0xuP4ndyAohUBq12565wr7GpEeuei0NtYFDOkGrGI2AHRIGvfFUEmF
j3PzwCHuyX2fY740neJH+SUHiI5lvYj2f6aHQTSw1mvbSNaSjiLoapYopm7HINHBswGOySrYszW2
TZOMLGcwBid9ZJ8KHoyiBKN56erKPK5bZSkm7gQWgNvs4+S5dRylI8c3/RcsNGJDkWJ2BEpm7ayG
amqWsF4rLKI+3IF+pYNYKbUQUCJPMrkgbLxEcztojdeWiXV84DZ8xA4qOoJWx3pPJoIt7zp4r9iX
kViBap8+9gg7u82craYxoqG28Fc37U2LY8UzyQpct+oWFATZBW4cWqz//7OLT98ClToUOpKbkaec
gK3OLcjQphsOkihHZe+VpUV16tz+hIZWpGw8jNiB9sGd/4G+Br1CpNal2s5sK97YS3kctEqAYL2F
E9hD1/STUZWdZjDbeRg+AaOvDTpU55OxySQEJbmiuXY6dNtSYmrWoRUEhLrt/H8zqi3WG+MO7WUs
N/iiJ8PQNYcvzaN6Xy+qGQwOEvOHbg89ZcxmGkjP1E7ycFSf+vAfLItwFPUjIOrMpOB91b01hwiS
MZ3MHNWA0C1e+bR1HFC1lI7SqUTP6aUXsoIR/QCX+sd11C6yHfcyoXJnDpV7s9PN8fqi8rh7H8Dr
aP6QPmYsvZJOaSYN8yLPRmvhT85mhlXbyxMObw02eQ9iXkIaZvxBzeyAYUlj7AmAnrUdaR8ydJ76
zfAA68nmfzSsVJRdV2OjaRrBJp2Hj0cZEcv6O4omszFyFF7mJiIFcbBjcKGYKRgworedQGqTwKCh
8ZlnImdxHZYEm69TRhIweVhKKIoyZtg/z+uIvECIqawZl9goM8NzSg9Ukmxn7EdGLEZ5Xzo0BgoB
XaL1lRzZbymMkZxhqrg7mTXKkkizf8EDE9jEaRcFht57oI34XKI5DSvHBral3BeRf/K19kQgtA9g
Ab4I/xGhBtnASC2UE79lBuC49AEHQnLrfNqiDRKNpxRFGyo3yww8rQZKXNUNcj+9eBIDCuypxlNY
5YQV6hIW+Q/SLEnAmXeyuj73ZkqGxW2cJUbSenhIBLRDGuQY55CGLfQzsUd8VWT2Cq0Ga8ip+rQG
+i0N0vwMCMFp6mWEU/aJrKEx2FqLEKI2pupLEF1kUl0gGWTUxwoWWs+R1VW3xrH0GR/ZyEv0koxk
u8jHigHQ3wpGKabPmH+zYiDfo36JaIARi8VTrxfyRaAhsa5btQWvoK7dJ6z8JvOjx/56AqGBUvh/
G3AiMQvF8gB9DzdJ8xMuL2TXyIHC676Sg9fQ0BrYb/yNv+j8P2etI/QG0FUn8LkjbjTzcJxTerEC
ZD2MwyjSeLNWv5Z17I5VjLXHXf+TfzaxriE+dqS4KBye2iAhnPMnoqKLAEe//6OHjcLgD8KOSNTr
TukVjk2EHAYropskuAf9poUCR2y9aDX6PeeOmGoeK+V3YXt88mF4ZuF97sKq61hMgKcoNoTbP4PJ
utD4s3cUwQ2xzYYkYQoPhx5gkM9h2ImA9X8yPon38LNkUI2hkbwbuEtpPiUmb6QQ4XardSqxLA/U
7cjgnTVuGR5f0NpjwsVXpOS0JNf9/C5gbbsBhvaq8P8baK6CPtSVmWe6uGYShQ98IA48LUWNO41B
bEv+dN65LUUFqh3MVG71gcSSa2naLWG4fB3+PzsGkACdlkSF+jbDX08A7Vz0O1CinedaerHEtzTW
p+I9zJGyuCATeDygu5AigUNhsemBNxYxZvht/FE12rogxbhtGQqD58tLshvYqkiUZNeSi6p0E18/
qgFSaRKZmbQMU7JskYmdZiSYOj041WdyZ3gsVRUNDuV5tl5nysGeXM141SwEoRhf6LVw7BzzZJm+
nDAw7FBS+17ajC/uAl4MYcdeX4qUHfD0MtEZFMIczDKt2izhHXlr+qsRhBiYX/rEkgTuHN+cxw9c
igcXclM4v8/T3FR3q8UALYJ6YzbAcD3/lQ6MiEop1ycyOogfKvyl2Ge51Ol5vcA6MXqt2jt8LSUC
bQILhP5N2YS+vNl7zTwLSgVwqttC+E0KENzaAuH7Bs8i6DFF2YCSaDk8AJ+bD2yr5JnErwDOh+QH
fxF6WmVZjyYYD8ojzuaw8RvCG+0Q3y+sJ8WISshXJJKoj1TVB/NYrOJ9NPl3+Ercjxjo5r3bN2wH
W6Hre0xOmbYF03oDVdRWJvhUuBRqoay+cJbXANQljpAaVEc3raOouni+2ti24+Wwwfdh5Tv6+rth
sQmX7dv/9XBSdC3K0vwVYNe8ietqRpTbnb3ar9E9/7rwDUAlQdjxyZ7UCcGuKtVUgn4Qdws4DBoF
SF41DOa1HOeO7Kj79+J3tr93vu97xS2pJJLc+9yeY+JRhWk4jnx9imSHESHvr+nAKhuYqEffzVfA
3aVc813l9wJF81jqhf9oq38YqCm5vAyMfLO7VjobtSg8iLW8yV8gMv0hp9WPBbfGrJjOzqwE7gC2
r8ltehsCqFs9iY5nxbhcUWXwpwdupzW8xWAZl2rWPuegk/+OUdI/0Z5Y/Y+cRwgjfBQxVzxcC4Rc
ssteO782Un++u4gn9IAWwXjs6WmJLbgs65buj7ToOAvtczFWvUCEjG6VRrOxvi0pECYCNwgvaW6Q
qqpDpB79vdoQmXgkNi9p/ALTyHHwjlruYjTwRB95pOpKq0i29JYEpJ1cP0csvxJbusoY3U1wM7Tg
izySUkenHa8ecrkgoKcD5SvVKweDbzyO36sLjIIiH8KhzwbKrSsNgJlDzQTFzUUD+e4JuSA57Pol
QZOOBrWlW7p4fuc5Z0WkfrTh/WId7V0JG4PYro/fUW153ict+/p1mZsOAzxQiYFNJuHXEPNUwvq6
OXpUIirMl2Bx+f5OKFdEJmxlrdIlkoKoEVYE8QUHokxoWp3TX4I1ITsjc5LIPtN1wN0Atb/FJhrc
F6VoPCo02OhtI4Wqm3dM+GjLP8u9rok7VpEvjHGOX+f11pQdPAzbZPFQAMDBvlhWA3LYywtWeiL1
qM2UuBXNTASMjvaJrjA9K8kMH/KVatDxfBN1bSQIFXDz+LGPHyqyrSCvkglUD2OdyAuMoQXCSuT5
o8L5kob0qmEakJgH+q2sdbfiasxJRg3P1fD7+9q2sVbNEUHXW+V0B6lORCIjbVu0C3onEFwByazk
dcHvcu0Goe3UAWJoa1DWWWFF+jm8QPfV8l2E8q2TGLyyr5jNV1+U0pvk8KbdnPCd7MWLMJetJEWL
K6rgiXcqXUuEInxnLn8Au+DJyeCLF+OfXzSIPPIGKVkD8nbcWPLhmVeUJeIrwdBgbA6xv+TckfXg
53ICVLT37l9yvKPdt+wBjLcsTY199lIL62N6OybXYplD0RQHUDcbPpefvOnNpJ/Q7f05YPfuXT5/
PCZ2/9mIwsTUJi+xmxructedXzc2y8okga39RczurcbBKE102f+rU5u7HBeZDtE78adwyWRd/Su8
KCkLuVQXSyzsb6C9D512nne+9Kv4On0tDjS5DZwlAGDNlD2Oz4EnBWAOOGPF+iR5UztGlSqIdAV+
nigTl0l0iZzepGrRHQmRd0iM9cHYYh/kr0iIAsBwHGoiMYuMmdGLhRBBJ60hKs/Z1gqlQUGidwZG
Jgxdb4acdIotrsRxWlY4P8eWJ8pKmUuJHsz1Ef9xhzW/hN3X0pqG85WgvcAjj6VMYXkbpDxhjZg8
UfWnM0qaVJKxoD10T0kn13XihHH+uhM21iVZ1KVv9RjwRFHJGaCUhxLfWAzrq+yCgx7EtCrh+yv7
dPspepWq0TAm3NRc+AnKztudZ5isOweHEKz9zPJx0xXkzymvLdrdOQ05UvDgTTSLLZMqRwV+2u5g
gvYxb2h6uIXAgD/U9uwpKKulRqFaPg7K8YXylfr/u6nHJ4ZN1ou35Keh3s3A4B4MX76CubBqMh4n
gF78BUYyjYrA1aMR33dSpnUGFkDj5tg2eSLsvGqflD1vTPzAmud/5lCnA+oRqD80OXhZEOehpkrS
Cy85r3XOSPD7mf+r2kb6afHNB7djBUusbjkVHh5FTUhEt1IYnBRPg/sEJcamNTAvxaQnpH2sjAYr
YHmNhXEk5kFkfMGjUyxTGI8jrwQiXmve0vwjFou1THMIBqPnx+qzIeT9JyxyEleGvTRD9LD+f32C
Hy6TvgJYxdZuh7FlnrtGrQNe+Y1sixcfW4iRoq5eDyJQsmbgV5Ejv4waQff20Q+JM6pJ0S/5NBfb
Q75PF0NNIiHwMpAFnYeCLb7T5sSpjNPaF8JKGaqQ2b36G3ZmglEuts8on0qxygvVLvLZJ4nJ10S0
NvckcPaW2/n8xGjsHfn3Pi/OoydZw8wGBkVvsnsLmvPTZ/pItFbbSym3hWWP5wGD/uenrBA+gIvd
FyuIxysmGLrtW2UvIo2bv5Qwp7X49kG2nwx1heFhSAtLvQPaykD4pL6AsGGcoJBrxoMjtNBp6KqS
LUXUqmAfFHxfCKLtw28vP7DC3j53OpIaGSuC7rtZyHU2I7LqCZv/W9+6+5UniEmJ3LvfTyYwfzUa
LgbeoJDXrtg04Sfy93UWk6jC5JhB4rmF3mUeFzbXi9DwG+UGdyOf3whOsfdkaIzqotp1nneN6z4Q
1BMycB1zegbYXl2mJEVjCnxNj5TGHyrTsot6cCq/EkqlVzlNRRu9zi6al90Mvxe1k0ji5TC0Y2x+
oa5jBrjCT05YbBaxl4man2gwrteKnRyilx5Xbk/PWdCtQVEmtq5KdfcO53Rj/59aNuYkz/lWjpyR
UmiyFpEIadmyvGvpO5VmDryeiqvYq2ryuhCR7BWR/AKw8clepnNg5E1q7ppODZfREJOsr0BhBdn3
VyWQBIMUrLpMAQxaIPCpytPIXWHKcK/CP/FUeVWVAhmSdnz5aesI9a4WfK0ngMeAgkISoeftckmK
wZmPhARstzLnPFltV9eua5EcXh3TrSVk6UExP/0TY7paVTSsEPniZoS9IEBZrEW0ancRmwXH6ONs
3exItXHG3xYsWuacvW1cOeOamXbpaipvQPsZJFPUeQGwK0NmLXd9Z+IYnwA6cDUeHP/wIAS0JvMU
RfBQK7FMNxCO1xAs63iemXqLP5PH5mi7eIgHWhvksqD+so91FRMMj4guPhjREdD6crTjbueDTuEe
etYMDCupjjHhiWrna35QdHDlAxJvrXIAvJ+9NqCv+v7wrmDtGp8Ru1lX+TTD9CUeCuoTd44+SJFd
G2HCDTg1m0nzPSqiov4L0Wwqwnos+YxozfS8UPZwiBSWPhBrDhynAGce3jl5rdMjHmZznMjqI1xr
7ww6BjeC/MN+6XA/EMDXOu13ZcmIM0Mib24Iz6M2Alj0dDoJ1K5qxTsARGTVjH6yfVkJBtmqMWri
KkeATyx15MwriK/vVadzn7FgYd1lwOFT6HeCD2kcCwWb7lU5RzZYUlbqacH/X1y/Y5woI4C/vaDF
OicGjHFEc71RkI6fwhThDnwWBEq16Qfkc6FMfnsEzsrf7/X/ylFFKtLH4BbxaZMgZLatPiJHEQaQ
dpYVXe9/mTFxfKvKQWy7jzIR69nnbEy64czgXnMUs3B5Qg1Dm6EKlD6/SgfQkiJbWl55zxQBWfPU
NNgVUJ2erabpIubICJKv0Z/DATXsUZ1k0T7o4zJCXYSrCVfzkleXTrS30t8nET2eVxXFX8Hfmsh3
GgQcvQQ7GFgpBUdtMdkSApIyFhJIJYzQqPYQ6UMJ8V4JCEgYFqAkA8+WPkOAwRh5DZasyRi2ACwK
S5dKt1ARfjroZCJBnPys0k9dkRDbLh4Tzu//ZhvpIWGrNbgmjKGHOvAg7BhLGWJr3vExB5aDM/5c
U1JujcCPXIavEwWqvGQzHK0yC3WVLcsnXQKEARRm4HdMGOuGJHxAfPmylaPAi3LZ5IZPPaXUYq6h
l45ToKfIZ/eH87dFnmwCZyb6l5dCUIY2m1APGZoBxvBdXm171kXNo6LK5ZBFliUxx8Ei24BitvvH
zAqkNYZVu+6UlS9DSa9LkDnBBm9VivQq+K1ktYDEgpJk+mEdl/PpBK8ukmEj/UrplDi31d6X5Dv9
F/Cyl/sn1k/ErsHD1UkUQ4bYQDJyXOzwxD4JwoU5tuFsA0t1/sn98Hkvrbdvg3RtweOF/O3A0jm7
ZbVwFzoMW84rbvleCM9ah+F7g6huCy/LAATyuaEzCrJyKH/iiywKc8ZbOEc04JXvgnQ58Tpy8iEo
iUwAboHbCGetC38U/HvQOFywWmEZuJfjpRUpaNa6IDFZcXsb08k2ltXB/dFy1lLMW+xyaNQCmoYv
b2LjFXoDlF7mP3Qcw+sMWcnfmOv1cD6ifbB+x1Tqu2x1rbfVllQxcJ4e7CHmRbeTQLAo4rmFCESd
VglUqzRTKyLvPcjEBTDNb9pUaSacGCRc7cGTdBKjAMPYg/sowgsu2KsnsQmbvKqYS359jeNU3mox
iOxdLc6vZoc03P31lrvAjXJD3TEbv52mxYeQPRtUou69l4ajknsaQZGX38ZClWejmyxNiVxQF4Ty
m0jgd84TpcygdCqM17UbIh2BvAHnfgG82ANl54WoFrk+Xz2jh3TULfykKtt0YMe0/P+Pl5rTpLMz
C3D8BR7IhyXdbcB658a9PUfQGiqODJjKDCYSZqBhj5Zlc+GiJ1XGUmM5jEJb+XsBZejp3lu/NNjW
EFMkIiSQXqEPmBnYWmatAHcAzQ39+YUG0/PwdmJ4f47UrRH1L1HfA5OOUKiLDQGpNiWeDoiE1F0J
BD/D9tU77y4RPoHoPYWUSTQiypdexuZ+UajdINeq68mNTNZpxiBCo4i85EDl1NPyPmRb+1JbrnjL
tg/VJ7Y8v5YDHUh3Tzj22fRfEgGbGbdzXeYbKfLT2v6nrAp5Edih2BqAXkk6ktjilknWCPnZxGAv
JR2A79FWcDf4ou7ZlJFgf44Lveuh/0bb1p1iJ2snYE/FXDYN3Wx0DSdqaXtS6QIAc3lWfYe/d66y
Gc+GcXI7Z6D4FdMQ/1j0bRatB91c6zuZ+KklSE173s5ByyjVVumqBc6f0UAx4LLwSWGTJH9b0TTD
g55QZR1xZ1YfUmvN7PcUXYZhAOiWyPLa8NpRooFPJYu/KQGtqcsUq00dRsZQdtH89Sdvh1FMbH8R
aXyfRm/iTbD52ah/fjkIMbpTdZdLa44zcm0iinApEDe0ONqe7YEflhoHryADODYaxyXiMOFv6weW
ZcF5vzBf962PB/H7ekU4L+BulTMegP3n0x4bgXuMKn7gyUZe++vOMAw0dG4Tk1tlXzhy7RrbZxqk
cEUbIAwanvIuc3CYYQZYecLtgwXS03PxfiBkgR2G9MWTV43Rn+jgIyb81O5Jh/5sf9nRHumuKMkl
YMuuA1G+/NEJ49J2mJyLmegnGAvSc07Cvc/LEgIQ4XcKx1KzAFQJ84Fa9P4hzhTWvrlAtFv5siej
ysii9o1AQaOYZ94PIH/5LGZjy6tljzvZmAULpyRwdVkUeyPx30xfOf4G+1kil8HFWgl07/7f+v2G
vEYUYHlOaFTUwLBPl7BiY2FlWTz8osFtE8Z7J8+KvqfJ/b0b1Whi5m+orHTW766gjBABh+8/2Nyt
ZS953i/g+tk6j5kExi1fNs52o58qo2vnrbfJO6FSDKXnFF/oIkRqHrxrC5gZ99N4N9SMsDycYLjk
K7pxMP15lLimdM10ZiIJkbI6TrPTNMJyTKEBtgmLA107sL7vRERZNP+OqO2YFVJ6gBkh84Uv4g3p
xw2OqTQwORyvHTRofOhG2GPh0gTadm1a5lcRR5vhDBV15uIjMHQlPDsZTCoKmpTFKkKNByru6HN2
zEhKwb7DEKN0BiXe1nldaF0Qy+Cwu9VlG4VF2RAEMVw0Gsn06hvi1ZdxpS1/vuEjh148/1TcMphl
x5U/SItzMR8FeCHZz30YYOZpf+yfERXU9jhkn/ILBbTUtWKkBy++exZaTC4v7r19BpuyfQSSjLef
4A5PnxDEWw+n8+zRWS6V1ivC712Oae8rL3H3+WnQg8oSwOk7fvNevibwkqiGHJhI+KelKauiRFGI
ii5SRMGR2+AidhDuWcRfPgCB24AhntzEA7Y441MDIVIU7W7nLxhveH3wev0Da375EsEZukTk8Kqw
i28QDAWKkhWBL2eE9454IimMB0V0KgyY1FIQbVeNW+HkxX1Q+A1vF1YypihmoiT8mGhuAWvsqB44
waWKtKEHMHN9AofKvzjPYW6PpBAKPnt7T0/LmuPo7MtqyBNhDZGnohcC5fiE84ba8BaCG2VWuTfU
E+gZZC8ogbTlTXV1Ivg4XH3tlgu/TGKK3LgVSKMDN6p95t3eSHj8wdcmEhoHjkL0k06mZ4TRuZZj
Uyx3GZh7z7IyDrBrKDbKs9iqrV23D8akwwMnDVtvteOtME+vITGhqBa5gatLKEpCba/OLXnL+ie+
FldU8ZxbqL4eGNzu2xv6/udUrMXPsuZ7u3D7lULI9FYxkIm8Q7TekGqA0SqMlzFCdFB1e1mWJ+y0
KBIb+aelektDOtjY5bgITl5/0TJQ/XGxAQ1/fz9qMusgHfzMiqI0MiIBV2S7I98dYdBEGK4XIH2f
qQQ8zZ9mMazXeBIsc4Z2bTu12MFAfgZlYcNhN31VCvABhM4nFHCtTcS3vI1W2+CP15dYFESyV1jQ
2RZ72kseJe8tMLGYIXUyek2fF0rUBrpif+z+F0AsehBUQ0hKHmRZglnzzirgmTw0BpFZLJg4v8wo
vA00yzBSRx8zu3QP4BoX0nj0eROgsvHe6XfJUDWZjV5YBtA3LUkV8JmXtjKZyNcYKfVrRQFnDmMF
YrgYR/3m2KeyGg/v4mQnqJyTLwvSeEDo/8SVO/Le+ZIrgYUx8LWVo6FjFa1Ypi09OZ7nMAZ/Zpzf
aMGyh2epn+8eocVs9aZvjz6KGqklJc+WyaQnaoqsyGQxmPZwCEWDR5JzOjHzha4XIxeQZPjcRSeH
xuP84HVVekF4tEA+t0jdzaClNcwn1bytq5TqjqrooNhOIoSrmmBTlr8nSFycl0k32NUkU2pxzbat
cXeoRO23Fj/uHhOL3U+GEsjq/CAHZZx+UQbMhsDipVHEB5ntlOM5wY0YAGF78xNhoMQ3qJ9EZUCN
OBOvozDs6/HB7/SaIqVWv1GYDubMZgp6bW7DbepCfxxhOxYgtiW4dRgNbIV7qHxRL66Xa78oTe8P
gn9Fzy7swHFcWdqGmluRTDKLIwcYRHAYFzYWSNfEcI8mfZJ4muxg4+N2hvCnPYyTrcr5HvJup3ok
s8zXv6tKcQSQB9RoVl7w0lal+8sKjaLFJfK0u9zMO21FNUEBF4BzXzgG+IU1UL862Br/q4JHSV6Z
7FwLhN4CdXn7tzQ8TAWMmwMMwt+ZAGh/PMu/LnC+wOxUPo0s4Ylahz4qKCwqLJNZk8qrCplf6JBp
uCxzLqeivHpeJaguCThu52Spq9h2szjLAwIr6ahWVgU5EOQ4e6pVnv2mk3Sx4Mouv/tWP/HFHPU4
o4jTAjGtljOkHy7uB3sulFHjBWkag+msHvJzikvNU7GrmlfKI2klEWgjv9BOE3qOV6BH9HMpQCPq
vDhjLuehStN/iYhlX3jr3o06heE//cZrZ8YZL/7iKiaGuKMnzp3PRWdQR93w+DoLZgghm8aCSxsu
Ve6vrfHQub3dVKONsQdTIEXfGqanuh8Y1A5BRhexW/6Ld1DGL6Mv35SHFjq4PbBc2EtIaANwP7iC
RGKXEAvGmfpOlNTbNTuBn0b3KNAPL3fG06r9NKECtoX1pl32u5SRS4gYa7Ddfw2pvKNhHlKqQMaB
fJ4ytph6ny3iVbDBd8d+VM4kPQQmyRTAyCzl2ii+yaE3JKURC0IEpcBKr1kF7kA/kFdRr34MpXGj
z09UhH/7+aQGq9TAH9QFii/JsyLTiE7cHZHP84CX4OTM0KcGPcV+LG1a0/9jA9D5UVj6jAvKB75g
GXRvhqHQrmL7a3LxaXhPJ8LBauLk3EWMzBENOiy7tfQJmUGNTPqRK72g+IHU9z1WICwy8kI++GJ0
TrQ8AYlHznNNC57VPd8sfbH9vQzCSlBuPRyjLkPcBVTroZq+G7u+rxX3ra5b8h5kWM02f98PEnDU
pBHvtSxDMftRWyoaki7mWVcl0mKIUtR146Y1BVIZYquA3GmK8sHPNfO8KHcJB54W64mrWbNqdoB0
vfJ3PaFL/GYSu0mO8w739cAWFwZK1PQpRqtc+1v8Wh8chXreAS5oyPKyQFWoalnZAHxeW/JX67mv
fyaEOYb1ZQAxVyVfUTkMIRECYBWQz6grQ3+wPsFSHD4oRR/OGtyssUCq6FqxMpJ+A3VNQnGE/Gq7
0TpITm6BnCbOcs0d+WJlBj3BfiuSlpbDHhrb+SH6IHPFsTvtAyo7KCR0x1ohK0WgX0NtEFaJLzMu
spv/QLEvXY6JC7o5K1qr3/lESVBIhQrHMRSUnbVWCOQtPAoK65THNwaXfpSOKp5QRkKYIRSRJrEo
1bvKjY3rlGegAxN5F5RDERSBWic1N1eKZTAMs7SfF/UAluDoJ4t+jMOVeYVUVHz09oMaJumFq/L5
Oa1s1gpzY30tPRBTeSBSW/eGGv7Gy8FL7hakBeiNsS3wtYSYCXCTVLzfX0R9yC4CT49tyD74kSSw
Hp9YzC2URG1uzY7UvDOZLDCeitZ3Q0dT9KYrB1Iod8fPPUG7PK4l6CtqXu73ef8CjXmGGrf3lHKB
u9d4w3QNLhs6bV2vPTfNKJpGESJyliNoe6Ybn+da4Oy5EgUSOAxfoxsjLMXr1/rtFtXRodRsRS16
ZUNWvs830xUXySmhO0HdRyR1FDHVqdDbt36LGB8naR8vbYbV3PtbIweOlyZjQZqq58qkS6xsxOTi
eyqHVROnORIBdZ3y+xG4TpfAGzEANX0u9LAA/m5qbixoxOu1ttjRRQP/nE6Uciu/xG+28V7TJdh2
An8Dy9/YineZggNl18U32oe95Ri1P7nf4cX0ipdhuAdut+dQTjixsLqCR23KMz3SY9T9glSf6ZIQ
D7SZuiU7mA8Tk0SZupVfeUCa4Z3RxrXbTR528XLloxmWxHJgVFGQt3IjOXZG+nZ3zBRWe7ZQZR2u
1ASiYz2h8akAfkKdLTDRZuJogJhhN7JYhm1jF1Yu3svIwZh19FwqC4Tbk5rj++p/wZOVYvTmR6Qn
dfr7mhPFb9SFnKtXLxbks39GMrZb5iCo1G6+tUFd8gbALDDioo0L718a4WMJnK4ddULBcIkQtm7B
aLFR5C+sWsa1TIIF7P4cbZo1q8bBdwgT9ZHI0xZ9t5B6u4GWS1CR1R2Wie+UxmD12igaVyDi+dNw
Cnx3l4XbgiEruCi+c20NKf0fRlmjYdcOD6PaxNGo1hT1BEK/IA2tZNGVgEwQtyQqa2DwQU3R+IVI
Ha+nDMjOBXH0B1FjH+jYR15J7hXPncT616RUlqP6WDuIRXvA9Xbt0V10U5GJv4i9gN7emU6/EKkL
i3ViVMVGH+pffL/SLS53T/D1spNx9OmXR5kfE5CwoCeBAuyM5bubDzcMNIAvx499b98Bn0XR4j08
VMrsl259ol0k1YpWv2V5DZ/EexvuGxogzhRXobb+C3aI9uaTueLOqKlDXuJrDK9D2yj32KbyuOin
FNl4hiDpqcz7mEBPF7ru3NoHWZW0RQDKRIk4itGj6HfxSPJ8DcBGTVYmyTm8V3GgaEskfHI4owBI
sSbiawknHvXGCXJmyFzNzTANJyuwgZ8q+mj6vs+OwY2r6UgSFisfY+WQ0ssnPsrM4RZT6U4fokd/
AYTqEpr0xr2K2E3OOT/uaxsA8i6SSYCA/MYSqKevlID4rP9J3NjRX22D/POgzhlYKglJwqZ4cQXP
NYCM9WexFhF0vEAumTy2LJWAhX5kMkipnePblL251XVs0ckj7J3A6DxKY1F+fcaTIK8aTO+I3z9i
G8i8PdFVfJy83fm/eysXsIIf0WscUntThXr8qDBsAfke0pVb2R5pS5gIKOXlzBQ1+JoQ9OWGp9Pj
vf7bcRKL9tdPG1pQKpn3mKztx/Cf3qF7x1FSr1LY56hrWn3Tg/RA8/k/9tzLqxIUYAJ6mfbuVRVI
+IslymQHpuqa1At65BSLuXWNFl+OxEJdMMEci+jJ1dCiKbC4/Ol0cPCPyWuIEzuCfcB6eLpJpT2i
Qavgy2gtGBoN1clBF8Phg/pBFKy49EcL80VSVLFl+4jdTMmfukJRDWwEKgbjxAP8pkC6q5jz+Nmh
N+9iVHnM38Q4fOgJDBlotyfsZLH2wn2YtnGGN4ZfiyqRRBB8zpNCxhbqXcNekQcN6+ksowMKcjP7
amzFq8vlyz7K3l+h2fjEPguO49Tk80fQ51+ml/2yJAaqs6j+DM+NSVBQoWNQzrqdxPLZn3vda3G4
3PTGB/m6lxC2RmFiXvr/AZi9LRRv2tr/JLFfVanWb7thcBYXu7CsTm9BWao8fIp2BMu1Nxh6tF4H
X+fJ4yByYoyZqaiMmCfBTJRkOO9zmVRnc1HO0p75J7r05efLr+8vNW5A39pIHlkmhaUD9w07sYCB
+Qa21sFqEiPthCV2ljBuN9H+UwYdETw3ZrPFB2Wp4wjhzD4243daWb6HyCIk6kCsYKLIoaKgVzf6
pXePMihtpiq4ETNuQrco338i52vwYfR0DatmQzzWqwkn2AGZ9fm+Iu5hslmtQ2jspgeuO3Uc6J/P
WHtq8Ph6v+5hXP/tyAsCuQXpH5MifJdYRrVc7lmaPrd/35anc1ygtAiAjjf5zuJejfV6fnXJHALX
jFe0QLnZ3eXCvTzpVP6LWLSJdcaBAs4h3/g6ReD7UKf3J6ken8bpGno2at15NBaocGMDEnsDSkoS
eLMbEDtbML85W/7hfhcAVvFu6EwHNG7+YZqF783ypzoo9L0wk/XlaeJemM2m/9NOPICrDtWw+goo
qYz1Vlz50jXCGfUuKT8WGZN572XW2s+lJVMXkVUEU0dHoGgCiX1JS1+VpdAB6KTFNYZuc7Yk37y1
9Vg7z21dlaEXDxCeaDAuvHrZbtYGqc8NHWYa+XYsjanWtQSIFn29Z/ymCMVqUcMqFkm/71G2E8Cv
P8GLlk9SfUG7uErmw6j/AZ2rVF7EGSZ4vgJKtfH5nw3O0+Zol1nFN7Csqmp3Calakkf43cw9EgJP
uBQK4camCTScKfqQqBgpvXQ53bwMopXk7axeGZyuorOo193s5wbEM8G4aEBkM7vWc3k4V328bVzm
gH3ZcwaLsx0Q0HHgsGN1ffj1gzefu1+mMgXD1tzMdI6IF5Qkx8bLI7vHf5ApLJbpxjpY/SIxFtbu
/SinIHXCjGKwqTNcH+/ba5Iu9H8qOhu50DBOlzXMdkrbLVGLtVMgctlyG5e1NnoZ57zVCHmuT4dn
XkoEZzJtIU3gE4tpqOWfGI4D9isvs4a85NWxfschcePDTt2BycM2IKOvVaaDDdPKQvmstrwm93DW
2knsopaZZLQibZPDlfF3QjiabNRKfx14/ikkU/9Swz3IZuMp+J6bgx28gRHWho8JBWMCqgSLvumq
WrCup1BWvFTB2RVwnNf3rnaKq9oMRrHYszExeyJa8+1v3NeLFpek9YhTxvrmWKGR3wfa+PhcBNmW
5nHZRObqIFN+SjdwDL8CFWh8Kpd+EKpSbStcNTbfH4rNVApoJ0exob1kFfkHzs+kkona6pg0O9aL
ZwHLisPwh2/a0E2IWhBPxh2w7BZlhXMbkg5Oo/K3jCX8aKDycK/nzfi0x/ThdZ9JJD9khdkZGRd4
HN4q9O+jrYzBzv7YOMH8uwWdMC9slaw3yBSG6acz+BMIIsbZH1euRTCyBJZ9erLLWNZaOPHotBco
U/sjleQ7Oe4xTbrlGSrrpZP7cOi12ywPkEj91HX9noHJ4hrXgRVG2P/fymSER5Ol1g2+s2Cjw2OQ
ZyjJRIrFqzngibauI3y1sGKsi1wxOAmelAWigTHMEqMyuE0CRq+MhYnI4t9Ymrk3BbShaJybeaZW
lhA7wbRo8m5HW8Ymu4m+lIfSpXaDEqvXyXL5tsHmZ0MKddNVQhHKNrqWNYN5DrG3ILey1boJe8iL
6W5eEOaVBjBDoOrzz/qr9Z+gkyMZ2t48BETjQFgzTLG3V+3EBArvXti1fWP2W7L53iGE6r6fSYT/
Nm/gKO1KIuxEA4Iu/Dln/rC6udCsm/XBz1KBhdmcFOyTl1x9p5Ns8SHUZVoOLg4WbrckmWQEK94A
nNYKHuwsvxExPwrKAqLUpCBWHwkGAUjft89dkADz3uFz466jxV6yH4sb6GA95Yb0sHtEfzU+SeVi
/Y3g8s+8BSotuXBKnAlLa1/rWvByKnvOwc6vNbWuGLRINYqYgwDJeqQyIeIW0vSGuJDqNgja2NIF
7YqrD2dGKGk7AWXf5fK1uswhaPufZJyWmuJfPJzjjCLvLTqNcw30RLDSn8EF/slcXiZSaPl1WfNC
X/p3AFRHBK/1z8NCb8kBaxLpCGOWy/MtFuA6yJiNfrFdbqe9ja2jUUEo47+39ep/LA8UCiW8OXwu
NQ11P5WlANL5pAiMcwQIwVvfRuZS9x4NDBaY3Yi24DkOYzTy/q9yq43h4gD5AIIzA25MOXy+49Iu
CRIyC1odSkCtjuQSi+6JnRXRwCfZoifABBJ9CVgsUNlnWIGVFx8jgKdcL8qLan7cWoQ/tDDkbVPU
EDbstde7lLsoxpljV/8jPIBbfWKYA2qYKPHuxet8t3QeKpaUNBkdX0m+kD32NATBz7ysfaEgg4Dd
rloaTj0RpdY/1Lny22cjYbQPDXBgzk2GcQufea6O7nH+4dlTEgEc10xWl4341GefmPbw0YN0Hz5+
O0ffg+VoDD50ssDCgHxvRZU0NhTemFxmAXvDhfvOaA14hVIfw09CGyNnYdXBxh4T0GVrOCsVBHYY
g3Z32GA2/g762Jegyiz8XE8gxm2Jo7GvlGWq2vhYboTnCsmCsymvccSIsyLclE5qK+RLcO7DNMQz
Fi5+3Ywpx/42OqJrLAZopOWKsB0RP1eyBdeyfdNEv6B49adRBHLgBXmIHCsVSY2oqqa+mcEtvRUQ
Hld+iesCAOqM7GlhznCagpFc3gfZjqsxaHfQSbnS4GbrHy50rSmCv/qq3xmJsdXRLlcBJ1Wzpr7C
8Tn5vAAdU20nvV+1BFFNx3VkwTgLbVR4lW7Gwa8+sqTnoy9vgF1B8UvMNjSZ1gd0HDVb6sQI1JYs
zNj4LwLqfLQTGUBp3hD+oh5zVf4vBg+IaBw5SXllncFTYuXKnr6sqFWMHE/o0tEHdXFq1+/3ily3
ju4CSEMYb5EaX4+dkW/5vwGuhyPnq80q8tdbkZHYGmBPZn4YgarFn5tQxwQZ7QbT5BD6NiUyMi/p
3SiJ8Bu45ass/WJjU3Jy5N+DMLV4NPiQdMPh1AKDbwXglZDn1wXkacBgPKx2dqz4n8ByyTYOMJZI
SJbYRoBJUbYKadwhUCh+5SzXNJGQ7oSVYwguQX0XJ1K+fNkLjKmzjg3pJtLPE17+ACLXqbeLMR77
ZDHc3QwPMBQ2mKUuR1RcdCPnUVJ6xdV4fgkCWDH7Hm+y/ArpEEqTx3K7NMGlK047/1vrzqG1b2ve
kvh1wtTyzGKPUP8eYR2ZR3cZrfEUkw0kfszimrO1n0W+TQaP5xLjSWewpjnpgvoehDNzsjYkx/vE
ZaS+7LpMgp7WwqrmsVn+NDsshs6ZzspxPGrM7eyuGd6HJKoGSWBE1DR6z29I224CucJqgK59DZgD
RRD5ItIp7tc1GHNSB4QHdp48MjofQCq72H56NNJ2ACTs2P65aWROibNyDhIVq0aPDzgqCf5Wxd4f
2Oy1i8+lLRVW7tPzJ5m0z3M5w4v0RfO88rVIwRjuzvtodTwdZrz/DL86iKUMqfM+WBlIjLlw/ma6
CcfmPnSRglQoI548Wm/86xJAnt/aEnB0qmGYYQUeavtkNv4BZ/rt6JJOtBH3OJyPs/Kqiadtd1AJ
1G6SLprJqrE8byh4HrJnhpzhEbMw34vbhdVIDnmHDrc6y0xTY/PPIMJne9F8LhyPKg58GWNckeQx
UIuujnJG3E8bpGefiIb6u6M6COBnPezB/XMI37jf7XRlYOqdqiJ5uNh/xVQpx+0fgemhNi1G/ldo
EJBa9x55qYlXoi6CM/fyYP7MIlnpZXshof71zx5AJ17niOJCLPp5ZJTKCjCqlpYAwPND4KQtk+Ki
nxutYqim4CJRJhMeqW1PlE8kMLstOkES6qkELYOradwmWw2gpSV+wKLa8jMUxVRPZ5PWAvJwmKGz
Z9beZ+83nDNJFfRNySjYpUPZLOyxnbdwrHst1XvJPva+NIsW4573xAD6vdeHCTX3Px5UXz74PKix
jBEnZFwyF3jhu/vlBh1mn9dkWUttT3kxKh1QBw4NFNo8Ee7DMIeCh9IsuZ5YipOSouKuOpfojaWv
0VkSGlwumPBZOKxrqIrE2QmxzhOjVgtYB+YnlZr7zAbaWsDNMTnug7sqwF9wg2zUSQ2f82ifo93L
MTVFsnOWEoOwUoRVFEgKuJGeXtXYHHuB99QctUJ4o9iOUuWM9cz6MAjGIfkMBoUiEsd1w0qyTfcl
J4ngqMDSK/YWjrPpfPhzV6gtyGvKda/uIaCO89wVAq0Q5lg0PVk44zq/yWSJ1fOC+4HdZfcskuSN
z+ZyUDWQ0fZAYBRtCutwPY1f4NvPbdJ0N/pqbCF8DcesFO1R9HfSOFogL2f8It5rJPFWdYgE7uKj
tF9vZ/yfPiBsA5GSULFxL2A0a7vhBF/kFwGbNVmSMu9WWOqxG1AyESdrATcCSCBs9sRLEcYvI78i
JRpNb4FwZODU4azpkEvvH5Cjzl4RfCw2l1TgFBt1NXYbmAQqfDK9an/WHpMfuNzQRoxCvhhaL2/p
eOzbw2HHiiigpkTcSDTA8E3pWY0mC127kd5hmJmK7zpHRJBkQuBZpJrQ7XWD3xAs4W7DsGHXIQU7
rHPEdrQWJ5QZW8BdO01rrLWbiJHH6bB5KcbgExQPk8DDW5RjdLe/9wE50d0LtcRMLi0F8CscvyyM
B55hdneqfMFkenVpEyNu6KAF1QUpPk4OLHfhksjXwCYzAysDP4I2Z7T8b8ERhGTDHcoXAjF1GjsS
DWoxutcArA2v7jUOXVnpcO6E4B4rKn6zgispAXqP4Ckrq4Srx/mB5eWjOjFsbuPdRA51fDzmxjZK
44xE71Y0N0j3LvzoB7Ux9g+n6QC8dMKfin5w1ZWTVAvSR5EF0L2pZpA2VSkD7pHrY76Bi6c2SgiN
Q8B3TIn4WXaoBUaJrN6vTVIFtPuzHsQwfe5FJuv5Ob1B3e8EChJOvY2+t8W8mv0NONKTJQX2bVS8
sAHJ/oET8KMBUAceMejdD0otxgKF+7btLUxy+tKxQJH2FwHHUgi64MX6VAQlCQU2jlvKpNPto1lv
NQNqyQQ+sEaA6RivjyEsfuCM9G015JlUxCmrem2n0qCZrMTTdq9CA2QacrH5YJa7AHwt3SkXTPnF
FErinxseNH169ImD/z/CimZM5d+9uY/+kzafSGYQMpnyiuERHg+Jn3b9716PFdHdvxJArD99TFZW
zdLqWXQ0LTCYc9CH7F1tdB3a+GswGtgB89xtUSTarDXaLIkHqCtNjSmNvnrTKF4VvpOwHSscoDhW
6Aqii2c3vo4Aj7tIsNxnt6bEFYD4I58Gtuj9rKd4NjEww+DwAQPm1l40U4mX6EVvNhbiB5yvznp6
rr0ClS+kCyfgKwatYMpwBiYcsQgOjw2s5GfhbOiHVyvxErM0jLSovRaI2nWaxeVO4hsxdrDlZ0Cv
9t2B7W0VHAswrkXpmpmvkC1cpL/p2v4NilytKzRFqM3sFZt5aKRDgtJOkVbQo1/Ra+5nIjfS+i4b
1MqmSvi9XA+Tb7ZNaCHpctASqP6K7elmNkpCrYS9GG1qTYaSOLfnP3q8+/7R93pkz6Hi1KIgGA1M
q/tvmO/9SE8t+WCapfqD1+eSPRxpqWmCr0IZNI4gMcQNFx0XGZwSdnhTOSXZMFGRr/ktf0Wwhlcg
Y2Ii2+w/UOKTTRRpGaGugaOW+EIuwYBn4LieYLHcX/4wE+h6wXqmupC9w1+ypPmPJy+Gj58GJ7zA
EemZoO50LSiDCrUzohpZNsdRhLAwd2RJVc0awSBpb+pEx5JP9evvPVSWa8uSqPk6PErLfGpO1tYO
+xCbya3pfoHNDBxvIP5hzIaRVQQSFOXso37hxOCTecUsNc+Rckkuipc2tqxFjXwlwx8SDa3Fkl8O
krtPQ+yIEnmObS1wnxLH/1K3hNeGSZhbmP/8BuQMZJjL+riUJDbMe0OvbuLB1z1IkuP/gOveb44Q
z67ca1BwuqRNKZAe1/59sVVYDDR6X8+erdPcQaZrgU7XYEtU3HMndARY1inB0iE6IS9UvF9/Fn1Q
jk+uxX3X82NKErJuo+X55SDbFmZ+sECzQQyNJYX2ud8Ezm0KELJLlK/gVaoWLrfigo/G9GyhyYO0
D4CK/5SvBZJWSGiYmHiI1Ro9rC6XhLDe8jO4FQ9wmdWN/4EnUH2oaFuukQtdEHNa4Gaj/EtcJr4C
qX75ABqKsVVBZPKC2cqiTWZUh4gbvx0boHmUfQUpPu74FstpBFs3naX90RZAzrgR18df19tbiXB6
2xVBljvqGVgrjYvg53Hkq6UTxXTS5Tp0p8zVLAhc+YaxGM06UouLfoOWQlCp4eRioaJd/jx2QRO0
OuqJa4ygcVwXQbiWAcl+ipVV9IQMGBY8NOEczcDi15orEsdR+plmBE/JXSrE8TyxAV8Jzb1fIcjN
myrfb315rjlza4HCPU1ry6mV9dlGtQ2Ib9H0sgZK7YA0L/iW/I/ObwQuN2vP8lwChadicLVOmV6s
ywRqRs7cscs+a1TIYJieD+vH6YGzW1VFZRLbOik3XzD1o/pxvir2dSth33NQ7I3Iy22KKoyXCyRD
lNxTdGpKRra6e1sZwJ8yPDDqaMerkkfwmqiEXC5icwyaYDjkfnDvVupt24OuoDg5DZpSPmqca5WY
UmZGH4Uzc6K1IBt4DiahcWJQuzC0HtbHEoyQw8BRO6G9i5SDDslg0M0IWKsnZUxPhMF229nbhnvX
94PntrFF6scHbuMQSHrqPH2JZPCaTge8/xCS/nRu5aXmJbFEv/1uVMf24ZVLKbeyzyf205JDwRp3
7i2RqaT3U473sKFLQrIuG6xJvGZ91R3G9s3u0FFGjTQ1Q4eW0Ftll4ZxyP4K6Yshw03TNkj29ClQ
8Asq4N7Fu/fTHM+S7r+DhWjRmEcg7sVVWuVT0NBdG5PcwNY3vRjz5zkPiEbsyqAdlrRI9McXASr7
tcQrgqFozWDCwXVrR71nyvblJEEaeSSU6oTDJFCx8gSqUebHihNJxyRCQFsGTsqs4gMj/OxxW7xX
S0z7Fow2G9GqD3d7wzG+o4xSO27dDbjxw4+exUIaTJ6UisD63y297gNrBejR8fSDYL8KKWabAbIy
1BjGaj9dOxR6/KEuVIjH98jN9KPrvVO9Yr7x0FyAoqHYTde7/4Z5BDkqpmxh5JZ3D5afe1H6Cfxy
L+TXgP1AkLyljGXJGshZTy3mQN0l3ZYAAMPYrQt+uFjcncUkcoIu8pzXRr1BTV762czSh2wcrTiB
cx6JEQes1PlbQNJvayde89n3b6SBKgmGgHuODP/E0kkiYbMN1yD3OILNTrA64IoXRBh/VDt2ljqd
8V4WActe0NjaAdEgmdPGZlYJfH04jywPRnSFtYpmvqyzjmjkFPWFjUpFcbZ8ayzTVyACey8LQOfy
R6Q3lyJBy6mTp8E8d4sbJTnqC207BYIrB8gE/fs11rLp1cBwI39fQTSuZVgfsKBtx+H2JhWNWa2C
ND2fQ7jowKcVY6SZVJusAdNCms7Zszl94gw97VzBYORxE8h88Iz+b693zI8Dk99f3IdbwfOiMTw6
NHlhHuxBQCt/ixd0IAdRsWJAl7TNWgR4yaPK1jGO5Q1Jh+VaY8VgP4ACouZJpL7FJy5RLyBZtF/K
LHYcb3ICgblsHFg8pAM5cGmZh+2pjNrWzxB4OX5EsPZLsuny3Ex9ZgEoJ0DdK8S4qxT5g+9VcmDf
yNunhGSQ5fuDEPSrZMBURRizbhjcxT00dfUqt1jQeoErk18pGnPjHmaiUIzzCLj5dlehIZMJBTsz
9C01OStfZDa4Jfb2htReBdEG7KiN/DxmhT2KV+DY0MYY5Rjru1yUcurloyAtlG269t3BQGU0Ary0
oraCtjody43a+W8r0sk99f0jSgMDFjgNc4WhZ9BT2ALHGmao5eOxSQWvF3dDWGlhUSmS7qLUiau8
PMFXaJF2Ja0JyNFx5WCfBpyv7KahQ9CFCfY+3f5Al4kYhXFOG90e4sCoGrbc0HLha20M1CEER4Wm
Q8YuDSZk7s+gc1Kgaer7pOsopdOiN8iCZedULEUGT4+NZTX0QzfJz0VncbXad3DrpB5Z4lAtpBLg
POiWxTBx7rNxNQzhbIziebDhsMbbG6DW6raPosHja6JJWjV9oozeM/E5XzzGogcwo5W3CZuaSTZE
/7TI2yiZmptkNJKE86Y9RsAZNRY2+iUXlMI+tKW3MVurzc+95CJksxk1IqGMq0AzLhqRwoYQpQZR
Fl8/esIuX45BqWJIg5tyEYG2dDcywdurW9bcV9P+nUIhpzLVeINYWoY5iIXtf152xzXzumjoYtM1
M6R+pUxZzFpq2Gaam+gVGuRgKXzO7H5T0Mg2zZaqJvoRTjjr854MK3A34M424dwxCXO7KIoCWwJy
1/89qC4nvuZkv0hPCmv4ID/v0S0tr5WBAAO3NQFXbM5AZu1T7ETtSQ2A8ZloufHUd2Av/GLz8lsl
6cPQ/OOW5lg7cBl41smH2lp24As/vzUpqCNtWIy3/D0Xu1lbF62wvuLGa0KowPo+DCnpPjg/ceq5
Fu7mGJ3PuwRFQ69kA9TwT62yQIdmEnMiO57dxxJ0kzXInHsVPG9AdYoeiTQ+qxKPtvm20uCt6/MB
xtXGszRtOKwdzKSBo94rXBlYdeecQBevsg7PLLqfgbp13Bykym3WrqCPEdAevG+UNuIwxavJngnI
3Gox+k5DqRawsiVQGhYUirmdNl+eC5qTkAOC1ORwIXIsk8m3G7Sv/Hi1Xe4Crkd9K6qA7HKWNjGw
dW4nGBR0x7mjIqoj0cNw243tDmEXGviP3lxJz787gikZJgkYBAzxjEzFJsg6k2zmLhaYdyUBslAC
0h60zU65dTcfy5z+LOlIu0lqq2UaHnlDklH7iheeK9hA95aHqMiz4kph5tJBCPia4/IO/7UQ1aME
Towbx1gt1IgbEgQYqt7hAkSz7jNysY+DX2O+bGwGjMixplSutOZlbKkQMA5wHQb/IW0vHrhjEulb
CoqYMfUT4angJCYC3XCQDLGqqYacvkFUcrvPVzuLHQELsljawcuXRAA4SwAkkcm2UzDdwsUu9KJZ
5a7GrmQUpLAARsEpleUGQg3LppviXxQts6UUfBCJeJPiFZdJig1LF1Lqzlm6V3aWamFBwIw8dtl6
97pUy7lT9TLa8FSggHinXkHiQxx7S92jKtMXfqm2YpALpmmtQP3IxGxlx7O1HFdPKezxk/ZIoquD
zYIiKROnPubyJ34h3ha4SlA4TsTbwoWPybzL+TYVCeQb+E/mI7H/GYtgq9CA0kupltYh0Hn14wNp
QygsBlXv0ej/cVnt8Jr8xikiumHfd4ufREUcNOKC8qIQpIudD7SWSmsF8UwtBxKgOxnLb5SiDzTI
GJaXtOuKAY5Hd/GmvH+MiO9ZaYyKoY/BQ4fKQgOGYsW0meyclJAkv7STOzN9PQJTMeukUaNfROIe
gNpy/30zX/XS6v8Q4O9n2pSNZtcDrBWrQNctIMCOebfvq3S8XKJSe9lN4RxhwamaUW86G49FIM60
eBAH0oTQkZ31O2doN2x9ZrnZ9Fx3TDg8HXJBOcujH6uscT03imdnDiFyQGe/KpotTRml+gKfVb9X
8NJEbqv/Pf+mIcQ7BJ9anLolqF+SAWpxFhLPZ/GVhgY1HYhK/XyT9+qsNBm4l7WvqEWSxpXPZQvn
snKKQYqSJLpdrNKkVO0jACnO9FZtatrDMKjld4TRlT2OKNOT5BjRU6y1v3fWxx1WDrsaRfXL0rOZ
0iuYcJ5daa+x3hBWzXi2hU0b5PIeTg/rIGSaj69/Z5H2Syfwl0ji0fuasJr8cz2n+HLO1h/oUN2C
qsBXaslgCzpSh+qlMYkSa8gXx1oEJ6Ng1L3vHluUUO/82bD26Re/HNntVY13ySo+nj2Mmts5chpN
32nZlBjf4WzmMoE5DJilphjUrathuqgBeW9CU53wrAFxPhiMt8lfZ10WyFMBbNRxyWxJBffakEP4
6W+tQG8uKu5qDKf3LsIPTT++miI5lRSTp9el6OOAc730aZaXtcvB+t+mfJy45gqFttEt67kLW7Zg
/qYuahoSpOuF3Fx3PUyzfWtoa0wUg6aQwk1j7K0E3jppf13bahfItps3A8Q4S/KHPP+f02WZh0QI
gie7CjzwsXOChPpzy1ZxoaXVfLDWcnsDz9PObwtQSMyqrVhR3RTvvrfkjuBBAqedBBAHdPJ5z/cp
mVycAXulc/TPDva9b/3JkfqCM/IfxdvBHLXZ2w0c2R8mB+2Fp/aoCg1oVpxTvZcfnojNJhWntGuP
llz1bI5XmHK5CCGQ9WYaSnMHwhVQt/tLHNVrdr4RGA8DjUNAxZQUv4M5P3PywLH7urUJUAH+1fpy
3nuqLdezknVg2JeXxEVp8H0cvzPzmXqN2MizHhuAF9myOV2heGhTKLm6J5owIZGBb5N2oKrhiY1t
gEv53Px1uXYFUw6gimophnfMT7KTQhmwr+VZD+ltrO2Ojbhbo9DF0jiQv9GzWvhl7+c/NEoCEMr3
CCwd88qIY+lM09llGfG0RLqKgTaq0I1yh7FqJPA0074bjOBkL/2lTAJAVYNp1Sqd9P1k5/kCYy2a
W0Pphi3p2KbOc72q2VsgtFoYr/KZebV0bxHSlEBkam3KaSmDofgnmtOQwy4xfQVAbUXj+NP2yBej
M2JPnshKxLku0dd4XOc6sZLIYUTH1YiL8L1VGqW8Pe5W/jGFwq6zQOnh2PEcQQ1qbCqYKfD4vzol
zCpAR478X3izyfkxNyxQuAkm/6lz31L98LTy3zS4ym/NAFOimDTfgm7FSS/+G6zbAvtAfNzZJOPJ
4rx5mobcLdHBLCegEpE04xhbDBRkcBWpLTgCC/tmktvVX7HiUS3d77kb/ZkIONa9gkV9C8WX1dCY
cz8tBZLusNiuXqaY0pamglS5cietZy5TEzzelJcK7wF6Psin/FMpvE8Yqjl9VgjQ0LE3yX2CStAR
lQ1KRWDAcKJsdC9ZGlPapuyEhJ03jJet6JasXlIYygoa6xuJAy7drBy/9RjGrDszzAr95NJDDePL
WMRC0r1/RqxFagFiIHct9Nixj0sVLBuxBtQx9wz3IvxNjoDhOSeb8fbwSSmslKUcENHo0OAny6KM
NqInzyJhA+qMY/yf3MOz8kDSzSH8EDEgL56vgAADarOQDFX2QAfaqSdaExffeGnTtiWKQRFDqB8y
iLuUiriDH/FnBqpljG12P9ytcJ0+m0eRAV7hJklFAbQI1ohNikkwAJp2ZOiRQ9uBtlqC3xnnAH1n
8gGNPDw2mThT1n4xCM6bbjcnrIUNzcQEPnz/i7AB/cH2Mw91S49oc23No+GGc3rBKRvWShXvKXwe
CXf5JtLthr24cjj8OaUn3x7gMGTohKj5e9wWWcsHSden+z83ckSUVAqlYUcycJH/qLNw0mp64VhK
arF0+oIRzoXjmcb9KTQvLjo6Q43LzcJ4ngGRrOzdePK+Af0BtQYSrRCfIDYJDhmUqOZUSPzmETDY
dXEZPfWgo2Py0QUWN8ZYrvsLalPVy+WR1lr1SUc7FG5xlpY0Ye6aH6ooy8IZMoRUY0LdkFmZjd43
WEZWucCYth/LX7d9YAxtiBthVyIqZUlyRDu02WKdX496mwW7kRfogT6QsoUEILO6bOstfmtIWqOg
H2ldfkrLveVuodDExW63HUrv8/hnb4VSDQOrdINn2s+lmQwFnRD6iMSm7n3DNcmEi1Oj0+AHRh8V
e2t0yuZJkK0pEBfOYRzi4pgC0yuI94OAbVD60u/AaLBk0V/ubk2U1S3dh1NpremRvBjmJxHFKqEO
AAsvT+7WJetUeIlXMDgBmLYNMUNYmnXHCAav+01Ynja9mxRw0WuJVbheC5pI1TjLjv+ROc8NJDSz
tUSGBJPppsWFbjbbHcYcw+fbD2IUqEhMPgL+I1shCVi65RzlvxTArhvdexLQvP2Gh7kvfL9Hofy+
4hwWVNiq0Xaz4YcK8eccEo40evuXiYkiLFKbdtmoSsjn0eG24hQkp6j999RU44CWxZBl+8Yc0XN/
BPBY2mqOWsvxDSISquirGDgo+oi134Gjxw/fml+qu38zKjOYVAA0P3Q3BdP2UODRKNxWntOoSIgD
xM8wlHWTMn/U2hvJhzyVTVL05PAxMzN6OUv4HLoYM3MJnRKjLVS/Tm8Du0Q3UKKyzDDKvz4mGekm
XCru7xgz9d7rQbVyvGZ2WyAfAgc2J20jH5a1x7ybxrFMg5dyOwzWPbBOFukbSz2tr29GxT/giTOA
PeiYTnlFwjuVVZdLG97PsTZS0CmyWbic8SLJE4WvhGSNw6pjtD53ARffawtGCBW/LtE+NdruGjRy
jc8XQdiFCdjEPB0QUppMNg1akGxn5ax77iZD0vLyhTpBGnVhQPZe30RRNHoBbBs16w/GaEnDot+L
CWB84YWxyOUYpvjFcCVAzOSd9p/FgEWCRoaAcJLoxbOgB6ZOQxVhaBKzKr8pWGFlbC5K6DhGgSF+
ssUx7MhQNGB1dg==
`protect end_protected

