

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
U7hExZJod/vUi3z5N4RSr1wa48P7uP/A8O0jgaKOZBD7WNfzo6GmQd7doggkH00XJgs7nLyNvPm0
0zWCfXninQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k253ey4kkVql4FDzRxE0SZp0nnUl5fXV3ls/4mgbh/6ghGRjfZ71MsiTZ71s3tpy77tZHD0rpNoh
xUysBr1hFwWkTjAISVTsWyokKm82DELzMzaI0lqt04f7kevY+q4XugjttAECZCOOrrnUQb5ODPuL
TN/5/7rekkgE3das7WY=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
WoA52aV8kh0bkIXA7aISXPgNn7kpio3O4wNzPv7z4wZK/v9qsQ4Fa+1FXV0tZ0D+Si1URd5Yt8PQ
TB8Mp2LGBm7aAfzTAAqLpPZr3KRYlBsnuQptgQwkquHJi1BcDR3dhZHYw2oUKeYXBoZJ80Dg1iyE
mKNc2EAX8dBe7hH745fnWjhDqr0z4schwVFz8IHUPGI/WDdrXtDdyYzuiWdux2vjC9Gao0MkqalL
zCFAkEPTT0xtWcvaccmMU2ICHf+NVjiwhEmFT/vt1jXBw7quncqpEDMuzTHteQFztMFqsgBfXXAR
/Q4rfhaHiuQ7xUCcTEngpAsL2ypgKweMgL0LDw==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yb4xLqu3x9ghRLjHN7QkYl0tDMsZMeJQgGEQuxDwwPb+acIMCaRAm0LVh6gbF0arOSlfOKBs+X6I
1sCY01AUXvqPtXEUt+RvllN5odbTYkY9f5RujZ5aQ9olezUe3+JLEML7oIeJ23v82E3q5lEn2hpd
Yirga3+XXZGIeEC2Q5F3LdU1PK/hOr/QQAn7r3cfSPSRAYJBv2q0KFRrpHEdaRVBAVRTnMADnWqM
+83djfdVuwjO+GhXELQ+rhNH9dkL0cqvHYfgIcRG0rYfPORpbXH4Uiizi44H6tpqRpTeCgmUfW/1
kW3FxovGX7M2+iedny4BJan5eJXy8iA1/NmnQw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pj6m4D23BtF6RtOvVlnmIzux1ocpf3A3ahzdQxUHuwpW9nlstiQd0oSmGGaiF66UD31sHUT6dfQd
yKhb6vxivgHto8LAAEiyTiUmNTH/c41wB3zGzcZFasAPOJZMvUysBGURofn88ip4eLF52/qIKVON
l8AKPEa6atmUOWXPGRix1yyvpjUnvxZ+wFAbBvP0ZsReS6AW7b6zRE+vUOJaMz0EaWEMMRdw3vLT
W/hp9Ruis3IsgHsdn6M611ZJnxSa2tuwXuWdXURUJzFjnTsi2R7EoD0bDJINDuh7T6iiDjBFdO8L
a4ER9/C3EG6IOxU+oP2sYgSHnI7dLthCIjJ+rw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
B2bb9hbJCVaDRqGS393PhTqcBLIIS3eowUvDjLX1RVvD9vYwfdlG9rjfAUVzitJwz5TOhOabACyb
mMpxy7hxgVO56ex26Ce3uZlntRRrSfXZFQT0ENioLNV+BxEHrr7uipCant7HxRFrLFt9nR5wi4m9
ZZq5zS207DucLy0jTX0=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eqzUQVv3z3gvc1IAF6D1gFpnG3jJXG9SSewyb0B7YFlkq+2WoV55oUnb7Smo54ZcwqBR15BnF2xS
jlkL+wI6xvjzAFZaDFixez8MkTdRnrNZscyGLFWOHz7RNKwEpAxAm7RSsBEcZUaS6x+lEu8Fai/i
gBi8OQLkjYbSnKt8sfNmpRhCWxhkRR0QylraXCBqvJVR8s/2S9YSm3zj5TqvYxlJahDh9O3V0iE2
aVTZ//VjzAQrgKQboTMB5R+3O0GmOfi7O8vgrOvK/PiOq6kVyAYEvce5/1FU9VRi8AQk3Hi7BRZM
1pWTxx+bC6qDX+NQvgu8HPGpHmqeqS/CQlftQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 506800)
`protect data_block
x6n0cBvIUxxuBbFu8KOr0mqMw6LwP5HwgAMTOncVsc2phCaE0eDX4kV9250rpBLyntowL+RuFs1h
ualJLHC+mUjgHzfszmgpMUaoPI/yTMZixan1BpMm+Kg0Tlr6DMKGIkipTjfisdEkM6CPnzrk9UYM
DLGyU5ustnvZ41o4BZ12AkGEA9XbPRbdzh6JGKMfA+aZdCqQYVBg6liUd1lIwREQ0O8uFHQKDqMY
VtHKaAvOwc8bvYBHaZaF18bDCUgTtUUE7qG68jxGGugYZfHtJImdlmY/eSAJdigY1toOi0zeFVRj
XzuxD8OcbNx2XizEA163XRrSGQYJ/0QQvulqZOknFFAFUAovf4ObCIaBKMzrBsI6rIGLcz6Q/G91
nMdULFijOqVgcYDcfi9zzzXSOcGZmcr42jP55ElWzGmwODR739Vduw4BEp+fNtx4fy7Bi902IXOr
GyUIHL1muLfdcPi9sUiNdM5a5ILNzMwHF6/1Ut3hWXiA+MHy7kSVPmqdO4aflC7ujcnJ5mCRJGkZ
EUUZ/yzVZ3S7Zmf/GoZkjl36StD9c/zvDJWW1ihSukYYLY/WlZLSXHYqoz6M/um+2V8oQI5TwnK6
vAC62DRBNZWo1VMMDm1hyl4ARIKW+PDD+JweBCsG9jJUc5NWokaZG5FMBXzrzKxrw+xB1WPjYmjP
fQHR3iV/bJiY2cGAQYPOwRjk0VHFUzEKD0z1ZqhgY/O43LfEe16Ka0njUcE9qwuENiJV492AjPQ9
vHm1yd8FZxusNSzLhZBhyynYapmwB6YRrOpCt923kOo7MKSARl94V2QVnR2HihXcdmgJLPrZp/uA
Xei2bRBD7Z352vs5TspT9xm7K0sqC1xCe9h/SiLNCxeNwtpQOP+NbEnrYL/YOKDMRDS9FODEUi8k
QfU2d/nt/mBr6G6Pl4rYWojXaroL6jNV5y13GOH7bV9NE+lWxOXLf6w3RECcxf05j3uksQ6dtPGK
qzboalq0+y15n7GgcWQry6K/hlGt0x8AvmjnNwGoC4ASqoEV4Kf+xrCZ0LbZdSXISXZJFvDGiHk9
GO7tDPNP5mYmuSmYcrOXbErPDdGh4sQBp3NzXHzHUZJaxF52WMZJSJUyzCaQ+mek4spyx85r/Rwj
Pf/Gu0RzaOdIT13MOp6lOuMhjBb2G5goS4qGt1LJjKV58oHAmK3+ywB1m6Xr16pZ2fVaFoVyPa+v
umNxyyUbWm9c7hpVlZ3IxcWcLEg+mMytBgO/g1ci9sOpAjEGCk+UtM0YChsOzuSchuAUFN2ynfxH
dSZubKdBHUz8kErSpX03BxjmRntY8uRTJhcesd3iw9p9RO66/DQGg4z/h9kndzVdNsDX3PT5eZeM
SS7ZrUDdoKt6D5mgt+Qmi8i/2IP04NaMGW3QXXDtSkwBgu6TTGciFsdRve5KxtS0G3mUbhbE/+2x
pVgGWnyxfZ84tq7fHgDkOz+Fiqe2I5eOhqQ7/ETvPYw7Oi1ujJOpaVhDuaN3Q3uX2Ukv+zHp7lJQ
woJpp8AcX3ToRaofF1+Nm2GLAJ6AM+zb8MSDrAWElnSJopEfEuXVhE85RJ/QGRgnxVKj08Un+SC2
lHSKFB50v5vOKr4QdrQXClQovSqfyVfNpjlh1GrvyEAjPVRPAl7YbKTlkhub7ouLIdBC74VFdj4U
DQq6M8GhSOZxB2qG8zdeyYonPdfaz80c+YybVcaSDEnbVrY6+Ii3boBNRiCIxrY08jzo8AvYKi+Q
EzGo8uV+ak6QYciWOrpnO61BT3OuY6pitYT9SlhLG+dfOtW3d7g0eGGy2P9QkoIt9i8tRRQHiC9/
boL+cJYljixN6TTdVF6AscFpPT/9+cH52t398UWNryRRG949wsuV+ci5EbFzf5vOMjutWG9aIO5R
V7KKGpKgIcXN/XtP+KVdtfWrNPZW1q7/4OUd2juRHJn/tzPyAO75DlKvWF/OIsl+/3UkidOQmVcO
ckhx4V6l00AQlmp1fBKUCwfnJVpG3DkS9TrJ9R9gZRokedTlau/huXUPHOMv6YJOQUIZLEPO84iO
Cu14evNIOTbkTAqO+4zNajxS8cknBlRA3uFTLdMnl8LsddvmyMAV1BquiFGsMxgdouCX8jcOOJhK
LmnPPim14fO1LYwvAtCLiB+AOnJdO8///4lfPZBRCpgCVjhDulOKpR25V42gntyNWhj7x1RXPu2i
NXSmLewmMQBUNZ9OU/SHR3DCG1AloUr9+f401zpU8Ft4ZEzNuYq0Y1mPzkyAQGLfSeSVcY0nOink
KEEnoSCt4v/hXYE1LEpWat3s409iqC3TeFJ83u2Z8uOXy2ufLMnUgQqosDZezaUsYUFJpF8j2Epo
R6r8kb77tUWLHS30HujtcmUU6feSez3KpV/huvRLrmJRZfJf8c4CsQbRE2Opzv+4Krvr1Khf/RUc
7+Ww/TnZCXR8PkhKn//O+6RAwYs7bJzYunrb2MUz82ngr7SPXbIA//1IObCDhNpSYhV2anUHgfnv
8ERj1zUOL1RyxKR0BhAjHl/WlzPb09yQnxGzSylgFdmM/TcrSd1ja//8NqzOLq5LXa16XPPDd1Oe
xjsfWzVwJdtIHWH+DE3L7t39bIfBsD7mwb5mHpEv1Opltv/qOLcmO+3W4xGxuTqLm8O95K+Ooul9
4OG8FfxKkVSefpy+Rx9AiaC7UdBr/3Zq91NqYeLNDYq8gFLS31J6HKU9iQoCJ9jANRWOABg9sFjt
zl1YZVdrSJkfKVkdG6SSszCIhtz02a9Faw+sEFUQqXT8dM7QljFJxCkvBTXeK9OvDd2RUOrTsYmJ
DcIKaXXGJkRxCq1vpldYgnUSTXH28+9uzbw03SBauEHjUB6PV5uUt/T+yauHAStxQ0dOhRXuN3wT
7TaKmOnwTbjIaJTWoN90/RiStcqaxwH0tx/zkH/SbFyucVfuGsv2S1BOzCwurNwEJlSuK7Row7yF
xk3bWwfNYTN0xR3p9LzAJ2KVaSZW/8s8sPz6g3jNwicIB++1DDXgo3lOnbX3moU4pC2msuQzEhaj
BD7pjNd8u/2RH+kdkV8VtUe12Qm9uzT20f6EZa1r0hS8h8Tyiohi5bHZR9rH/UFz7QFjMb6XRhSV
ZH9sKyQhCPy0bc/q/I03SJOPlUGKocIjHXAwY6KUZH0EDEhf+7IfHXPjFKqLALysmE4FJtqn95Gj
V/A3RyF03bRKUJdSF2jxWb05EVO4VQboBe+QIyptOpcGNaPM1YYz1v9lL6XcQEuVye8rJqqx2SWu
ZYXg7TnV7d1vuy4lsdnjqaNIDJlSxIKgHygnnuVJs0bAegZ64nKZd4MgkRqvWxMDEfFckk2szpk3
yuhq1bIZ5uom0eJYna1hF7rkmIB0SjmvJky/bSVhqO6yNNNtqZiMhl5U8d4v8AQRH/1RbO0kM4KP
TihV7+77YEVcSvf7ENtTLSJN6dFLPy3wH2jM7d/LhUWDPacRtppRGbQZX+qqNUqSWorjhUceYmFW
PPUfr84dE6G/wmb2wJgE3p622km+WP5eg3tKJ/iZk/ucboiTOT1x5O+gN0FVII84najRS5ZyjSlZ
PrvMRUtfs804htp0dF2gR9vIrArhuXZfo97V75lrcSCzvfkUyjaR4fcohXG7w9MrGScRG5Xh4bwJ
NP85i0vDXzB/MgD9NejS2tBDErYxwXzycOlK/YxRQsrEF4+VbPF59M6tNO1n+xEnWLxX1Ve/yfty
Hnl8YxdVqd3FgrPr2o0Wh03smQGVPf6csyapV5JcshBcyz2B+0h2rDAhkfgkJw5F4OUITLVkq7ua
YV13m2Fh3geBN4OrgUYRxwU8yc7ABFwDiVE0RRLomsUEI2D6l4E3B/SN8p4DxbZp5Z+AOadY0+PE
S/PnW+k3UBy6lTYajVICnuALV4wPZMpasfVBVTZerBqRyYr2Tb02Y6IeQ5e/6Yo/OwIzOSMF5a++
rJ5t/8NX5OnJZpMmHKu/fHv82ckiNfeJf5lPeL2oyM3t26RxLVgHEuKoIGzBHvoQTUgJBtUp+WgY
tMoxli0b91utGE5AeftVTY1tC7v9ki+3sJN4zy9A/ykQEFLnioKiCFjvneuYLIDcE7pqhmHbEV5b
8ujYUcbUF5x73zm6fHIM6Ybl60eNg/w3VqMgdavJqlwzOsxI2E+KtBxw8oO0U1avzyZ5f13vwIfv
iDP/BbiIGvcFsJoKMbU46NRt8hxtJWBSXR7MxAgKZMx3LrupfYq3pfKzTaoV2/v2aM+rQkum5s0R
ACXO0nIAG/bZbGvYG3krijj+cXvgPS/21+tFK18vtyBM1AQ4OB1kqHTN7PFWfvQQwYMpubyzNjSW
5MLRgMfUEB2P6UzFpSILFDUgyjmGI/vgxm1vtVw7ZTq1DHS/JsEwxZ4bDH8u5MJbzVFZz95l38Tt
5f+W6spntogoLAYJEjPkDx3CxRlPNoebgr4Y4gIkGm8sBt9MLHPj97bVz+tEVsra/Je/qv8c9Gd7
5T87C9ZMLazeX9d+pLFNsSEx1oAalo25+Ry8rblsYg4Uv5sbTL4WPwwOJxA4vWFCLtTRQHSOBLWt
XQr21GNlvWToogW6H2ik4/AruQhSsGtcHVSVmzAgguypU0Wl0z1gVHDiGWoIm3dV6eBr9slxsZW/
/3yI5Vixo57B86eC0bE9LOX6N90nHE+zH9OPAjWf8k22QuGgmpWWGSKcADen2/+LI0e5gbxUae0+
uyQ44/sTq+NlibW5L34Q/uJjV9wx5BRTd0+MO9DaQZ9I2UdCf2UGr+VL4IzqPrwMg0fT8l68Xbjw
kZd324uLpQoZkQcHh01gVhXkYSZa0nDuvoSwiWBsEPamG+yVfzUBhUsruO2x//ywhTXhrn78cG06
L1Jw1j+ASzitqkk5CZILczIS2NN2G3fkqZy+sHety96aOO/UsvErXuuvJ9RcaSOisvGKCRqvy1aD
yUrbNkpMYoS5pm1p/pke7/DOex8w5i4vB8Q4k447HjPO+8AzLzeUYZjFM2Vd8PAo9dnsceJHcY7e
81NR1ei6IYS6J4O4MzbzksEmElyXYQ9D3DbV1fRBrP67+e8OrJMj4oL2ytCKrUbWBrgHnrlHXqgI
NrGg7A+MNnKyiiUdjnTpnekCX4x+0EhxfYuj1IgLOkwHhtLEUVHI0Vz5oZlemPzAoIlN6bVoRGED
f98yxoWMACFIpk0cX518KL/yNkIoBGo0rUCTTKj2bBijHXQvK07jxeqdRF13rAOMBD/+AEB6N75y
YdjuHlHvaovthBEQlyTMasQX3MnNSCc+K4SmRL84g+tVpFMVJF1zMd5rgyZ5x/iveqrjGFIyQOpG
A997vhri+9Y/E5JxX+GpAnBYJYu8OjBUY6RwSABIefpiT0ypJEmbwLYTVkYuNursVJ8qrXyL4ptk
NVPy2aGSds5rRZlS4knHQ+N4pWM5q/LE8PkM38X4Hnk1T7RDxzCYhI3LR60D+GLEQzNZb61ornoF
ANarRErbnXu2mRSHomnvzVB47MdH9NMjU1RNQnn7LeaQW6dsf/Alo7nFIzZIPsmpnZfhBjmyxPb/
0moQhzgq0Fgu3M2t2/9FGd4V/RcOljq2KReYIEig8uYe+tkcIgmJwx5koqKgja+5wk0UJfsbpec6
tvKbH0UTib0KLsUVFG3YQn99rHW9xQpBRMWTv5+Dl1hCgDqKcJbBmCYUUUFeuVloYOV0x8TGdwYQ
qOyUE5OSvxfgmv6s5x40Fn/46GUafGETKDAtmjcZXwL4ZzRWfoSv4q0vdx1Uz0GZUY6jfK3xQQA4
sMgidzIZiC1kD865kbwyCRNWhPo++ErdOIamhAuAjXjKyAHH8Hxbd1wiPe3VnmYV1hq8CIYV7xYU
0zclBznK/HCQTnyJE8EN8MmKzJrTzrTHvt9NXG7Ecs1xFSiRwqeDK7oBF1OmEC3smH1OJZq82RNi
f7n7ye5v7L0PI7MW9KQbgrTU/er9tqAXEJKKgFWRv9hmCv1VKZ5pBCJ4ikdTKrHNYqu7KMf01Vs4
aDpqGckDbT8VX4nxQ5a2XkvQfZRutKvl0aWuFLY7JUlAqsNyUjIRP4OfGLZJM0WSfKyNExkGPyoo
gq14uY47K8OlfVngBuWjM9A0gR4qfFOXVV/JORxLI6PE9jt8ftyxBzc/zS4Z2H67ueDz8iE0ZDO/
k63PiMyu4J3wZCs6aDNIKzhjWjPncqSrFs5lR8PRyNa9S2ZUq2LwYFcx5mvvZ1bw7prpFwBENm9/
T8kG1KxR3ZsePTx33JVmJrggW0Xs6o2XlORAGJAbasXQnkhD/U8xzLZ16NGLip0JOIE1eIscxH3L
f9cUIxW/o0oOBk8TOZ73vnLmLJhN9RO2JRlMzXSO75pWi103WZG7IGcZVZ18LvBTDJY7EM0/GqAg
FcyYCnPOdi/tC0KfBQzm5Gxtpnjpe2nPgE6AsdpCJJODxsbWUr6PdAu5j0HKmMfhOBE/0nb6v0VI
930YQAh9JqG9NfEhMpURI4sZRtolmXchk0k6AuWLX70KgX1CguN7Pkz6uY/neihSf9aSGdDiaMQP
9kA6uQyHwFYPMzVg2ReRxe6RBWgtbXj0Eiz6i2zzQTt96X1PXae+5VzkuRpGB3YyDWapCWDYp4NQ
ZcnIBACIMnMRprDdXaON1DUIdndsHkIhOvks+pm1HV0nhdjx2H+lt5t0wx+nnOQ3wrei5O9pZA24
Ty/IZ3GZou86ETimEbs9Ebk3qju2WrkN5ayWw1noyt4PwH8EC8BbyWXLI4G7WHeAHSBzCvpa1+Nl
pm/L2iQ02A4+mLSyXyLkrQtG2UPgOPvUlkUggvPDYU0nwGQfRu8IIWVnEIIPCzZrSKDhCYDdlzaF
KpgZYxW7t7/0v5MW+THORLCEJ1p7ehdnZl8GsSPuFs3oqKE38olBXPwds0cJdMVVuqT/Pz4w4LN/
+wpzV+FGFfBAUCuoV8kZmb/5PhVOuEqCmIbhoF4Xo36RurF+29k3CBmtida1pdpi4IJnRorulF5F
7fumDMkS+TkVDVtUeo19Kc4ecQ9k2SXTZ2lamUTTHmksoNDZlCVGeWatB6mFta+/HqVuoEQN4gI3
GqHFn/L6+PNBJW7toETro1zWT2PSxdqOIPp1K/+2DSgvCHCQg4RXruAcumY82biog3jLuMoWBS8a
MTsCAKfmsylWaxmEobjaag9hHtdzqhVIzIoPHW3p1+Ow2s1utu14r6+MrAH/cztCTqnGtswa742x
yekU7WK9kGUT9fYAtC1dqm1Yu+3Wr03/P0KDX5esB/3Oj6yyxm83acS0cpD0iBmkufQtw/Cg6P7Y
hknzA61Yp7YuZFyoNKHCJHSy9sKKU0xriKpBhMEtCaXZVzxVNiJhNADI3Xyqwzh+lKBexhdJc7jQ
YJuj1kmfWp7QrZF5Fe81Y1puxzZDhUeRIcH7Qod5Mb30JebBzANgPYN4frFdjffnsRggSqNC27xi
HIrspATRvX+Mj/KhaUO5CdJgeGC/Ec0ECVnnhmm5Yl2c/nQa8IPaJrIEnurJQuBc3GvyVXucIzTL
PV5zHLbcaJCIZ/LrDD48DDWUhTpdmx3t79aNT81hyOdapX1uMcCKvLSnt+VvUc9VeLfanXgZXV/C
WhgA0rYcx45Wi+0EmNxHBAOAh0bxxqJem8BWzFjkP7jBXoUDQQvU7MI8zLXlqL++NwVgMf8KypZ9
A2xOVrV8Wn1532XVq6d72YYS736Jb/5s9vP9Iqdcr+2bUpyWb8y0kFkTfTa4LvoNan6C4yEHcMKJ
oRJe1V48pN2vq5FwyewinvoAYgRf0hnFXF4PWqDEBFtU5+OTlInyGonBlc4NTkUiN5TDjEemxTYl
AIOelRwjl2KgpZndgO1GIFb30Uk2sohVfANb5XESMF2UjgReDk0Az/U8PxuuoKeAsYLb1MCQF0sI
0NT1XUrusoGUIG/03MBnIWnFS/Ro30rauQFwd+YE17B0nW8QyzDkCAG0AaeU2ejDIlOu5DoG4rQM
d9UW5bwFIfCT1D9+vnefjzGLMm+NCDuBIomebUo6OaIxrm355QXKv5avYApXY6jj89pDsZkfHar2
Ej35qJLQj9j5VReZVoyvqYI/WnQUTvemwiiTYdQ5BdQxMjYooqQtkUS98HW6W4lhcBiin9FzKIH6
9N0gEBPMbqbsG/rubi+vUOJx6+QC+QOYzbkmFYK2N+iXeBe7Xk+loA8dO0Y0CatF6go4bXy9PL2t
lhGzjafRXUva1pnlV+eW8BcxeAELeZicb9m3cPTRsy4oxKIGCtJo9ICaR1nASoErzEGZPn6T/Hry
YP5F9BMXshVFgKPK3qmbueJj7N92vRgsvrQQjnKI5aphpkWcUCOCzsnY0YK/IAvWoFMiZyyo+hL4
TnA5eSqBWIJg1uIB9j4KdVMVd5n8FoWU5ZpjweomkUZO+wMPZTIuoFaf7IkJx7Q9RGFRPjBjIl9h
6H/HSVnNBPr/d12C/bxjYlcvgPOnWAI08jvcVAmvvehRjGpobsb0JqU0AaLbmAX2eds+J7vuE5WD
v4ZET+gXTPCOKz8jt6P7ngU3HiazVoqs0UBYHHETWiErRVkHc/YhcXcq3NvQebP87ADXlS2/DkNM
0G6wcY1fynoMvhW9kelCCEpNAbsPqNFnnGeTgJDJkdJfwaELnib3Ji2/JiN9ey7ycpw7A8T7ew1j
iRPTXuJ920CalYwKZKqGaGGPfwfGCwm0AfiEFjT52i+/pbdxFvLtRL0+Vxore6yg1bGpM0MCY6aP
NMmGUop2zuFf5wkJaixdDWz66eQ/xHHZFXZqeMj/t6jLqRM6M69/MNzkItPX3x3pygIGOrp/GvS2
i1EqiuDsC+nT/Zg82NGZWn4aQY3EjagO3mdDx3Y5YWot8Vosf9FI1rwWerq36Vl4E7zU7QVoZWDC
2jXh5PhQEGRsz/8FOYfk09akJzj9aXtE3LCXligaih1cgrqhjs8T1hlR0bLzzoeA1FSBqfV1FbuJ
oOSxic/cuA5LGk6Qcj6uOsLHXUqBx+qeiuPNUI4GYF01cMa8Zp05TTy7NGMRsWdRL2cQZazdMz5r
GaHf9ZRvKduuM1HmhbOojqaXBVcIjZYTfiUXAzhIkaWqFJ7JQzA+qqo3NdEf0rX7sxwteiamp92h
EZy5+oLftkkOaAaLbcjzrNRxsEoTvuV75fgRmR8fFgejHYh6MqOOSx8iOhiPtzXaMhM+4BUmwiIj
hmuQgmThoPEufC5R0cupQlavS4iImlKNn/vzcc9OFBY60/AWmRszPe4BMUCggkVL8aYrdd2ykboz
3EreHn9/OERH++BDdz2M7TIxMgi8b46ycOhEzPqLys8hQggqS0FAeRU+fl1JvzGPzM36i630sCqq
2mfS6zAIZAerXKnLHZX6IyVZA+L/vAJXUfMXiVDDosO4ioR6l+yNrElWBj5YOz3KX8H5/gweTXvg
sN7iFFG+YajzyssphGblApbiyVtbzStrn51OnFqhxPn5+s0YZsh8S0VNo1NGVdn++U6RJ/5LwHvt
8JowwrXQvc0w/ON+6jVnJ+/ii4EejfBZVSn50HPnwZFjOjxSbqZPmvA0/P0jOg9Cv72ja+fCwzdW
9oJZBtE1pojqr1a5K2J1gxzZJjIPOt82q83gNAnntOsB/4D5scOANvT0arvwjSBJacg0s2hsAm9m
jqH/L/WwHFRQm9x4zljADyVbZByOyYo+HbHQe+QenTaAsZi6734M0QYgqzl7ZioZ1cvq5hQ9mehn
oJ2253IumoDnUcZIqKlLGhMxo9XMUcGiCwvrf+fdkkaozIr9ZbktalKmlEMjiw3+wVGOWxM7b9Ir
wtzzqkoklyJqEpo9twhU9msm8ljiQRp6Luw3Ikx8cnKRqDZLXXk3pIJym0euI6qSQ0M1+AH9LuaV
k/x3P0VGbjM32D4EboBW2zWY5c+b1w0HIYt/6D6+DoVsDq+O88yUnEYbRZMJIezYa8whhPTVhCdA
IJx0UeHiPyrKn2qnzo6X3UOLjqv5OOncg3ss/ouQI3rDfdvgwuBf6Obczn8f86kUK+chLmlZ2ioD
vZihr+YuHKwedwtWH46I/VG2IyCC6zqgt94RR1gb4fI8CJswPwuaHtbEFlyVimw2xUFDw68IcufA
5lJ2oncCB1rS6C+jIW2HTb0JSymbY+0bTRJ2nUH4bUZPUWlvg7SLU1dsq/R1hZofMBhmYSMu/6dz
W1HggySYHXTlcKAywTHr0hNVP8pd/jluOQE2h3OEzcvy1rKbYw5STZoMPWaTvcGDR98xgFEllXJW
xQ+GM95bJ7459hKN3jH/8qLnC3RQwv4Zk/5rZF1hgy9fQFxUBvuNg3Y6dBBtXQYteZCIk6mlIWBZ
Bjc6AIMo+9yCXdBak4plGHRiA45c8eIRm7A3s1vIJgTBhM0tDy5r1VZeRI7h4ybOcyfcz4Dy+h+0
AtwTV6fNQCPP85XvfRYlUyDq8u5/LZJqchEV1wfe240gXlommm0fYp0WE0NxD5Leg8/THxE0WYjh
5rYiNIuK2cYfxpc5nfFSulLoNciDX8L2o4yrKTywU2hkGsOJ+PqZ3h9LaxIvGyfQguJskX7KGbxJ
0Ct8UnVmRJ0qD1Y9Kh6NacQIgPowFWgWTwBsg0CJSgr2N1k3JONn8gHStyLePkGZN+7yM1PbMM6v
ywAOAi+Mfexnj6Qd1Y4QscpgcpaRY41S5AxP81BQp0Zyu8tI13tefnOFkaIJyZhhIRSHN+cUXOmv
k4M0/t6WFjoM/+/kQyoAmQbITlWsQONjOWs4HwuEals3VkFLPuuDMu0Zw069bGyM4zTI2lmxT3o4
fbkODiIamC75oSrqz+6TK8Bk1RbGHtNtXUHIsAG/kb0bjxRz9qGKXODrk2NG5/Gh5kXg8f0qRjaj
1Y5UOgX1lI86SU0ssUt1KqqnrB7Wib8t+ceXVkyWNA46Dl8qE3gNofQ3cAm0Vb4BL2XUaiES8tMj
Ah8fEeGiHZkFVos/JrXcFN49GTwW4vU9WKbxUGIEH8a9O4gC5PAnmxv3BIWEMjnzKj7gaoKwW++o
CYGt+BBGFYG6Jl0dwSpZ7gEXDFU/l1tZawmFoO2gB+CYakYxhalgVquOzYGme4FumuDLec4HOSBF
oc5Z8NAI3IM8lKWdnNpnzaDiyvdNj6YiUsHCxuUuzw+QzzrX5tkAA8tyBbTFYhc2vSbf2clVxS77
JksNbFziQmBh1/tMF2X4PzqBNCcJBiFHksgMDVdweDqpgiN8StiNgOB+H55KkNbYlPq3IooLOFKA
h5QQUDDIpz3kGU5TK4l6Co9vZsXy5QU1shRHdL578pQxsUuUoZM24icZDxlg7ELpMrOKd80/GxMw
lKWnDW2VokTa/LEMUmradh6hIypP/yCwtGB4rlXbAmEt52/rXhcTOgWfMT415P9vaXBSl52X2qpf
vGhrVQDbLTb7gymdXAce73uQCs2OmdhYqdQ2x6k+/tIesCl/lW0CmtCkPKtyybVbuUc2Mp6/XVgp
r7zUc1422Wy4lgi+qYMfsDR7G+VjQcek5u043DRWMBbZsCRr42uTrUPbKL1PgBcPGM8nP4sxAYQR
X8vJK6U2WDKPNxTXRbvLFpmNi9jkktmxkchvdDHTVvucEmd58dCA1oHO/mCZ0ECvR7L+aVX3EQkz
KIfO1BngBd5iwKlf/3d8G9ZieEToePvemmXWk5BJztCGubkh2qyHu8g68U8JsX6AQAaMELWinK+e
3hf4zAkeg5UcdGNuxmzpIQ4PlkreEpSIZT0tuSTSCG+Lxe4/UY3vWFYaQSHGlB6BrdcTwitDnozr
Hz4NPox+L/mYn0x/zO9B160XJYlu6u6A7p22+dSk0ldCtynBRGbwtFmiQQzzSZkpjYqkjdMEcmd4
D+NTsg51G6LUGiz8Q7qG3MEA3KFpbCRcntrHTCIblATGufH1QXOVQXUoZLfP5JmCTQIHy9V1gcfX
Ay1Z+SKgud2vp3FPQqGQ/8SL4hbNaHkEW3jLhcxRmLIW61D4zHpIAEckBkv8TyZ7FJNmYMuXCNdz
XFRLDrsVAv6v16N7u+42Lbx0QflnfV8ia07cI+Coh9/8tZBu7xfq2ySXauRwLtoPw5kq0pRS+czh
w1C2Wov7F08uvin/OW3DujvXa2+6wJt7fW/W3DH3udSi4JevF1225ilf2mzVShlkad/uKQIjie3r
eQFVL2joU490wp5XNtJa0uD8dQGlKW5dRfIIQ9Y200IsXpJGrLSOKLg0C4ZH7AIChJca/cLYc76S
5TQd7yIIUCP69k3xiVGS6KAvQeyGGFLXU8nQ/rVMTVVKXVFqTTdMn2x3gnpRPNuSBwDnLef02cnt
piSCQ5+yqm3xfWVheXHMbFf/tHbs5arB0mZOmUhTRhQpbwpnDNrwxv/E4f8ZWgtvNbLS/yk4UUe5
f4bfSM9inpaXLmiT/ukUNGOKGs3jUaYQBwivDg6WwL8/aHhyg3fjODQoqGlkWEwRsNtF62jRBwg+
zsYp/foP4TbpGhqEyTnHwvV1oEJo4MVRqeudC0i9wz1zHP2ABUCmZ/Tdi0gdoyEqFROcVmAYkSjm
7c8KR5H+HKMmKGERLHRzPIwLidMOXqjCCGFeQLB8Uyg2jgnoaiUSVJRotbohQ6Apr/KeFwfLkPO1
S3XLn4KVU2QMBjBmYv8KFWzerK2bPYiMXwt+TjgFgVJEG1RjQtVpkND0836PkFnTjOWRoERSEdDN
yd+vlyivZu3DE01wEvWWBSdHtAsUpBSpfpWh84nC4JkjLvhkwXmbuwpvLFpbjStg87Qr/Gd/D7Ff
BYmU9Kns+1ptezq9UlW/nQp03ZrOzUxUSEwMzjayazbcMH5kHFVEY2Dx08/4Xy9WO1e2BRrU+46P
O2gfUZoqZ14NjBpEXQqMbHUl6sKVzGUCmFpJROnr5zDZoO2kpx+ZYZ7ovofUcT+ZbKG/LMV0AmO1
WKQEH/Ji8wfRiHT0ONI7/XzkYrk3cXmhPo0Fvj3diByQVZNR9d7fSu/a6jn8xMfEqdzS8aHFLBtY
S93EgIEF3qqvPnLq0o9JVlb3aIZr2rq1Mbypytj/K/Oj1j6pUtbYDygQ3P/5jBVTaSUUBMGk2Wkj
sEDIpNsuDuKoLdLTfdqdSm+qiVWOfvLe134kUlfwc3vicXhZVvSbwC5Wt6JB6XlcF1cuxLWN9X/P
OHCcCbOtxb1+DKq0k00BJgh/6NQQdSO/gLsMfDmyFVwlnEGwcSooe17emZfpzLdniuPpahFd/2EM
JiDNiUJ1HNt2AEajwdil1SiCwRshpn9d4MVv79cjN0sPWZP0iXNohSDz3c+O8eDVxHBLdLmuFCO0
CvBbLrtO7boM8DLP57RC1s5o2DXMsvxcbtpbBimNdNITObNkcU+hXVI2ZYTeabRtxi/1qkKvktMp
XxBuloE1S1fzVE5VyR/spKn9bh3UdH2ZxDFGgFrWFZiCTY+zkRxXs7aWbw+2V6TyoR2Cg2QC+UB+
lZDyifk8YumHvyldmcn3xjyYVncPr9lVPWSMCf8Iq+nDQelozzVWM82IFfF0P2Gkmm+8TSSqewbb
EDjfV8YVnR8BwZY24kZwOxIhYxjZGejz+olfid1wQgI/jA54xWQR9m2WWjHfo3b5RiLfBszU7T8C
S7eBbE0k7vJQv0Z8kF3hzcp9LRaNNXbE2bAw5uhfnDT5oMir8kOCtyTecn2mjw8CzkXofJ7egVH4
aX9s4foqbwRgvGBa5BkzRAZOZqto4EOyf0eMaHghi0My4+GvPXE4CgDnmDRSMvKyTv44bDay8gzL
IlU1Zz0r7GORuMuO2qmU572d0Pt42M6xKrUTKV/Ktxt5prVpOux3yLkW3UFDxdMXOSEVlAkfrRhz
xEKvn+FAXMS1amzCymV5HnVvq+QoTtewUmn+8TkquFojaZpNwTeyHygcJg7a33d4sAnQKQf3nb7b
0lYk8+JgnP3uKI/e7x7N2rkFSXgSz0yB1QpeV30a1Z5tlBfXMVC7YdwrkZRRRcCJiwEzgWWIBysN
BBw90DwkQNt4sgtHjE8ggN8TY/sK/E9fwngjjh74uRwLk9HLHqLwsFUAui1pUvOBx3lgZibu3QzM
0EW56S9kbaXKe6m0KPhzMGMtJs9dojzBh6e2VYS48taqfIkAuYdLOx1g/znVd9yiNEPT2OLTMNL/
GPi+JJ/WlNltB9iUjVyMToivXOU27MaYA7TB92fWBaZ5Qm/pQVm51qG6lKgfa/pdeoByfL4LfU0h
9T7wehke3yjgqbSCgJwWRN/OvKgQmDvzYwBXhSEx/htZrGM1slrdS4Q/5+UWj9eCa1wSvSC6+9aa
UmBjb//b4ZfWu3RVu8QQ/JkoTBoncQQKkGgTy5AbKfyCtmEkIP8q1+AoL2wzTgeHRDl0mu0wohRq
EOkuTXPQarNBwtp9cTwZYK6eUT+P9dOqYmEx1F6z9CZWW44XIsPT45qmhmJNgTeeeazzgOOykmzq
Kyc/yptW2QWGbq5omNsgsoTUeBjkED+z7knEaRDbSushlLklJbQGjXunNelywituVGOJzKpc5zrk
C4HHlttSIHVrtXUr026JaIszgaoy8Fmi2GFSFjIDCu2QtZ73lhQNPoZESWzk6LY+GxQDKy8BbRKl
Z9RQFxMUDdtcNWxh101SKy0RNJOa5/coLjADwUA7ulIkTnQK0XcKPc2u0RCNpTzC6+fmE3EMgil9
QX8sv8dxhDRUzWtbroaOZGZDKO+rs1JqH5b4QSSnCSUcwUzS+moif3Cgf+JHTvG1u7QxBY1+kAA4
2wk+ws0V9IwNxLbsQJdGyYRarAVs25/VdOKj3bYFaaSJw3n2YI9YHHBF+TinEuWqxn7Hbg7nyJrR
VoPkROK+MvKfhSXQhnszraK2go8s6ypyCIcmR19HnVCTwJF+6YeXSYXS3DbFQu09gw/ATD0q5vBW
qeuX61cGGu22M1+aRdko6shn2Y+52Q5hFiKhEomJjs/7JHCNaN5jFuQBM5A8ANyAVPr8uy7/YtwM
Scxrmp0mJHODTwzmtJ57PxgdXdM6hBQuouQ6jZ0JdBh+XXmynH+1FFve8NRjp2Ow/HCRxLES5G4f
O1v0os+PI+BcakFKj1c+W0YsVaKSRvX/YUl1RnlGitT2GZEm9xbGfLU+7m8FW9jY5IXc4UdyLOB9
CKDm+qw1jPVjtwLkxlKTOFmol5jBnQFG0LrKWwwhRQZuBjbxrL/5pIBp2zviv025m45gPsDnxOhf
BY5Z6sTtbk+fAEVIhn+XRmBc/I0gUM5pp5hqdCtHbuwLdvH86zu7zriBjekUQqlohiJMyj74l6kC
2a7Cc4HJVzt0xQscLd9/xCK/tRFjntO0u4LUrsoiWlAGAuwFrRXVPGlUy26p0oBfFOoaRs8crude
aAZ9EvbU6C7wlhHVNeKtUj8D/WxQ5kynZSw7weC+Pxv+udxDqSEmoZ9RH97B4koLQ+Q92FEqDaVs
lKiWEOh5tsUdbsZukEhnvw8dWocmPBBke0u8XSaiNuLKdGjQ8F4r0iG2/vQZ0oWQm0iYK2t/a5gU
YNT3QEis6nUfVK/6NUUAQJU180bMLhCprGyphH+JbN2LnvNqKHucR5vsASzYVTgQ5v3P/uUKzPqx
F++V2J0rpyUIcRKThiyy04SE94q7H0RVUWMwcHRZXdUJGeYTncu2S7ALlbwqm9P0RB66EFTsYXp5
gUd9ot0n4OAm8HDx7iXRNA+51OBZ49LX3cGvF9A33HTydDeDpcvW23q4lfFDm0+W6asdlJ6sOoi1
qUiTzMpvsKPlGmoRFHfciVZAJZffjiSqnl5OhwxdBputmoCOolCI05E9ExEShDsZdvK0ikc1lphw
dvvHkqWJ4ltuHjYtxMwyZkwSSxoKzoAbgClhrjsIeiWxkGje+B0xtdt9AFf7ss+ipNGzD1ON6psB
+WkBN1A5wSDB4OavjZF6GabYB88yt1bSHL5F7/IGx+N03g+sRmJGbk+e2g1H/+XT7aKCkNtH9Oik
LwsV2RSxcDPqYHrXwC1QvwV5MbxQZQ83juqX1KtQVouv06pqhv2PVn4xaEBHyDT3pnec8pd3EfQk
k0PG317GU3llQ0J/YxW5gaAFSgVda45ebrE4W8EGooJbp8nq9O2m1JGw5asaNUSv0qhZx07B97tC
+3yjqD+eZ1INX30rPY4crHVmDmeK5lbAzRhQOEdKMVA6UrIiOI+ATwmt59PMfgS5ovOMRqifpg9Z
ffFrUfnQEBpV3wrbMgkWEnbUZssz6E3iS/sQGNBNyOrr1RnhJA8JODf98inoXVWHlpKBE1sj0Cav
Fha8p/BkX49nrOpgtHrJ4TqNf7y241l2Wc3nnI4qoux3FbN+seK3lnvW48r93GR46MiNrS3XbEOl
uBTlrdEtk/kW5y77x2DZ6W208KWcLtIltifABIAo4SVVe50RyN5z23NcVYkRAi/BdCu08OfuP/VC
ITT7gKykh1TBUXLdIq24Ee8QnhcaOVmKb0Yig/uK4fmY5d7CirP/43BWOXJ6jOxnX3D0lBVklrBT
Pu2E/8I8NLZfKWmJDANFI9AecJacwpbgrFdAaS43hGSXYuhosJ/2aNmSWS60ugEls9FuJwDVPbN6
a+lk+FWeB2pE+pMwg2drNmbLSoV3k4z+pDINS1wX6kb7LoYsKbf6My8Tm24datIn1t8IBRFs660E
ZfjDsmsSEr5qkeGQdHhNmhoK6nZ2iPhN890XqqGewmAoIa6XmmKg9/zmY8BVmoRB6bZjoa80Au/U
vD4N8kajebJAROV8TpE8itXyx2R69rRC0GInj88qyztgA1tBUpOkaq/flAJMRKMohzb2uTWA+P8e
K9Dr89nQo3BMLvw3oaNcUVgJCPU4XyEfaJtXSu0/h4+PqkgSSsw0XRIWqBPBGwjOBibLDhjgfT5V
AsHjS1/5iegNMzunVr06HTGACISCrRXv+3xsX/NrEEcQMFP1WghkgJR1TZmeh4oUDSc821LOM/xz
nDUtkz5nRTI/bW8fpdcDfMGX4IDx94roFk8Nq86L4rfjiM3zPuArb+wbflAU4iIbQpkFl5Ku/IcK
BMddEeAsHEttU/qnPwF6vxTH2J0KfCOOFRYOyCevfdiopU9d1EOddXPvbSf9nIaGV7ZCEb+5JCwk
JGXCAUujIEqmD4ubKYv29dcax+CBEGYtREtYx4sHl9UOEr9ex3aO9nsf6yJXEu1AlVjoEAFFoMkr
ME/F5lTHbPpPgKo/EHfikIzFZ5hgrYVdbpUNUl55mWph42KCJ65R8Tp2CCdm4lmASTrhgQUWrXHj
LgKmQexQlL5uyysvNfOIJAmoGPLItyQXDauKBVRCCD73Fp7CgZzhoFs++bihGGff092zzxIgRAa7
0Zg86NsWiN4ovQpwTuChMT+Z/eeOoYj3axRVj3dWzlL65VCMlrNddJV6Xq/Dov3ICTOY26eMmV14
PDAJcHxwbx1oS56Lp+9AJ0ZBsCHTu7JmfqBK0RRi+sply5ODdSPz7v2RdetaJoJOVjNs0eOXAU/E
cAEOHWMrrmDv6PWs2sRmT2d/mqNUTEchwB9Q/TySa+I2UYS5NAa0f8k96BqXwOwXApnkvUpVrgcE
ZG7OJWDjHAN9irEjDJcnqOArwrKxpiD+33hMJ3i6mbz1u1HUNL2jzKqQKPmI6TxPDDBmz+3JQxUb
+VJ6+jsSFXRQL3Ek95EOyJapAMnQDMffJiWWnIw4B2qWDaQEbgLqPHaHrZmpMxewz1o6+WVZJb6X
gKGH99cljSvYVrM2FHOEvW36Puluq7SSBSuXnldzULdNzsZJBKjPFZ7IK7nf4XXiBHynWFgFLMAl
rwxgbMj2rOF9tQgpvBQOvnsMJg6f7kIbKSjyVgg4aTFIeIcU3mTVD3vLWyPiFEDyyuwwenm6d5WV
xv6HB/woxXGx+ZIuJ/D0EI3rt2Wb6jg9RGYj4oYe03RnaGN1Zg1nBzjlisNQSBG3bSNFqcBw1+2i
AVPh5yj2d/C1uSWK0YJNst0b2H/y2l1BgNSme0i8qEKga5pnkhsQEbQmDA6ocPj9WI1wNhup+Li4
ja8Az80oDBFAMxdXV98fSti6JnEPr0R4R5e+M2vnuIDUt8tTkfjOHXJBf77c/pevWj3g2RWUZQbn
xxUdDYIEIiE1WRmXBY+vp51c5P6RCfCt7tA4XomHG/XNBw7FXm5mppXW97c8yLxCxdETx4SyN0BO
jRpjczkiNIf5jpkB0SH9Em53eFiLIi/VZ6JDgdC5EU+Oe3ehwxPmSk299NRErUIpAlIaXkYiyZbz
2MKQK/WaA3sTwISEhhLTmsyqW+ZaisqQ5DwuWcmknr2HyAv9UtdDFWssuk41XKL3mqAE3CIoh5G9
BeNHcwY5ocr4ZfKjpzORQR1Axo501jncS8FBfxzCw4udyIX7Idy40/v/bhlyeSbOXIsxxL9BaYLB
jOEducUml6Z05OBy60FiZheri4v6NrCJiUfk65UO9FPFE8LrnhaCHoBDezvnsRruGaQql/tSmzzt
1ASP0VjEnivzE4CY5u3BJ1ToOKLlq4+tQgFPIsDidO1iX+EBACa3ifoU6LXP3qLZote7JTYxT4GQ
k2QshYIWS06rz2PwEydqFNCS8OGzkFL73KHjJoaAaWv+0sSzkUEN/ZmbMgVNIhGjuH9gctJYFweg
yjDnDRfPSVC8B2NNEwCJeNMFkwFRq3PBKXNAWJXCLCZiK5BWRQCUAK0lrfPanfw0oTtvov6AjBaR
/B5ivngTBsNw5+hq8zHWF4NgyUSiopy22ee/VXXWlv6gBgJbHzLtM/qPJrnzEe+13jd+wwpP3mjG
I8yZMMutLtBIRpVcIFQewSEJv7iCUDjjEelY4pAOY/Cu8yGi/jCqjZx4vhydOL7OiT9c5Czsqch4
s6eIZdIiR6NNg9DvK1cYB8syObYVzJPf4KEwmbseSHEpzZpbvOIiYSgJa4cHbKc/qAUz7h3Rl9J4
g23UPvC/CbC6Uge66J24dgsDygfhrzs2tBdXBfjF8cVdtzGdczD9tLCaxbqK3T+UpOv2Xnjm1p2r
vMCs8ItM5rD1XFGn7KX6aXaDtZ7Qtgj+FnbKdpxvR/ld/1s7UUyOOhhgX/BC1iTJJWoctIE31/Zj
ZMRGvIX+OkebgTqeXj3noz9zl783edLa5kCZWSZ5Nbe/TKDucyMnp09mStQARlIv/uKgveogfNKp
Y0rGnBcrfuOB5DWiVgkDmvPmdQtr9NdC2PznSyRKn5EhQ/xlb1eUKsadElyWrix6cI4i5tzRwd6F
MZZbSkizSJM8pbXxiSzmznRhB0a9lrw7qClu9gFqZ0K5sCe3m7jgtdFfPzUyubFWqsr6X5QebrJI
pSo72DPBaWUIocUlKbe90O9YJxtClgvxvwXFMxvLcf3SlkDFYbM3ao/4pAAQACNOysTndki8wnAk
+rnUIz2LkrU+R7M0i7DhIdJbsPEOfNIDhNxS1U14UkXrahEfgzCDqnKnVWw6afJehhM5afTXIzW/
8uoKKPhrERfhxe2YzdgflH7qA/fFHC7OR98AT91WTEB/ZHnQ4RIAQloJWsgZQppz/aWYaaM4CVck
wGC/GtmU8z1P1PCkjgTjXCZskiYti3LBGj54DRBuMa01XrIG0KHsWp9P099LkghN/HXx4x2qhLHI
Xv42CKXQLYZsDEXm0xS+j/AyNxrBbvp15aC/PL//HIlLL6eVz79eHItmhgmox/bTH8A4ElycoRbB
aiF3vdCAh95gmtU+X4QvMJMdSeKb/cml7loO7iuMpS2vxdr9AEeZ+GD9nH4dw1EdK5sOMXK1xjtX
g1o+X6yPKSh4YuVc7LZlFvU7s8OkBovrRewLvNdWkX+UUuGUaKPSt3oTTEzlaDvQc5B4jtHN7XkK
lhsPOci3+GxTefH4MFYNzDjmIfSYOwJYCAFZcvBkah/of88JHbGoiSuQlJ3x5um4ytNZ1+pFU4Q/
H8c7kHb7GaR9+8gr7+Fef01JFcL0Bmf4NMcJ5rojRZeDl2Hliwd1QVxZHLpchZoikdIVB2XX9PJ/
xoEAoix0DvITGoZknSBT2OW43z9r4iLn4ojv2Oo5JVK/LOU/KibpXSbA+j+EPGiAbStDyx0ZPQ3c
OzvSt/Ho7aOQIE59QV7l3gZH5YE5BOHi4yje4OCUw8tF1VZYL7P9ZnFlWDcP0O7ijQPGrX2nwazP
N0sPUDTK6IcVSQQMOwnV/fn97+jNsSF/zyxPQdg5zEH0h4R4GFtRuj2cUpvMG0dgYW9VHom2BQ1X
6rUECFKtpdXX/HEEAAgQlfqrIL0E2ni56LR2S+KXEGFtfb3rcfH4daY9D8Bc/6c7calIhP9cBA6J
C+nJKlStNy9XY92SZBLbknDI9AJLQMa01DfzD4JnpBSiG1rWEChJqDyfg3oNcmtSZlInD4UfrctO
g09WM78nRG7Dzd+ULm1Kh26BwQjJM3eCFOLksvqReK506i6VAJTVC5lObngDyVlHQtYt3wrLmg1W
uQkpo7lhxeXol63vsuAnVWhSmpHTgyhiB4qf5XHH7Hbp6n/4JtHbptS/PqyY1jC9y8S3VsS9y0WD
8G8MRHw2497BlpuefgN2d+LbK2xDVWYe+yZycGKfYe66rIFjBjOAo5s9YjcbIoq30WYg51Ua1Rnj
w3WX6xI1bahErhidtaq2Et8y3WYDzeAObEVqh2XjSx4uDQLTImayqi2VSZCPhHLlQDEdWF7pdMwu
/faA1wJD9CjHl0DDiSwKo+vnBzdQk2whsd1yRr+jQbCxTiY58+3oSUh7h/naeRGoK6mr4WtUhcel
iVr6LMuED6dgPWChqTsuhHj7GhEt35KogRwrDU7pXfSy9cKlnsLKoxWCuYWShRLDhSKZzS/c6uEO
m1iLrcEG+IDIxYwvXZfELzap9zz2O+0fwoOWg7xBgCg/Wixe4zQjNVk6xs/IG/dG68WmzHAMrIQv
PyX5xDNzkuza4M9ZV4UNRHNDu3KWfs4ValTXfTM95HrNFw4RcLvkM0obcH9if3qy1cvQtzRZhKqm
qYqrvUZHb5meButi1xKgryK8cLzuD8Pcr0/OcirXsVMiJW5yOmk8RVZFy+6u32MBNgAhaphwQfgJ
mLQzG8tuY0OwGwPRJSS6WL4KgkConhjA/NKowhJDumwm6ILSkuHX5rAl9OiuAz9MQg3JOpdGL/+0
9t17KfN6ItXDm+O1X9lwbjpF5MVNx0n+QlHgHyGBv0qm7nRp4o13QHXmChx0N6bxOa9wYTJLAQ+g
9evPwbQclzWAz8XYNYYQE1RXVpgXRm9naNcdY5HA2CtYUREtEAwASmXNTwemeJPDD2SXS3vriSdF
55L+jqctz588HFwNjcqzy/Ilg6qHfWIW3Hkb3gjRpJPC9MOfttcNl3QHdYpgNcOHg+3nVmPOCpTH
uDj4o3JJW4JuwnirlRKtD++lIdWDogwwVuwyqH0KQYdTEgnpVjfQN0S3XbMmZ1EOlMbhNvflM/UG
WkwNQ7WotgcjQpOisGo5tsCWEP4B4tP0KxC0CSZRfhkWzjsnb1YLyfZnBokEd4r7Zn4EboD9U4pm
foSxM8Ecr0yuhHnGO1DzfXbZBHw6HBjfZjLae2TYTWafPBOkCEG5/aeujHwJrShLtiDQ4//Henf3
VavJAoYPsshZDa+8k9jUMGw1vugt9oy7ftZ2Xrq+dYtrVniFfVd58im0iAf7hmkj4oeW+O/sreAL
YUJw3wwMr6PfN6VtQx7jHU11gQd31dpWgi7ZvfghRZdcU6f22LvqA/IvvK5jIZ7WfNA0CLQ5wLAJ
4ue7XrzBJOdALeFHs+IXJYOsNHdDQbpJKg84RAAsJWwvudFM8IxtakrcbSdkeEm8kML7ZxObfNJ9
/ESimgX8o4aCbAmXtO800Jk4n2lW58zfOW/S9CVi6TF6MACl5aaniLg6KSrYYNLtQoyS1M4u7/J8
hAbtv67IqujkahCv8DKRJWjDsp21zWiR+4OygFNT5DLeWdqouR5LS61zJ3iGiSpMOuO6OdSTnLOr
z/DsIQG5DSsqrxHX5/9E9M0BFzM3my0JSAPm0+E2+rUbRpq0QjI6kAiskiXrNC1Y3W00RV0y/smB
IYX9oBKopZ2eCkvc90NNV7THUs7HaKCowD55WxdOFhEjfYQwBgDEuS1tHSe36F2weDd+zZD8bFGo
a/AHYLNUP5zovcgtccO8GR8m1+kjsctiAdqskqRC3GLHPlA4rdK4Xu48uF2P0g1XxVrcCrVZr5J2
bIJOyrhzFIV00h8S4BZzFI6ZTmcFgR4MR3h2gQVGAc38gPg0o/e5tn6EDOu3ActNDRm72KDJiAWh
f3i/UfVv0mvvHJWTGrdvTlUccQY10sVrZfBaktHGEk5AUzFdTmqpqF1iN9D2pO+4BgTF1nZgbGH9
mARtTZFqVlBLgy6wQUL6Zhg/EkLMGh+PMc1qzlTwVnPT7x3NAkAShDtcG3hnQ1OwWmQc30cwZKXh
DaHh/G6hxqKqkZiZ9YDW7TmpvHIHeSBpg84ioj6TS3LRBAPO0drgHkdb9paHLFtXH/1WowF+GS5N
QKPLTDL0+SArTypvH2G8uQ38Z3oA4kBif8xh2BtG0zyirKZXD4rcQh27l7iaU/wONYde8YI3LHta
LWBMtEfFsg0bRHoWZjsWZAbpkic5XwVaPcl+DaawppcX8dEatVXfTl63uUzM3Q59w+FQv2hf70UB
tDQFi/bG/bnMhk5K8WvZ1tH2RuYm8KUJud8Bel+/Y8uUhzDS+vN4TQolpAi82rWS1R2CV3tLTj2N
PhosMvd/pJA7/JCZWG3F93VT/MASgu8kalFWaGSnvB0lU4NS7/qFFfkie5VIrqzNkvKmqyXSY0IM
UDhwjEv0ocOohz5NgF3fI0r3lpxhye/G6L5ke4W3ZeCsybWwEzgFB3BZqrrVupPrdThXtAOtEKK4
wyiIbdmgrptxNxzD9URtFQ0m73DCIAnZ2R9B/Y9KJzhhbyipIb9xB3cCl1eMAiNsNNBQ3Jz4jR9I
WlGbqihA1KvhqqXMMei8tB4GP8jm2zotj6VgVaFo7dbKJ4Qik9eWLQUf8TvUvbCLI7+7IgamBeaz
3BCW7G9fl83XCfvElWWmiyKdPq/0ZTgphI/DBjKIe3AoeRjmmEvPWIbwm+odZlJmahc5C7STvRHy
9JpSWadIutku1oup5brGvJvS81Aha6RwxPpbbMxPX1IBvQ+EIrNZvMWgKHqlUyBRdf4jqgQhafGK
Jyjzx9y+59A4DzxW9k5hr87ZjUUBM26MoeX6VkywAU56IlXKD6zhsJujYDpWZQhWvRFJl8kRPmBo
f6DUrPrhTY5KTkUtT5aG73QHeUk9+7eijmaKL8x2TBy7WSUoIetSrTOC4ceTGqvE1XCrtLFErEhN
IpEyQ5qnY4OdQPOCYGJEocfyTvj2I5LWTJ06wYYfmEwOmx5tPdYyN7jFRwa7MQ1Ca8fXCKccRcze
HKIe76J+0ah7YITMyXNMby1DppgoPxFL65L/3C0av0N4EghicZwsnHQNRn6AmelPtQ9hbQXQmO8C
T713kSVUw2E2t43XoM/vS+YLR7JAq20Ak05BVCSebFaVOah+1XcRRYznStk5nQ2UTXzIUwOACadK
owNzMKO1NoIkHY8FAOZ3nNQ4hsfN4iSnRjMN9hfQKX2tVMaKVcn3/WdsYNRHhWj0mskhaapWK8NU
7fs8xUEzSPHIjJ6cJhRbnpa8wm/K/sHg5DUsel1pm+MSIAWc/LGiXKuhNTmVhcUcBpwkIrVkUkQw
S+cHfAwKN2xWq5F+0gde19tuhLLP56B1MOD3JABK1WfM/HtVAcozVpMto7mgywdXNsWCdn+/OPFX
TXTTRWzcQ9qYz5S1nc1F4wuPEYSGeMObiK9V4IpiOdYpSqYIXL5mU5i8cb9T4j8I8odA3jTpSq4f
s4AsUx/yTijZYHHKUZJAmOnseHC+DrxTWrZep/NYbdzLCX8oqJ3DsNWwU1sLUFBzM8Z8kdaFxr2O
2RBJ+bL3DZQbF25k6btRIeZ/9h+R/hAQJm6KGH9yFnWqlBJo1rCSkG2ScRbq8yNjtqYS565Box6X
oW5l77KFqUi5zmeQ7Gd4CmTSB6m38oMExJ1C3y/4yPxK4VuV/s3oaU3lKl46wj8f3oTB5ttJplnA
u/Hea8E7FdczmjIA5ZHZigaMTVR+bzCCUooy7l+DXeetmRIGkAnaD4ngOcbkdKZKcywYoLWJTSDg
0Shn+1oqzqAZACaYyWlFjGqQOBhS8dFswgNS1tborwhfOfHpX2o0K2XtGFvvWa62nmJYet7m4ItF
iYq/JwZOT811jee3eBSG2xH8TTL4YyqywALudHL8Ltkre0UDBmwElqgoS3w5lduqB196AKZWUBMr
+cZyxuFU+5hX4qv3AAi19hKkUAVr7B3C6jDiao9g3vh/hh8gIGTlsKueuMyw1T0FjUGnJMHsoCZR
/BCZsTlRpaS13IGsqIzBJwb1tDuC8aPKW1psuxJeXsYMGGvyR+AuG7BIMnu85OmytWp/JlL2ivSk
kGo7eNMOrAruKibCRQMvmG/jlQxWRfVJbowh/LCMq0vpHvJWyqn5CpcLHqi3gvBdN0y42PB35Wh2
q3VmxHORJrFHa3AaH+85RhAx4h4gwyS3M2I7rFKhWXrSkvVEFYAIq6AQ5XOITlzBUBpfMmBCDr7c
gpjKu8xVnO+PpsZgoYYS0DOG1ZxeBvmtGHP0BV0dknEVlcgoPEz4PGZX+reepSSTHAjJxHHR7MPI
x89VELxaYCP/HTjcpKEZM2zuzqQf6zO33j0Cq6DqlwtXcZuEg6en1uFB3kOVRDVsofcQ87H7sbWn
bnf8N+0VLWGn/q1w/Tud+PZ3THTLWOVr7c4i48/gVvHrXLQudC0/WMXIDKPXUQByvQGLk4FsPNbi
YUBXXiRH3nPbxpnwkXcI436LGk6iH5Q5Wp857qb4x6mjC6Ao/yFqKEEzl/xJsJDsFpIBk2WqB+Cq
19hT6RP195iveDn72GVG5fmxat/4nkfkwy+TW99tqZ9eodzwYHtMKe+mPgnlPb3fLTAg/nih1xlV
hXStfH4PdQgvxpwAyMTaGa1OPeaqmVALcs0y4/11X3BoEF/6ZTD06KV55czeJGf/lXvqZl3eAuGd
jdso6C4jxHONQ1h1DsfkfZ2iD82jmuAPzxaofQux7A5HELJlGCLuUVGPbW3/Os5FkxNPigS37Jf9
U+BVqD4PV3friCTHoojzDMiw8dC1HWgx9OBP77y4zQ4BPhliVLe3aXUZqduQb9AK3SwGL2HYubtL
yUH3EEsqaWRpS6xcC2wSOMCI3AgtT5Wmcb1l0HNRkV9r6ewfutW5+6SM9lsu4czzDAoXhfEekymK
07e/JdCRih5BaMzKAgu2BJmg8lUYyMJfjwfsJqtOQ/ynYXhsUR5T0zQ9oy/geKEE7Qw3waNlqIN+
9x7qEXcEohH7JsER9s8z2dbvQZ84dqx60OSlp5C3UrDn/s/r747GGFfKjeBqpgm5Q8iPOeRPIIUC
0DeqrCtPXDj3lcZlEabR2x39mnPMDg1Ti52iwfXo2QKwS2LUaqYRdONqpbrLhXkO1GXg5cucszgG
2mkPv4DUl6ypQIx1MgYcjTZIvbqSBKgUHGOx7kp/XaRnWcX56bpCCB0EaMa0KIP5XDvwJYGZNrIj
CGKvdakSzJxByCijDcUZWowcjQz/xTtXGsMcMtFy0qthaovvFaHEJdoucrDKwev21R/6YJx7TepO
mP2plICJMMqxwG8dH0l1LEWGNqHs8Xr+/vc1CD5Ju8iyAym04Aq0/ERA7qULWJuJz70Tt8SHCRR7
RUvjVy1r9/6PSv2Yyu+4msYUtsSQynGYrEYcLEjrXuEPgUTePzOWaGRGp33uo3o3FlXaQZRm9X2p
2Nvjo1ODAS34Z4zk4mqseDjrQzuAxBFUhJBGLryVtbnUfxbuF2ak2stkJ1iVgIiFnb43NgK6TNaE
cgh9GvUB6zoprmp+StutsjMCSLSWNRvcfa9yfi2CKP+2Yn5tZAMUnMGTNlE9Y+HJmbV5jigi1oT5
jPda3v4e3PxOhpS9hLakFT4i0Ml3aNkXzKT19s4HrB9bw7m8wB7tRagt7XS0VEk8XQy7uGB6Oy1k
nCimeATaMOFa9sw3hIw+MzVLqbpdbGNINLF6i/guQtvZrnqz8Yb1SbuLKmByLhVh2zezn7txfhMT
H5MYYxU6TsI7leVHogt2QnNrhLB9BzPEbVmz4sf0j2XAiL5v4XcLtf6ygIJjtiD+BTjgjw4TtG9M
5i95ePtphh7N6OenXMDAn/2JjJ3e1F+5X9Ft3ovWEKXmUeHUCM0Gw1O2wBxHkXLhTGBxgjEKalkg
J9RQMI+wFB3OKtTl82WzIq/jZ3PgnCUsCtR/jQAaxCxy9m2gvCIsPx+7mPmR5XMXXELAcHk/lA9d
1wBGOvZRYJAmmkr7Ar0WRbTtrNZkb6Hg2OAGNk0N7G6WuvI/Rb6Y0+zrwl01GrfNAzg9LWe0+mVv
v1JJMcFIu41TjXkHlrPiQdjjae5Jf0cUXOhuOC/OLtdp+cHfZOVRtul1kfch6KKBKV2ozT/mvZoU
d8yyYVnVHgsRJlKvTU0YOhWZPsc0Bnl4pGQyFdd6w4lkXwZuYPoRJ+LSgQpbud2EnWlWw/ppdYCr
b4qgLZ1HHT02Ez5nxsk6ZAFvmwdPhKmiZfYM5bmcC2oyZHP4Lm7ajqIuXf+gdS1hWg2TmbcHqHls
clG9URK4HRNucNc71WBUQtfjxoBe+MDqW3Psu6Pe6AFYeuI9NppAsh/ipw6f1LEVLO93+jiKuIP5
G0BlAVX8h0Sr6fBpNJvEEuTyVHeeTZotDyiWRfKIxMz27ON86kPHz6WFMNX4mm75sadd44LFp8ib
BHAhsXTi31meJle6xfIadjyfM1wAuO433JPWzB17P9UtLydwS2bbjBuBX3+XGXPUcYUbiDmQ2SWw
2LeHRjRg/TychdvMm+z4l42C9A63v3GzVd8fKxm2EG0ynrc8juK+4NA2sBMm4oOJ6hjBBRnjJUsE
3TwuFCsqEvQawudNC0Ig0zEggSP66oONo9rAvGzceQP6qmnS0UYIcRI3gEJMbU9fav0Audj5EooH
UyNQxVvA3gVEFEm0vgeuwedBv+Xa3ZKOzkLbjmq3TG3sllwAiLeev4oW1BkKxZ6H/9rgZTuotb9X
Q/mQPxnsTzdAei1TumSSlX6UQ/HSvvlCFv245nlzXXgIsNJ+MFRDG+zmBXJyBJu/IxgiOIFtvEP9
RauvE1gc7cTwzOJbr9Dh+C6G3EQRQXa2C+uC+B4AHNXHr5J6uJy4vGL1Ai2fTp49g201Bf3j8UcM
/VTyfjhLRS09bmGYSxhgBH3S+qtbuiJPY3MD5MEprCwKlLgOeTxHBOsxQz7rY4NpoynWOl3USDeR
vGbmmo57eO53F/+ltU/7l/wQNpqq35UCUlSRe4ySTpx19CozRJRpaDWPHuDduE8xUcFOOqigrQhH
PzQEZ+fq8FPRVyCkD+x827cnkDHjk/ROB4mMQ0OqWYzSlEEjolXFYfFZrAZWGzpCDaXIcQU8m5Rt
hvFovnyr8lWzoJQk2YLt5ck2w6wfYZfM8qT4rr64KW+MHzpVFneO3RW5sHHSAReYELg9VoF+EKKn
4HMwRUQV9HrajOmV4BKu3rp+Zxa/5VBD4Fs0VSoifPXdffQ+ctoQL9ZmcPh4zMFP8FFCsyBluCqX
lqLeHUaFny4XdckeI4M6T6/pmMi7iRD6kSkLU8VI0IulvXkAUle6uk2lb9mrlOW6nn6gxWDb6+eI
UcxckoAG6eSYFIzIi3eyMKySFKdM6mMiVWwEkKQAuvb+Mss88FXVY19FN1GlqbSLaCjqpe2vbEHv
aUWsxQdR6J5V2Yx5d0XqQ+7NzOxxp+bdrHk1YY/NXniyEnqebcr2EDSIkLTLA/Uklp9yGuaJ1JLz
+60o1WMRC+I9OTSk1EZmErAe7tT0MazVHl3pa04JfZco7W+8HOL482tifAHih27bQJXFtg2iXz9F
3S7CilrRQKMqlunshtSfvmpv4Zmt6j2WjQ7TH5zveD32AwauWTH4USXky1yT+6jV36l5Rh+OngY3
iaSqTp0lyY8ulF7CcdcaqcY8+AqQoVUXPJrrQNBtDwZyy2p0sZNCQf7LE0PcDr6d2vnl9u7PjP5E
W5HuxJRoiP92KLCK8rKL6JDxP/cWbWL9DArULPSXcAvHi3sKupF6E5xoZ2CXR12N6gNcKZ2SRJrZ
DJA/jJGl7fYafFv/uW5wfBmRd78n0wqin27rO0G3ucSJhZrn2JIHVandlnjHaPuERx8x0Lulzd/7
1bPtqji4k1haX2yR7/6AG+QbKtMO6K/bYKnF+E8HLnxcb6HdNsnOQG1b4wu1dHyCNUgPLe19e7XO
n6NJq2xgoaVmYVikN5UBCVi1f6nvM/GHDOflcZvOTqxEyaTIMahAAOCpF8+6nm3Xq7iyfEJgn37N
6XqLLfihduakM2hWnhq3VIxGb5Ci6tLmAY4P+3Aw+wAvmrB0F2FSDOibx4HXn4tnW+QFulIcwWSM
z4mkszJb0u9jveD5PBIdsqVq8fVqtkGAxIPwdY0loaGiAMRZTuHbtqZ0t6eARzAYwYWUw7Ej8w1j
gL/Rc+kdKU2AmFX79EUMyIhryM/5c2sxSFGcTnwFv+PnUSg/T9/nCL7mUseszVuG9pq67vaGjZN8
oJpctQ6zRMAtIEvXiAG15kd3B1JGlzykoYVftuKhP6gd/CUq+zl0TCF8g6SUhW5wur3nYlLEaplK
bIl6Wf44NW6WAxB6VhtGUMw/ZevSCcfr3MxyLFnFz9FQCw6lBJy+Rjf1WPmCijH4yR4xI45Iqx9m
O63bvh/iK64LCReolVTm5VHEfqRFS/8ZP+t6lBUDhn1mHfhTtpi0uX7a9aTAIKwRNXmSD1Pm/o/E
hYMW+/kyC6LF3fYAmmJ3TEPHmSGkIYpjFz24WyZYSYOQ7meNIDBvrqBvgah3aah2OUEhLsquwiWO
bCaLWWq/CUB75Vrb4Y+n5UqNYkTWSGQ3UPhfakQu9wANWIkPPW2QJ6wkEkNN89IXKZ0RSoXuLGGl
eCGNZ0gxAHMvsT2fARdocCT1wkemP4hnDtyirm6ehQOWeqp5CwoM4T/bZexiSMZN8g4Mb3IGuCBU
tXOr38samxGm1o8SpVeqAS9GwS6nO/IwDeYGxwH1K4jT4J9lU7huI7TvTZ6LoQR4xPoTYGFkCUCy
WGTu1OHSZ1iKX1pazWKbq39dGYdTagZNqqqzfDQ5PgsNxqoUV7nWR6PKSFKyUN44fVh1gnT3CU5s
DwoMp+HCC6a8vdNRjF6j8yvZAnFNYeBUM4VVYaxJUSocjeez1wiwB83hDXRFllGbMrnFquGUuI4W
CR+D67yi4Bqn8Lb8OlfKz+WQhjSsTBGpINeO4ViM/q70/EXQJIuzVyz18PfD7qekkiNKwqKI8x9m
+OnTRRfBN3S+zPBZaSHXTWfXH/O7mwwRflN3YSGz29O93NFJ5tA2IgxFUYPG+9JPA9SvH9rpV/H2
iO2SGLDpWY4VQyK47BMJS1LGXjBFMneGjKD/cD/I+bBYRc646uUPr5uiolfwFyzAE3zbHf+Zlr+N
xjnQhMFuCeZSlxFkaVB4hYY2qQMRBBs/5YiaTRYfUaj9ovSAC2btANox7pDDStBYzNuyp03XHTkF
fGVzLnpt14VlMaKNOswg2SWVDPmPwrTm+7CL+1M0+UyDtGjDevo9WZSvlTwvafICZUD703cSjZOY
USmvRkQyzTh7z3uNmCf1dhu9ivFGtcjmB7+tmcpKNgFZD9WuI9QKIn2ELyX/4jBqpWEkggbIQkt+
Bnjv051r0k1bqkA1VMiyLUx7GQR/Y/2NHfNz43qUwrGzadAkNOz84dLoWBFRI/11T9/YnyEIj2Du
8jYReCQcDznVOcFGrri0TkkG7fc4YmEgpGpa5xY/uO6HpobSmyXijUVg6N7xm/wqB4o+k8ESKW4H
p5dBUvPkOArSnVjzDFpPAPgpUi93jF9jaJ49GcC+a0Iggt12fMEQqGmTfrnsYw0ADf5I06N0zOQc
4QSSlyDm/kzelaSDrZ/Tb+uYr2UFSLPBL5jPHPQwGjd4Ky/ZCjXJeJyAJQm3pJUSNa4gJTM5txeG
OVhFs2/BuyS7yG4eIcCs6l/p9mAJa6uz+C+Ru1Ex+pidAhUM8dgl3rmYQcCdc1rSI+vpExzd2456
zXsmHIfb97QMHDFa4qZHx2PcSzxxV3F1a2SdvRILpYycnyBWuRvDArbw/DjtSpyHIZunYiwGmw+H
6gelZYP0or/6sXrEQ+7Ig6+sfBfrRrpMA3O19Wnv0mLzB0w6EkWtB70eW+h14400XTbR0XyebEsZ
Vd6J5iK/kTC0FHV3fXmnZ7Yxm9WpqYnrOXFAVibbKs3TxLb8eOdeOSIWyxuUHi4Pt/Dh7FFJ9jgy
y5PymtnPVBNpgo0YFFGVg5n6oNR7+r3scze6MztnNI1ngMdRySnlJURwDRkkvGfzIAY76Iv5fHA/
Ga1yxNG9RGZZdONghpBIxmvDPuuCTtuqQx/BJPk52wcsTDQjVDqeApHUhMj5AUoOnN+4oByYMti/
c3MW5ZO28z3iDddrWvLATMBxFbr5xcbccZS6Y03tpP0nY6387fjZMQ5NJ3PvGtiVPHynyrHvnmgn
FZVGvpa3K++KJPQvY9fW5vFA/HVptQjA+B15oa6ZOiRGbCXdFq7xUdEXVbUATbFcmII1CjIQdLRy
ScZVpC+enn8Wxr3JgqcoRnJ2XpLTMWSJ9BwPt/C/pT/7mLyEkNHadQlHAtyuSzkZgRi5AI+eheRm
cU7E+dLJEXP94Kn2pfcHYd1nrAusTSZOk2ao7oBWYweKDwDj7/Ob2W7yPWQU8rMkaDx275kdXdf5
GEeiCDKcBst7y2AdiG6OPvpaDs5gxOqCKMU6l5mlmQPn237iNy4B0uUzehezqEhthcow+Jm+bprB
J0BmqlFpevFTcey4ABjtiimIJfNtidt1j2o7q2z5GY5Exx9GN0Jj0rL+ft2pnE/HYGUhl3MNpccT
kJ29LWmAbLTaO6rxb/rhGtGRLQWLtY4BkDUzZXyvZf62KmNGQsaPQXv6DQPVBRyAZc/0PUkaa15y
7d2biWeilZlr+UsI5X+dMQFZTzBL12OprLfX7MRFXtLZ9gGGNRRzoN8RF+/webSUaJeYzHuTuUPm
csMrZrnDfSWeuYpSSdHRRRC+TLyLe6WI2SwE3r3ffsyZXjA182MY54++ImMwzzEn+fgvgAH0Fk2Y
SNGmAOrVXleStcJJ5kVlRkJFJwHNxeR2mkrHF4WMXr0p67oXb3pkLErCjs0jBmpR4nbsbgLt2Tb4
yhcqhbCgfYzj6rvR6QQ7z0xOsZSPsN49e/0kAes0NNgCruW7Sp4aNV10EJNSp5h10zO105StYHBI
L5Q8jHRdaOA6vpD7dqLP9H5u+hoexvYT8Y7akSnFKPbkgGYJx9w4RWZ6zMYNyp+e2kE+Y+3ZDwBy
vq6jcaJRBLwatiRqCCdSwi4S3dhMdkoK96ckloD/2YFrJzbpvZ5rQNJm6liCFUDS0PLKCj8eVhgA
dgjvDA85gnmab4tvIe4lf0p2fsroXHXoGy+0mvAmjqk9P9pi3lSO9lyB6Md8odIw/SrFfKjkTPpY
+Pycf4pBQskaDB9HIS/5aiDCo99TAQPPVZDY/DmXsslemKAkzuopnJSuLFmpx6oUgfYpaH2PTSnJ
S23+sMZZG1fHL1EMT6ycvu0BFbdkHU4Z53BQZhS6LC1vZQsVaSg2FgIRCVJHepJ3DMjqGpMUvUMQ
U9mKMKZBNoqCAL2OrjzA7E5EKCW+RIiAFFEQC+lYYu1URA2Qc7dJnro/YjB7PVqC6K9Z0B24LOGa
455KVN3/99SVv9oqorLK2l+7IXgJIsPAb8xJO8795hhSBOo0M1fE5dmtWLcV16NX+KI238YyfPjv
fqEnykVn4FU4hpzB1BqTo/ULW8DtZAM16Sn1FcrQisQPiRouR2uDtE/MncyLNXkVccPcpcvDCSdv
HPkbsephh0Ju4xFRAyXU+rp7xQ1tdhzWXhjF2tx92kg8Jkaq8+SSp+kcH46TpyR1AH57EJ6StCyZ
u2vr9n8XDRfK4PosgGMB5w1Y9/UNeDapA5QbVxujZTKJu15g69xNhfwxujMz+gAdEMNEUjmzDtXm
gAPyyVXGyvmyHeUz1njHDsSQZC1EKITdwrfrlxCTRBpGRAmHSPJTG7ij6wlStNvkkpFyV7PBGHXc
zxruNLgDFU6guVjtiAKP1nEA0BJ/AAUBL11HG8trJjZ5teanRelyJAxpUeN1VDAMANeHMin/1UZ3
4z9gUcu9jbIv1eoylHVUdAVB2QOhTs6tkQxEljOSxsgNzfAgUypOk6mByGCwq4FMsLE5PBlAA214
JdemGuCs8SfES4d4l7wda85RkNtF+C+tga8o0ty9V6vbCoHs01SjgrZTyFS2rNxdQd/BpdUKzgL8
A4c0dIckobVewNhbgcEU5lqhbTQccIy8wemm/Uqm7wvM7HfbvCRfG/ub3CQxcYVjbsZKENHlOBDR
LGIUJRynKeg9/b9GxIG6ltWadqvDBcMPfObYFMBYKO9OQrQCNn1YlKFpVebs+J4/XKazgP5JflzV
Cv7cRZPgJtThYeRPwUNWo9ohpzWzLkaHz3XZK7HRWuG2jXZ0d2YGM1J9L2DEGHUsSjoq95BD4Lop
iMguDexezz1XHJ7Axn3BXHJYUGmqp+Vqw1ifPVg8FL47ViTKUDqDfdvkD4nCNBFg86yo6YGfv+LA
W1U+ZmwmB+H0x4ra+hPhWqUgyRjnlaEPw4Je+0wh0AxsjfiRkIhaAb0SXy6w15/v6QvnwArepi/e
62Jbvat3dbjnZFvAn5RLEC51AP1x+np9e724INHJ9yWLimF5KbSkhPJp2tx+egw9Bj5oD9o2RQ4P
rOcXdMQxOnToJMHv5ffozrveegKPTTDHVLnq6kIIRLovMejOL5dzA3EzvY1qRnDT5JcppVRAeto6
r4UGHgPpEoQBV/xNQVOYkaSOGjy3LcSsjwAcSoFTsj57hj2uvJWCJf2kPyM+EUP/yCTC9IWzeyNW
ONobyxIZlrjq7c+pMk5f42MwO6YXX90WPIKhqS7KQIbr4utHp9QwNNUbHck8bKB9Ptbmpltwmnof
kHKm/ID9j2+xhSUGKpAm7yYu3YURLH4qbM1dBKvGzFZNSI8yMXEihilYMn7D+zAsnnszjiWpchbW
005nUwAnVGBmnEaLwDFY8iX5iUbfBqv/fVjPB1uBPszWwK36D8sa0zcaPt23ar0bcNao6tTjwdpD
tiphr2qcSEls6e9kUYceH7NHvlWEpGkO3emiffn7YAbHxvRWkxDkfgwhxQsUMC50Gz6RReLRk0ER
F0nXVB9TQHWomIsJGNdY1KfX30CroQSRVmNAgC6zdcfLxy26jktulWucpqyp0Reemd4TE9/gCxTc
q8TmnksPpaTJOgWNLGnq9ikIG18SMRYgiapXtBTHq6infdh+knwikGown5/lvICDESR/6O5bHQ4D
jPc2W5sEOjf8ZRwjXnIF/lDAsPLw0uCN9WZX9XQj2d8ngTyqdRjFoWn/nyJ8taYv0Iv9unR9J2Cg
XbI9UPzJCJbhJAOl4U0u+MqgDWhaxXhsjdZ3mpsJ4h8x0DsV/9S+i8JgAxuVude2gUdTIe4yisgT
k4CP+YEFfsDhdoKk5ci7Y10+XDJjQH59CcKKednEvRMo24hld3xozbCOhNqOMs+LY2yeHt5mNAAW
7QsClfojTzbgYHYb89wDZvz+NGKtDkUROWfUrUMSP/y+kpSjoUuiGWO6tutUiWkVKLQrEYE1SpKh
ZcFAkk/twKfz2AdfPQKWKuzXOsGkYk11UJR0vZIxM73ULMnVCr0y92P2v63zQmiRHMJp7PURSJEY
PjedrxP+TwdISu3ODZlWT4zLuil9+Sw3HINKqhK0tdCIvfV0mRl2Q0rdtrJyS0YxRVkQlSQhmnM6
Cxp6B4aw8+NCcpaiiX8TlwXdUJzwfYZZoLxtpiKIPoct+0Bw6Tv7N+IwuJUQiAZ53Uhw85ON4cBp
tK1NLzJq59mUbaPW9lHawQxfaAjaUyoLOKtGX3I9AqgR1nd++FYGdmtvTQrkpuH0hHbbTBUm+wP5
g4dq3G2qDWPl9GFCVN8/BTdpbzvs9nDxiAJUyakOb/OHAMdHe021v8vSKPzY0AjlXoFaUBshGMdr
CGZdRs9t47nAa5PCGa40s5PNtDIf95hBE269YRPrqCZ09Zs1epg63oVlh37nEr4b+PTnnG0KWalE
Bp3PtZ7a5zfy9Mlco8Y5dQkkFfosLLlEDF0hGXzjdliB8MS1/wjW1iKEj+TPULwwkyQ7+p6bsWgb
YfvwXk4fihT4KM7fARf8FXcrDl5Doy4ZCtBpTR6AZXGBeyCu+fWA5Tr8+LbJiku99AxgZitonQbI
z5LLWwBitx4pk7UaTbSCbrDAqOxijh4xdkJ4bzriWELezhbQRL2/mpLmYUYCFYUB0Ww+bFWpZmkG
KVZvSUG3ZCULF0sbOQTbNSxBaCnL1MCdxBTF2H++ztzYU1McUcFuzZqYOqiaLoDKSLPDgIV5GK5Y
J6nRleGeOBItMtYSxj29LFRLWrAMxxVjNxF1xJUWr3WPgf65y/wc1isYP5dNBuzpLJKH0QI7kWNx
jKYnBHXtb5jNWKP6L8i/B+fA0ROqBZxhR76jEE/KTEsKvZ/k6quAUiNFLAgSmlC6gLzyXVzUO9ru
5O7cA82BJFzt4tnpj7/z2KL2DCBoqUhPSBueLNWOHRkkrb9FkXTTAusGyYr0nynrKguqvR9y5b6p
NtV3wQOlZJzftjvMDqAE5GDYcGMbd+KSevob4B8KXzsajpgf3hUelLxZ7Ceo9LS1Ah6439hGx5Ut
kUDZX+YGPPfXW4LJ6kfcAZzZXjd7cjWaLUo5HxwCaNarc0A+PE7RBeMCiQE7AWHcvOn4upL5RccA
3IkWm6/wyJEtHUCBcQtzcgef0p1vzIYXj+bf2nvPoVruqtqcQlbmc6IcswRYCQ66JqdsKsLHSBHl
4V2YNTVdW8ZaUk3ZAgsZydnMsnclABJ5gOGC4E19SVk5fucvBX5as/BhiaAICNrbWPR8KsK4+Vw9
BB79suIiN+w9wqvpT7f4RA7xzbzkihN2IRrqUizADnlNF+rArZ8uTzvaOVKUIFFslVP8hAH4rxOQ
R6fldic0q1ErfuAoA718FaW9dlyPpISux7f4o/baGs0Sn0w24fQGv0KHG1R2RGYtIozfvxc93Q6P
WtmauZ1CXxnwnXavWYcq8490P/0eaHbXK8rvP0bl4l6d96CxijwWV5wwRiOPyZoCjsoaPLgj1JM+
bgZ54iLE84CSsY3nDhezdGoQiWfAouevmCmzspdGb8iLHNYIq/9RSn6uF238Ce7PfpN9ZVcj8STZ
zYkZKNNgnDsVhidBV47N/9TdvW6qE0HV/60r9j2F/6z7W5L9BySZ0cq/5kbNOqqIIoEsihuEdKOb
HacGCbdj1QjZ3zMeJIIbfFR2q98RArZV5osA+X0Y2MDnSOEdgc56nPxhEOOjvP/Tl633fpyvPwmG
ndMs73zHWHQyMEZEnej/N4RVQn0LpDZPZG9NT+2SK+ne64C57cTcLyl2r32UBVUqp2GjK9PMnF81
0kBxwvHBABwP3kZL/qvxbWetaJ6eT4WGlZOR6JrtvFOwbY4QO2Rp3xEmYTR58ROQs5tZZh5yO+uj
i5LTcH1kFkxsvABaWWq1hMjIq6yphVSmcDQW90y04I4QbbfK6S/2PnqTygG4GlR5NNJUJeI89wGT
jxkmFXpdy+IRzCraCA7MlkPAy5578g+JxrRa9WhZYexp+MEg1+5+DJatEBIuJOlvVZeewVusLVrB
132Ctw31ajnw1bySGf49dwz344kJbZEYuVokV8FWKHOuurYvt1fR4mUo+wEN+oeZYuOzY/FgLpaq
PjKUXbX7tpeIv7h2Hs3xRxyfEc4bnx+1EwYgvc3mLJVwPkcjKQmoC84hEZkBorpaQyRPinANCUWZ
fiVm4+Hs7BN8zuUwBMgCsIIxb8oLyBS7NLELVu996UbcTA2THLMOqhDbYFpcdwPtZo/+AX1wfXKU
9HwRNLiwy514bylU34Rf0/TuZr8H9TpuIP2qnDYby/15VlYhMX1wXG4Lbbsa8aNXFcNAKQ8u+CcV
jtDPtrAxs5Sb3sqUAqXQI4e6F1e+IobS1nybprdYHt1/CiSVFVxAW1uG+dUjSC+eJ+tepm/1ZrVL
5enGvCxp7LWRoYgNSTg/0LKMV2OUa0OtIljhFZUgKgrSHW2iIZhG6yZC+Cg/RWLdyDNQQg3EKEf4
EF/HfG8W7m4/gPVhjPQg1dksOYsRjiKV6AsW6fYe+K67pYOYjaQ4L7o1YFJ4QY37EZimSGjLIdHF
v9TlRlqnunf7z8zMzzL09GhpkUxR7L3z8+WmWO1nTHaWunCj0D4Tv5enHtBbXrbdMvaYFb3UYk5S
iuoK9XIJ04FDkBMkxwpN5LQYTS6UGrkQwSgW9eW+NYWF8fgp/vBAQXGEEMv7lHFpRwCv3eIG1sS1
wiV+4Iu7E2W2Cawy7NGNHntzqgE/Sx3Y+Tsr2njfpibDz54x81wJTnLJLqbbEueBJkT8OY49L/mF
Sdw3fMbltQ78flNCK+eUPbpab3mbBuaNEB9MkUD2Vj58x3erJZL8Nqpkl90FpZ1Qbl+ffE6vBJKm
pwtaSzL7i1IwIs4ssDu5jyTXtg1NsrtyYr506ZNNoxQa+dZ8sPtqhm6R8PwPdA0avRl6ZfrJuUw9
Bm3+RPimOrstBplGyuriFDF4WdodWRxlwv02MTpQ8GYDE1vJ7mXuSTLTdaZ9MGdP4q9fl0vCou22
Aj+FbGG/RdVWV8OGLUXGJp1/ipt6smX/xtsrP9vrO/Kp9D9JoVUmBnahZMqim8CIXRxTdAtEILiY
+eBrtrYVRBLYHypWBem7Ft75Log9bboBSyZ02xQiBPkpGQMSsbfFuBJn6pUtXjdm+4l61wzyJcQu
Vuf8tu9HCPwkxTulBKk2NLLuHy45xaED+93BZTH34iZzyedLXLj52FeRtFDqeJEeMqxkDRWTeqly
xWmgarVjGWWMm3HtJC/NG9lXXyWSpT8bMcEA5uqedMfdgB5rcgES0Q9fEIOpmMu0bLte2jjgf19q
7A/wF7k0yF9v/mSk1eT8CzXIK1rAAAFlul8qAPMn5TsBX/ZXq6ydchWnC6/F0iEtSsHcEWE6kr7k
tKIFT4rveShUwQNaQlgjlEHveBZJPB7EuikYUkYOIHrLhz9CshhW8/ShgFcrqsPLg/0NhYz/d7RQ
Hd0gi5u6p1ingi9I/xY46rDmKgB9MdyB4ZioeqL9r4UHVqXvliX0ki3kIvkJzFWV/rGbo6F6Eibb
on69dbjl50cy5HGsbV7kVj0oSlPvxVZneVyEjykvgxDAfUk2c0cKb0g22DdFPmsreYv8pBIqQNrF
KMDkJA9/6IvBtkq4SbmFAz4c8GEynShXyXwGP6Qazd5vwvfz+7hq3TeZTamKBAZZg4tfvwaUnyGK
NjJLBnBsTvKVns4lLTwxG/UFn5MbgE6VdMPhlp7p/faeGmOzpAJGwYgjQOrXyaZpQmSdHVTsg2Qp
JuZiiMcAKJU2wsnp/Rb+hPxubJUBPz62l5urvAuQc8xHAudjbb6Yi7edoysvDBEmKPpSS4BVpBks
OBdoS7W09+r4Ct/0sD/6a3sIXYzAE151xnI3eg9MMlv+uc6xLAFg9XzHmXFsefqBza+MwRTeV7Qr
0F8VjlEzBmJA4TfblYcTR2xcaTvd5jgNfwZPv5BbV9tn4BrHrs8XwQ8Wb1wvvkpHdPASZw/jy4Fd
42ldmwCtWG5srlwPalvl/JnSpuPsys0SNC8FunkUsUgsATsmBo49lNbljmPtavx6TP7nEWA0jKEq
f8VZq7vKgfo0+lNu8c+c9QmDxiQyQs4VJvpteQrYlJMaD4DeUwHt8GLkEROYwxPIhVDgMQvBr8Wa
d3j3mf1dDR5STofFWzrVxqdTuO2xFVdG/qRNyRFBQXKqgAC/RqgvctKXcNGeHmsnLQ3aW6l12rzH
QIigareWnZmnCDdJSclYPSJN0b7ilKe6/c33FtjOMLLOVk1L+sMxg0S0qWN8WN3m9I59Rwta0+0j
50biOXsKRUE84ba3RSVuc9wdvYkkeSdoriFPblHHSB/hKkw/RIX/Mkw5dDVFQO0bHdP5gk7AZQrm
yFEuU7OqUsbw2KOKZiKTRVUdcrrqnU6iuk/lbC9QGlrLpAlpokAgfvdM1MjX2aeZ2gntJQTG+cdP
ni4jyMB12AXC8UQKo1AVsmvuvvE56R7vaTWmaZhcjBAAXFO6Gu8kYxGRObIzm5lknxI1fX7wlai6
rQQRyoW51SUwJkLaPHEdz6xLSwHGQo09DjVMEOsRCh7yP8LS/zet3qKwi4mH1u5V08MlWr9AcK6K
hcXr0voLJMDxrNyKJWLEZGcHrgsEiOi6PFyxYjPURfr0Acg2aY4brstM+suXAEjW70OV/cIAA9wK
H80FfrtBmC3mIZt6oV1zGbd5gnyxH2jFwpcMyf1LkFtf7uZyfR5KhukqIdJcPGFs3KT/zdPvHwJ/
3Oq0Z6w74uy2D+LvkRplq3cw7E+xn0jrGH/8J5m2U3I7oMr5EaEv8QOL5eYx9MgQx0RRJb4EQ8OA
SrnG7oYhaM6PqdVjN2vnybbL10Yq1fEY/7patB20/76xK8ywFcplNE8srS2efGhfj+xfmzYcUaDj
V3e6r1tmMFdnEJv3rGwv8V0Chp86F7RmBQNgdSuog34cCnhHcK2kC16lLkosqRHx/pcVkf3g/bJD
YI4PI+j74hCQ0hUQzhui51F14vDvmWp4Dvpipc3E5iZ4l2/1474dcANbM70owoNEuMwc5KIbCDmI
OaaGESkU+kG89Dvzgf3HLW8Ly4ZgLmBJyDWuWyXJ7qErnk23+htZKXAaP8PgQqDOpHGTP3vZ8a5/
+aUO9WdJmGX/GPZYuQ7tGkAYKIjk9/jfUifmOdMdcDQ+HkukM4YdaG+2OBp7lxKKNR57Cnw0lYDb
bvRYRRlwk6lGLBaKS2hmJSjy0BH8uMejIgW8yLSouvT8yiOFCIhWHZhK9pa3uefW/6tFtHHMshBs
CP4RtQSiKnFwcVho1p27lr3hwl69hItFva4x6C4RrpBWH6HiX393kyL6Eql4i9Ei0VccQFOll7lp
hcK6+oEgg6bHrB2qhCqyXl3BPWI1DNjkI8M6OflkQQ8M89rgESYaFCK4UObvONmyOvH8nGu9Vptx
g/m8jMax8kUXPNegeYP/OAOLMQ0S6ZSS7PlGrt/498c4N3hssW0EEFQXJW9IkjTSvY6sOCvGG8fh
W1k8Hsiaf7o7CAi5xt4S0pyPWXfB7OAcu0VdLFXi5KfqUkC6BRNcDrjlfLDCBSdOuc6ZXrIFmG8U
LBohEYdxloQkX+orGd0ysOeOJZ4udo5yYdSykzifX91cQKL+fVTNJ68H0Eexe3ZAdKek63wCAz9/
x//qNSYrMyXGKlXdNnWCSNlSvXOnvL7kDwZg7ewXkLk+86FZG+ou2vCR57STtw4oYJ7SCWokuM+2
pFL4K+wvCpOGI1UA9dEexbC1mP0R3Wx4OLmae+XcntEN/+B0oRrz8TwWlBq25mE3rN2LyK9lo7aa
DS4xJhymOX8/FnWqaASqu9DOpmDOITXaOgQgUhufIB+8/Om/wJFVgoQGiUEL7AYRNm5a1qFpvKbw
ZpKDAg2iDuTRSSHAOoOGHMoaA+R0gW880Wu8y0SJ1AflpQIA2Ne7TH4UJDVqCu6migXpyZVJMQUo
6wR0nu+MyOu7yAFxcvfv+QkBRdqeJdnKlyRmwhKMr7+z1zMhbpdghSNj/fpQgYHhpMwFDs7KFdg4
I15MnQJ1jhZ75Zvs0oZJxKKLUu6wJQNoW7+neY8I7M82TKNRzv/vhx7iSRDWyUWB0AWrD/Fdaabu
6e+wW1qiXPg74lk6o3wtCDE+a0hFMIyFAzY/U3IFb3bFxMjjtHLnkNsF66/K4n1XTRilpXZwcCRl
OQK2MP4HIEy3jVcF60T31vQ0YV4L1XX4ufeQt6nEh6mi6a3ZupHkkptf6dmAuoDSmhLU7NeB7uaR
hbx/wV8DYKPabzUqeQYwjQYllCmYznmfOBuG53RG4yl8CfZRmpPGPG58zpjD3PjPUL7Y5iVolSf4
ulAVub8TEbGpOHehvOC1XaCJCuCw0wit8OVpdvnv2lDIxd6ExFJUyJuF+m2YzutI6FvrsZTuTghE
0yuETpoZ4MkgioQ4L9QjOMolgqWThRSC2D3VY/NCB3YJ24xG1rr5az9oaNqEibqzOfBgW8XCxP8v
qwsKTWKqdxMZA3FMf9p3Dp3mjYOF+5JHxXXG9FkeIHJTQQE3fOS7yVDwjPFW9Zwf3LveB4/oVwgq
uZpRxm2DK1OJ3IJgX1t4ybmQiPmRYx0DfCA/G1mXr5Q2t+kdlVRa1QdJ4DPDaeX5rb4L4OKJt0uu
Lov1rDCoYnfV0nqwRQeiDOJGhX33xhO2R9ywuCk+Bvs21BOyO8vMX34/H+kWtLN9mmhYOmPaojvl
hhc4/WGHll9t+XL6kjIif7bLRn94SbM7753Svf6YLl6oyJ8kBuPqWyXET4JOjJbCrtPy2TAikGFe
yCG1MR12bpVHW2BnpVewfDqv3TAjGi2Qxolr6o0VQ+0Yczr7Pqmx4nXVW8YJO4X9blbsHbbpyakN
1gVdLRFm2Q/RPOf7nHJUA8EN8uC3WQZeMK4QLeiU8ZRrfKC9tohg9Gs4iXxCuywjFzSV4YWLmMfW
PthGOtoHTn9sw04c06Ni+qXr4izG3rKwpBZqUGrSeiYbrterzWnajrwiIcLaIQ42AzSYdJQg6yEe
IJnNDuWmYPa59q1bJOQs0PRyRmmzKqdwRzX5yHzeHrtCva+PaiXUlBV3uTFSuYpIU2LzrGHo8eWC
8YSDvC9QX6Nwl//TzKzUJukUTNjhZMrwMqWjXLrNwOf3yZB6sv1fjMyylp9X1vhEikHDYTKNRjCa
DXkk8QT4CjxRWZ5u+jmXHw/GItCAOHjszS0KtIx1TspOnz44BBw0DubOUGLy8NfDgpYvKLscClrI
y0sLRKqrKqRk3F+4yyt5j7QzgCyKdUspkLGCVzoNNeNv5/4RUNEf9majigk+NpHFSgpcJ9KIMvHp
YLNyUYuRkSTR4iAk4bysttGMnn+0rpIGEoYJfrd7fqXvXaLPw4QRHVs3wvSjJaI3FQwBXInvtoMO
VkretRjW87XITiuPg5UzvnQ/Z2NMaNJuKPwrrweiyloINcBOFVZi4T0Lq+lVlqMXC/gY6blNZWZE
/ECTVZvziiihGykuMts/USQyAFBrVbURoO3L5/nbO9Vbap0aJ/0U4leI0yCnLYWhGP617zUjl9Oi
ANH3x0fETCQO5k71J+6aV7YIZ+Ua7shY1Wq2nyARuan0vPINh0AQPoAl6afVbWKevpkTeTx8QFHF
B9vtrR+GktgeytP1lpaHZNdjdAQA0m34jJ93KRLe0JlxBL6mlpIoXvDHxdPyCBi8CYZ9U0uCuUeB
NO2RkfPpPj9JeSsmQL2+FDNz3z9yoeDKAwswIjFyQXMzav/3ZUXK1/Nb6iaKJVtr0Hxe5D0uOa0y
JC4z5RjS0UDssx7qrNZuPFXtl8hBCry8vSyxkG8RsHKtbx6w/uVuMtdS7TAUMGekFwISaKiAQFEa
fNiohubz5c7koqXVD7V0BfZeXZv/vu/fl/HfiUnBQs68PjS/M3xsXhLZj2aqjuU29+YGtHcscPtS
L8WnsUhmo8seM22+pVnN44nnZAfzavjr+PsuGEThpQ5tpQxtJKtdo/ooSX8XIIcQ2RBuIUAdR7er
AI8mMvI3ttwCCc3pjjhErY0eUNllxfrnF1Uq2F/ax6G1zMOmB59b0hx96vA0iYnj1EJjV3Ny+J2E
Op3HBmNC2K4rxGvpL+Kah+4bP+viOwiJE9Fi8skj19n21V3gPI7CEmQSwAKV1sKlKeN07V0qQBjR
8QrdVTJEwah85Fad/1J7mwTBslG7roOSBs2a3QuVXTy/GNKqVUhJjTVt8t4DG3Ye/mR+84IJ5kPe
0EKtOgkL5yWXWusY212VnZIKoABnjgP/wAAuCa1uismBM5ggQ5mF1vMxslHvp/jkgKGlOM2na0RA
bH/0jFXjwx5PiQ5nyBD491U7QVkSqJLcjGF/zYH6BQMnoo+qUnsas0Ju1KZlrKiHaGyFnn9tCeaB
+gW/bkjVbOl1wd8nFtdlwKogt1fKw98lxf+3VG9wLcrzF+aKDYEKP8ajBUcaIDj9gbXltnWRmJVU
0NQodjAmWWniAIjYUl5c/055BaIwVlwjkwjlhdX5F47Wvs3yjdzlRGOwpw4pKit4bTEPer7/z3bD
fMRFaODQxTJFiOFVlvr5foE7OkU6EjkwCL8Kz/4qvVknMCHJdCFR9sAQVElj1nhI33y8+pAeQ8q3
vpRKdGH8E89KrrvF34tCyT+ADr3SvshTcSZ/N1jwmqberszDQF1Ku628NNH2Cw1U/bPMr1nmO2BL
54LfKW2UnGg5+ygMQ8Gc+Blhwb6X4tGzolm5Zna520N1VuM7Ubh/NS4A7STqjVTDnT9+hmJOY9Yq
UAqxz/dkq0cM7W5+ZgJN38otcWsM2yvaejcgvjonJOygtqwcF/mxN6Jakv9QaiqQeT/AppKzgGlU
KETlk42IhXKqmJcyCOSLimMseLqh2m6hKWgBh5Hed7K718a/YLHBJRX8/mlye+GaQDhcjYNOh1uU
CaNhGLHh/lM5ax/Ny0Uo9XgVlCJZaln+kPWi1gegTR9cmxKmaLvVgERwC/KKrbTtZWKD7yGIv/r2
GAQzi9LonPbOWxoVXiMOTViau+gDvj8gDV89s3Bw3lk9fVawEaUhbD1a3tcI5TJv2aLHeRvcMUtv
3L0G83iVWij8lGk2ApjAN7dC5TcIeZGrv6R25Gn+mRYJnelRSLanANX/t1iWkxboxEYIWpzONequ
AbsjVGOHEtvMtvv9wZyg5QuQo1pD0ZonNwMeymnOdq1kpVqqLFlNVaxT8iAGA+/B1h//I7eR6VZE
O4svlxJZKaD8jvRHAvgHHGWVBK3QIx1aJ3o2ogvKhXmYp6LnqgGlUPKRmCMgObFHiqslr+3mV5yG
U+nibmXUVqcB9RDVWI9YXi9jeRvdt9YmCR75z06wYAZyoAX2v/j8Z+WxoYb6UgIGjfyfl0GwM8Y/
547mOek55gOYBIRkMh7NX1NpKAsfoEq0XvnX1gmaUH2H6/Bot8I5i9ZKQr6TmBHXxbZaSanS7gU+
UjRveIyLi+rsGlpGmgjOrUzy2WtfBSHY6b3ZARCbevCpk4n3W/mISVeEPbVgG3T4o38Lo2XluA1N
95XODny7vr2dQLmMOe6BlrWOJyQoQb5rwV+aeOyb17IkFbS5AHcjVK30yU5AQDzTrRb5CmDybrzC
+GiOqp8y5EJvbZKgxdZ6oDhgj/xPlQXO+yH9mCZ58gqL60t4xETJeRCEpGyrB/zdHojNHwXXM4WF
pJsIdaWcWlsOl0zln0OtP4uJxNG1cXvOfy5NV1Y+86Oi6bd/1mnT7i02lUuIjSqwFh4/rquVUrGD
wtX8EFEHlk+GWRCBmeyTy4AMCgB2NF+4CnBcMp4e6ptMjs/3tFeRYNnGgRC+Gw94eej+Gp/Qn2F2
eEIdBjj/FiqMBzl/1+okeJubfFz9QEAwPewIRAnUElruz44Slhg+LaO34dY4baF7m5Njrg9plUcC
9VmzCTtV2xSWpH264wwjUW9JAevrqGRGlaf7oIMjB2Plm12ZAgOxTZE7yqTheDveurEcTxofBh9r
h/RRS00PgfOqKvDs8W6ByIDozqgQ6e+vbcOcdVligX/Jyh5NYutd/yCs9CsnoanLvqSJasKQvK/h
r6fnSPHfFgruLMTS8vIYIXwWI9rXWJxYUAaTZMD26plk+N+PMzc7QVEBRoyCLZJLXHYp85CeMDhu
77PHd48Nq39UeJLE1poiV5Vh+u5TooYWVV7xYqvwHxAvetC1heCv1bC6jGltZ1Ypzge/qZHAReFa
ugTTXz1kIGi0tEWpvVXSrc6/8R4i3F/XPxtxWmlxaOhEPrWP6DUK4wF5ZpfHkEmmLo315+F5GCXP
ESJ6vy/hgb7uFPXYwfXeO1KTgYe4dBcLWpT32EpzUiZWAfKdUPK2y1O+iMr7dPj1/p97cvDSORZp
FZxkXzViMd6vHmywt4mL8psT/txDz7h2+1t+zEpEJCdNrGQkKwgBglRWbdhghuM+T/tq+EBU5Kbw
R49MuYQqIE3os6GWnsc7lcnREzT9j77B4Zgn/WyYD5JHAVZTtpxHMSrEpSEm+dx75m8PwOLgu+Ua
bVfk40mpBN0GRj3H+UcffLIYdxk4tOZ49jie3haE2GBdfnHUhmwVEepyFR/kMtvKShUTZ3SG7v9r
G97Y9b10gaV15yDaas3U5Wmsha8Jzj4UTnJnxHmGC8Z1Ddcmhu9fUMcD0p3gEz3OhlLuZQvUVqu9
6bRx5wQ/yu5zFzKBlro55sdgCrcI4Iyzh0Kzl0ubCvgTHj75T7WyI83388VxdSfVRJO59ur4XB8t
FerdKIXis9gC7nTwpGIP0AavmRoUgK5PNB9cyStzWAcH4SaDjgGQw6G637X2cBD+Sz7VHonQitjB
B6nMRT8mvFqgYoXNRYbRRHOLat+b7r3o7I3D9BxIq69vbwxlxUZ3j13giKVqXrxEdhf5SIPkGetw
54liOsHLM29rRX3ziGviqoelR6w4RYiCh435gxiYLr0MYRCs6BOfpjHzFKFfBNlVK8dVXAiIgpkn
Nbwpr7QGZ07Zi61D7nNvEPtnfizSROZ+7HDmVMcoqzPIm0TbuOOyVthLWD2r3+M/kCQg38yU03GP
vERBG0ibBX/Hvyewzb5rNumlWcL0YHMMBbjrcZptLLUv7OZjDbAzLlUpZ3e7wG3b13z6Bh64SgUs
NfETAS6vbIu/Uu33jT3qREtWv7GIW4//ltu5sG5LjccXG5lOxE43P2VB0Cbogiefbt9jnqkq7xSH
bt3l4gTK2X6SxqL5EaDBTSAtzCEkyWY+/FP6O1xXGG8oyHyW44J2gcqgnQNJ+42m2y6mfhoKg393
8dRrzt7DFGkrtRi4ZF5PTyV8cbJjWC8Tr1e1QzXGMzOQSiyIjqyIUwG6N0KOSrFRbEvsuxpBpe68
91q0tOxw3baFyPiDe7kNY3cj56j5k56mRml1kRjIvMcaRt7pfxg11rtDQDuEEZXot00/wAxRLYXG
TvhHtmgAktMDeLQYgrwF3t3D2JSHRh64akhcoIRtw/yuztm+QxG9CAiTIXEMvUn8tqfjjEtQ09Wx
5l59tTBwdjVpokUbm8GAOCp0Sfm6kjta6Q/3omAqQMyBE9oiUcW8tTpH7oLIbOs2wpsta72qITwa
NyBMWdFZ8cXe9JeMCimjkqHAxHswScBx50huIC+yqRyW4SCVdUg4R4AP8VjE8VrP+9AEL2OmQceo
Vg9YBqJRcXMyg2u+LV1cIri1JA0Y42mSbHbfXt1WUl7Y4sjZ1NMrErxaxXA5eFfNbpe0/Lw4NMIu
1AS9v5HOjzBjaPwIe+OSlsprCpOCOwPbBVuF8MSNXT/ssBil+2hC94YGUIZBzccoIPriGG7E0VmT
+xPG7F6ydsD0nUhQcL0ZQwKMVEr39c8yiD1itY+Sfu5W6gK1Q8/P7YQFiruWj+uBPJNtEQqVP+As
vxOGGG2t6PskcVxlkZmp7SWlYnml7r07vfmN3fEqBYP8HxXDUnFuQKfl1YfKTberqYBtoumAYbT/
vm+hoK8ZfMjx/L20tZrCcZmeukP6o5dT3WT9r5JQ9+CU054lWARKAQqPFGaZxzjM24tCZi3BfQoh
j5wm0uRaAVVSfRboUI56Z623urWsvwergf+jl8rN3oOGQ6M5DkPswzzY5TdzpGZsglspBZKyZYfi
A3+CoMYejXfBZjTxKKLpdpHEj2757fbTWX/zRFmzao6KL9U+akBKbyCACWXWSki4/vJudPUTWxWZ
/XHI0UwALx5DmGpadX4EWCzr9rZXToQgpyYJiIXwzb1TlYnv9Wp1lTBj2o6038Kpqh6pBoX8VVUb
Kqm6lfgPp58xnUp7JbCTfBNYXZFVgBgKXe/Hwg8rhqwRxm6GwTW5DCuMY+/J2T3cnO2j9hRmi1N7
NNeuzqJPaUlYTV3xsZqkcbIssFCWpTiwa7YPz8oTbORM0WJLr1k+KnGKYrOHfyyk8J6BZp8EHwiH
JRp75hqZ0ppBOT/BfcneKe4bZYrtM8PgmESPYBE1PyuJjbVUvMWKaIosg+OlzRYbtnzLFLvP/3uF
tyBdxwtUAxk28+O54rCC0+RRlTa7BBFbJcTsiRkfG091EnyyC5F/YwZzWOx3NIzDtWL2sfzAwuLN
/TML/dBLLvZtBeKAb4gBWHIHumjQHHOeAqUMV4Fh7BM7CqgyvRg3caLM6nof8miyHdtm7kKedLDG
gZ1Wr9SiBgHz1veONeWdMo881ibH3adPf5VHUScxZkuaMMkvmqZqSoW/onpp4or6g9A6+MiX+zwV
RiZGxO6jn3GKb33HfURt9+315JCMsug+F6PUUXc9wQBwmJqk+3q9rd1T8XTq6udnH6GMEcqkzgtO
axDgzANXvgF/SvtzW5DH+iLvtM0YIBTGb402QY+qI/RaFusOU+b/7Vqpfe8ZDA/LkepOhlXenoUd
tp9cGgBWFZtf8r9xeIwdUztyKUGI6Ke4CW719tpVmYuj1UJka8jAZmdIT4+1lYP6yx1saQAKhFrP
PCOeJ2tvLa26BBtcHIjIInms6ER6EjaTjl2jQEfn9t8/3bYJyiHDSPPmJgdOd+WR0hnRgnali9xb
pxxoIq/59VaIsYHi2aDNOiUeRV5ox31HrxPIUsXS23kinMd84UBkfDh8NJXcL12/qXmUJxXGtGQ/
7lcCIj2HqHJArtJTRWw+hmWxud/ltl+hiMlV2xb6CX3jY8iDbZJwPX4KyUN/ebwsn5XsRTWoLb25
9iiLt5ody3/31j4MQHH6sT8c4IohJOGPlPv4ISdwLAe5oXP0HIZB/N3VxBk9VK4eyxYClrY0TxnD
uicwc0izylNhxXaSrwL2NXNjMVC7jBTH3Vz/EDv994e5zmcOJAovX7COC+mN45/CoagjyLcgBDxa
HIBQRXidYfladY6ZQugu/J9DNxoWN6tgXVP6aICPN7cjmfZXtSoL49RdB6lshXaogyrJo1T/gWqR
4sp9SrCKoBSn/A7dgGtPV+fCbYBn5hzXSFtVCjljQ1UDSZCIPLAKyINrl+NwqsOycaUzeQ/lWPkI
jv9gbWyl4bSmtKZ2FXCHF4tneuqky45aIcYicDHebZJP+BUq/a3k3kdoYju4rDplbQMhp3l/2HtO
ryqg6RZW5WciG6rWBrfF2fd0DKRECYQbl75cuxR9ewR65DChHYbb+evUXSOAi00MgX8VD+aJgzfn
GlZ+sovnTADjCVr5U8vrMhM4BKWbsPjxjdb8RkAovVEuIZtznUVUk75PDLiDaS1xznkJhy+MSt1U
yF8IT45wGK0mFRZHbh4KnNQ3Fj8HSQXxmZJGP2SInIJnDB+Swax4n0B56308jkom35JRyNVw7jFw
WhkSIr+vy7knrTKiNAMfUQgOTwSM+WZYyOwfcbMBuojJleCYE+HRoaYMuU8porjKhCKsfAwO9D9l
EvDNSuKFRKbVwFr4+AfWNUDxtt43tsMrZCQx3AccHAOlGh7/ppOaEXILGjmliOm/RM0IwWscVIxz
DpvovSFmmOyCtM8jDGI36y1OBhEt/j6L6ey7PHC4M11gBHENBvmLETH1T0nR2jYsfoNKC5b8Vdjw
6askDu1OL7GTGbGMiEvIABLFXFiTxpW1R19K6xTcj2S+d/nPNkSRBujXb1t6FMeu3EyxL0SA0ytd
zPEjubqaGSyX3OHAoOM9KhFDfE83pCAc2wD/ANudlt0EPefp/KOhXiOxRr27yImEVUMobLQIziL7
CcQ1hglPLUJSoB1moJiuQYJMx2Nou05qJptR4DByCBBJR61SsuYOKrlj65tmQm6htjwPh8P9ZG0n
ZcrWEBl0LJJZv4s7kPhvrxasQ+smxNpQsrHAAkheTM16UlkMlm4t3t7zflqZGM2+sNjtrUzghGt0
LHmFg+ISWKy5YnhE69Kzlk+xrGVxenrzF6p/OPlYmfmhVW8wGNn1obpLvkBXK/JUIMSV4IcxY/11
87MRdoADgnzgUiFXSTH2uOcpFFWL4h+GcYk/PU/pqHzPfDvwcmZBUGZ/adfRJ1Mb1a1MwkppMQ9z
pWmgoTCGZzn0e8ndQ/ujs77fu7z7cMeZk/BgHsIhCVoOoBpHknYjQoN1CLEE731PLSaQFVn7BXYH
COq6w29tQ8yv5mveytZCuQEL2TDtQtQ928oJeIFWsGo4wZWsM3mUYutMUbRRv1PG0VDzQyHDRsnM
T51U7/PiNZr3SJb5zd9DFYKORnQ5VWKXpJxHWUsK34EiGgn323ojOA8OewCrQeU0ygd3j6Msv8eF
673mMrmZpxLF3v9heHN7eAcl4yFv14RrjpwIQBJ1/YK409snUXyAUqRxntnqa2KeVDimfcnpV1U0
eMW/eTW9AG+jY7rPP5cnZIx8JzpmEo0QZvr/+L+2cnr9KbXaGRQ9TGLfq2woCkDckB1ezfy7UknW
87V+KFNfmltCUrO9CWafPnwxeFUy8/4tt9cY/4Zv89H9afy6Rfki+Q7hqOpJ7Pvs8PwFdTvsf0sZ
/8dEf13EyTsG2S21G6KGbbEcmHytrv1pKu7akDQ6HCDtlFAEbrTDc+aYW8mjc3rzi9xnGsESZjwS
BimxSrvtAnO/ESw9Bdcr26K4NxFL8hLjdbUFK2LuQH48n03WdEDCy36BqqgXETkSRWQ7iJJ4aSAE
Vg3Un6IP1ZP2H6foZeHKtD1JQLA01EDqvslaenFoNPmy31x8XThzNtr2sFN7mASBIf0g4vkBlYW8
U0wGRHkHnbd1Tjk6+RBMwkiyLPd/O/T+D3NBUIgBceCmi23u3YS0VTRPDKFIw9PkxIHVr5jvQUsq
gpkJxOsGQgm4esxGa6hyg89n8D31iWZCsPxwqjzWFEK9UyjtItcpwv1kcJWCrcTcto0i0etiGW1B
se+DVuJK2W9GUpWwo5Y93jOQATE9MZhdLVjS8IpotIMUPY4/UMpwE92S9CrhkOydfgxXFakISnvR
mLTLg6IUfuIrHwS4MpY0r3sqaEbyNe5eY+zi+Zv4iYUHdgSZCLiDVrxCCeqCEX8F8shB04iaeYEN
3LC0eMRa9b2uiDNBte5SbvYfsmhb/emxWsZ83U3YRf3jLOaaca/lXYN/IXUBWqVIWh6AYZetumrP
qlWMake3f2+ZQdARw+vv6+xm3nfP2t3PEPRevNDEeYDLoy+BM4wsm+S0D6wVqcp/AeBANr+VI5dG
tXvZ9ChCYtnp0iW5pkb37+QPnkqqJSvw3r5E+ei7XHfRnYWUC4jtimF51TvMQZeQP8ML2H4X83Ig
1B9psbRLpkpegcK4xGK95zhNbfW7ex7dm1XhbM09Wvbg3LVx0l7KXTC6A0nv8m+ynGWOat/Y02Dy
qRrNZWB/UpfIO95Y0JCkdYeFg6BCosFrSl7PT0Tgx/Uqws68QzM0zQEONJfbUREsy4rdALAwqOPH
RzqQWTMLkWE0FxoE//1gilH0Voj5JSkXD5afvj9/hvGRGcsuK7bvdjP7AhjB3sLbPeTDmZbihtw7
cMX7dtF/zfVbJXwbxOOdhdATIIS2RYIgDfVTDCUPtbTnqsFIzkizUY1S0OSa+6khEk2YnQzfgQ4p
cgOZHrPx0+jHXD6WdCeWz2cVE/RDiT2/8GK2OcVN5aQv6mHd2zHq1gClERC79C8b8d14N/uB5ZtB
H8m9ETQrPd5gZdWgpjfsuN+n9pCLl2gKQ/wjRU8sbEbEJ1X6UiA5HjLiwqNleab3RJZ1M4wYEj+S
wzvuUu4DXKIFmn+AB5hZGQExv2MsSVGgWBA9p9XzQWa15JHzaiAM/GGY8kiOxr9zaEDekszrxb0W
WStlsXbjw+aRFiqar6M1C8C8I22qE3WpP/hdOyjxZNh/Ps/Iz77nZBQ7HtrL4gq+/7cIXI15qcPZ
I2D1EE0NYWgUt8+bWf3xebIl5L9VxC54326Y26PglfSzw4Eww+z+ViYYFj805o/AvzH6mURV3hJo
5Ir/J7PJ7aQJ2ZOmIf+uYJzwMwtq8e5sOtZaqAucK+Sf41ct2LryX/4uKIaEeZalBgG+1gcrVq36
iTF+7ptknQ3LDFUfbPTM1s3kNFqTfDZbvUtNjG2iky1tggu946z3t1IdA8xfk6ePF0aJQxtFJMSb
xrmbpeWfnZ4K5H4ZYoZncRE4js3ft77Y4fLenorgn2KrcvOCDYZJnTxKB4OdxGF9ir+1DKKPWHMp
SOdxYOVhj4+bDuoOmGl5/racBZYDWO/cn37qTBiI8yvlxFxuWsSPqooH6AWw07+RAmyFx+f+m6zQ
NcTXtnl1UsHLDb0UyLaW0/qhJ0vMntq+aFq0e261oBqdUCfeN8e4eQ2EVwLEcV29kUbIVyzD/99A
qNbzlpFBBFilzwEgeMVh05mlHQc5mIWsdZfp6a3f+85pwx9rUDsoI+thNhw2Nr9T77QbpvjoM0AH
7gPZvoD0+3srxgDtgPsRgICDr9C4JL2Pt+WIUSZC2Ab91lz/bqyAHAu5A4OxCZm5Idnc54Ne58K9
7nx6GhusP1O7m2znZoDDxANj2sAmjnbwnAwiafeqx6uvn5EKI/VFd6AfFuxYqkMiNmilYPw/kXwE
n/Qw3+1rhfummL2f1iprzyk4YGopnhN8zRRMiqUUPGkdeCv8LczCqzJNDNRryHuuMIjILuOVzEws
yWWPbHei9q/roa9b5CllE8n3TeFojrlfvaLq/X62gM1tPFpkYWSkoEq9IJyUJJTWVesvI7xvK+yC
WYFeKUnfaunJsC3D0yRgww5UbkHwpMkG+/Poe2huncJAuktB1F1QHszYWXLs97ckDBgoilres8cS
uyHt+KzO0mkXnNcwt6dhWub2jFwcurDW3xPFhjS+EZx/XWkGg3oGWlLjFON/GpaBVqxbRne3mxj6
fB2g7tHs+Ba92J4DG4xWHzY7WUx824sm/jBRBQZbBwN7Gy4/IrlPkzAumYxnJoA6k4qGkUu7kex5
IUjsR3lwuP2o7aTfwJB/SFx8VfEJnxbZxFV//eHgq6LLiFcAG/0eWR5EvwxWx1NXXanxaweGVfes
TdytwarO2kh2j+0fEM0Q3plYOnkF7lfe74qo6p9nZVvVjQGQTa3Oek9twe2ZCS+V0zC9D6rWhZ9S
fGxABKWacIxM2SH2jgGRuGbi0s8VrlpVXjvV2q5X3JCsQ2aAVRwmrCvGdx8jmPpClUSeoUA7vDSu
JvhWMwZKmnGqcNsXJ9Zs1WlAmOTVjyCMFfotI9K2vKjxtX9J/sMrIW4qYGoQgjfZPdYd2S9l844j
anzSKNn9e8nZVTN8+qahzD4XAVGvPqPxHTYnPn7ITR1qoHu7BHKRCTCc5TLQ8ZK7hB+KnBK7px6L
Oxo9suTxuZzYCJ7ZV+/akldujw5NDwPzV5RVmP3GX87tWPPk59ERh0mU3ehyy8xEGGmyKm3JJhx9
2eoVTeDf/M7GcCwmO2U2AHGHLcHASE6upuLs0JO5xJDhn9dmW/vk1QuOc/Q2xjhQH7uIPmHQJ5Qx
cZE1tT7ydKuGb8NVl8bj2B2CG4H1Km4RLNBOIz4wM6pKupw2ZQqrBqv3CP0vpbKYGfd8KOTHMn81
ozc/Dmsn1YfK1Vi0MFEOL9O0K2Cwv7DpKSG0Fx8nVC/Mwct+Jt0U17mOfbG+Ri82v1oH3ZAazmLn
iSGxOnEmnpAqI1fJ8uEL+oAyk+MieF8aQ2XGl5BZseI3q+WscMXwuH7wnzaVoKfoxPTH7s0JZBbJ
lovAmOQuDrZKQUpg6OrwfCvJ0jHwmzZHjTSvJHfcWwrG86SFjP2AZK471GCvU0Nc6/K6LzArdWPf
7LVjMIa+PlGd0VYudXPa7dHfpWchF8k5ewazaf3t0BZ+hDnTbQTwBnVBrn7WIAbyjJYOYRj2zHHo
aqbMmC/vlLzsNqmkVQ4hezN1GEG9cp0yBGCYcG1G4h0KiuNINZlxskIKwlvFN9sbD/kgt85SKRlp
D5dH4cIcGGWhQw6q0cFDYJFsGdY0hxoqr9uNs9VsRqXhmQQTNZfCgmk4JAB5Hc/LJxzLrJUodkfu
vflaY64vaj9vKjZGqe7piebT+YG5KUPE/qmu1CVAzH97MDe76zUbFMJS+gLTVXljEoWLGiEkCim9
jzkKy5bdO4B70vANvZm88Kl+I/ZQv702KyEdGv1qzCmZTtxeAalNlnho+w3ETN1bvei6kIs2pA4z
WaK8AhMq9stkAVHaVqKz88L9AmxcZdqOmK589rtuTSDCe735wURPxD0Z0Ql9HW2Rvp7BI5diWoww
AcP7YzK0keqJLIICeoDZNm9Bbi137tIHErwXIebMekJQnNSFUXsSrC2XnF4Na9i+NTAyURNqJZmr
xTrHITLIL9Z6OcP65nQm1vmeST68IY3AXV0R+y2o8IHx7KEE2X/Qbd3tpIsCiCyUgT0+I3IOkAI1
Z01UkOX8VNb1XBi03jVFoCIcjYVUAcQJdeAuOaoEfI81A4img3W/6drzVdKdJXrPXXzN4SSZuKUb
LSCFNRfPBwqC3+LUks9W5SkeFZW5tFFa39pLJrKCMGDgji1pjkNW6ppslFA3mytdbatc0JOCPkoH
Y1jag+saApwHKr4Hz6H3FZCDgikv4kwi5LywuYUAuQX7VHRHgRk4alBmeQGRFbYeAz1rWzgxihdE
B5EEt68rUV8I4bzApRJ14J0QG0f1ScWwIjh3v+msk6JRVloDT33aPL3nqHHgBXXOQ+B1F+4HMA9r
RA3TJV8fjaw2zlrTvr844d5QHgSxHaPG8ZTLXJvStPoyLUA0hH6mVyD2swnGf2TD4/BI7nNT/iWd
Ey0aqhu92o6yZRYTz/eiqnKtqQLKBc/BlDtSJyOUUuRq7afp243lGK0H1L5f6imaO73EvLeSkdZA
dMFPKkBhCBnPRcWZ+rJzWzCB/N/1a+riCEfGzesL+F6LoCx/rwOxX65t5OwoT7u+3RULGh6Ul+ug
wrp7HpD19Uz0139fF2z9706iQwzxKapCy+yzY2YJZvhyCAlVw9wxM/WM58NE8pzF4OCRLHQdISZ4
eytrMlDsuAaTIwAfy0hk6TuS3gN+0O2rpKuTGFREgQyxgK4NasqZIoz6uxQgMk2ckthmSgktdSLO
wmp2O7KTNK9rEYTnPAYBy1sCNZpWqvtSianX2E+9YqKUiBS5ugSMPsVB1vIV4oZ/Io2Ubuof+5x/
WOJmXYt3u/1E2V6AOQx36tPQeDipzL0TJVQzBMCat4NVeUqdWA2zi5DgaW/rPM2Rbhee4xAV1/hp
YAopISjfacjLFmOHx4q6qx0AT5AcyW2uAP65GkIQ2FezgUYjGYKvJODVkI3YLiuDYmYcPkX0WVnC
fcSJCpWFAdsY3PLpUGWsfk1/nM8GK96CFDtwmD/yqF3Lz9RYgUxMiZft59ts0zfrpZwX+J4X5WFo
Op0+gwCbXGX0SwotVvsdPJpNsVg0RQwvgpygntGSLV51MqLRY059tnYVlKDzEEkJ2dUh5hgNy59/
Mws5ekjiqvYmoM/Zu38StFGL776QqQaZ+EkYDyNOe80FuHWowp7GbB6Emw6tOg6wIhVOLewK4N7x
BjDViz2fe/ZKZ6J77Dy9FidCWOO7xB9EebCE0fmjgO//OhKzukkl8NaouRpLMBzQ7G0bstbQvIm3
FBEC3JlUMIAp+WywfSI6zC/LN3ww0QrQ8UYsHZDogxZg/jzm8ArB1M5TcDBEsHIEwi4h6YbO+X2A
FwDNIPgb2shn+jVQd60wNG1gBrAa1xo6IbYTnpSFkJDnHI1R++Sb6EMkHRPYogBlW7zZsanp17Qu
n4TZnVzqAyazSEaE2dlgMtF/YnRU9TnaT8efOy/cqnijOgUU+xqoVwPfiK9QH5dFlARgfGQ7JVSl
Ga8ycq4drqcAM3LSnl+0YFwgqNQluz0v6sWVKI6ZbYoQUEn0pKzGM0SyvrVf0edhJ1RD26g5Rg9L
TmmHYmUc4Y/yfjXGn0ilSb5IuWV+2i51bNyL9vVdoVkSrXh8pcsyaRBZpQBkbl/dTZTMldsRTC7Y
JZHHT4wDoAIi8PCAiIKWXRkRO8kxZEAXKc6G2/lltES7kLl3hyRUibP3e6Ard16QrupH9L3Y9R+z
mTyq9Xs00QVIqfUSsVJPe1lHCHbADH08zdo3/tLruDWGMy+MxR1c9ghFFVMy4PtrKJ0De0GsEV//
Ni+dhTQV8+hEuw9iCxB6QLFPwAFevRhvO4kiglkPYGDw/2lVH2DAWhIbBjLf39lOG97gpL+Be0KE
kvy6Uc/DZ0mL2LfIdhZGxS6SvNdoWHF9XbpdivlDdxmW+N8w401KJVcN8vrlfLxfKA6aYAwymJWb
iXCPok7nJHv7X9TPO8KQih9877srcQ+ErMegJz7hF9LIBKKt1MONM/ZVfLU++20MyPVTJYIXtSHE
NgcEkGJ1K8iAZUQwxI2dZL3gR9Mm7m20+G45iHi7LEbWA/5Jro9tbkn9+1cz1AifhIEgJEcQuD+w
bZLdsuuBBJyvtUn087OkX+fOmIPZxg53P/u9hmhsUbJS+izGL1Kig/CEC0/9150Qas0saw5l9Ew/
U+fWoSN/+s3fDvTJtj9j6TJOSlP3YAEV7+c1m4buaeO3yMmhtsEGS9iybHs54ygsKD1H6XN1I/ln
OeY8sqOg4dUO6o7heY9Np6hJRMpLDAqXnarELJh5KqSvO4kNiKpV03+cWe5GksiQz16gxeb950x/
9IgRpgMtNYKK4GkeP1hb9Belvd4ZuumREugLZzltpAA5Pg5LpkgmO/WNhdh2nAgoM2OA6bn3wt5g
2JCIdCVgRLdAu9JW+3m1x+YCv3Q3GPnvAYv3s45ur5PMv90CcXJAAadYDvMVhfaE9IcU+0miQ+hs
Ja6vRDsnprF9XJ6Rjesqh6hR/6EfkW8abC22xJU2D/x8U41OgFQ+jle9hH+2Uo7GI9SsWT4gES06
w+UJEmU5ar//8sMSZo+mp+3tuVwpeE8eapmhhgMKNdBaHa0ufFGxgTwptxw3Pl4Y8xqDNTmgdfab
11XSg5PLiu2LH+ysj27mJimwRBoAe/f18L1wNIxim05b8teJzsz5GedZvFukL2Dzck3q+ELnOqTZ
FMuLQYPZDJW0Y4kXb5lzEDjCuPchKbFRr8RDExFnmWRPN9+t25MRExh5APRGBPgHclNSKfWacKnR
UmlKGEGYMNsdRCfazH64CKVJ3IxeEBc1OYbsOE0dqOPeUHrZAQXabr4vgMa2noWSX4eLSckmsEs4
CBjZHZcL9GU+rjBfoLu7HBgBRN3Hmomb9MD43o84h5otJjiwg2Gt2CEmwVVbEMoTIJdMOIopoc+a
n6FM3JirnpvLCWJNCALtUsHyQuZxa3Urj/HOY3GyE62Lbq8UQ7e0l/SU1Hvxu9O86rMZs8Ejino9
7Jqj8lfn1jWZsFYtYhfJAKpM82H9zwJx2lAEFBszWcZ8IK1PZgbQqn216PsD9E+xXGeKgMuZbaE6
JqeV9jcvePYVIR1jk2/KIrY/fxMKN2yKPlO21qW5HykYtzxvRHbdd6k/khy8cQBoaWd4X06sfgvy
57AfJhahaqSUvEVmCIjVpgQ9s7M/MkdW96ZWJla3NCpMU89h5k3HSUOE60NBWIP+NtAMUtirBZLb
EYWFDFXULOo7sEDzXvBpEKIVsyS1PT1AYj8anUWulZBvPM/p7uVpcKTlPQ7DPJ2FgafifHFAn2Bq
6sRiiFd+vHWPuSo60NWzGmtON1NlGSJ7bRHOuaW4YGoflIWFkql1dE2piEjLfaa47VVvCay73H/+
6bXCibbgpRDjMD9gAeHlkkEyk0L3lWsRbv4p/smK/TF2eh5iX+FhtrWOMEVv52b0qg0mSZFPSRwI
BWvsDMxSZiwTr0Zpo+02LpUbd5Kat7t/2nIJvomrWFQO7mN7NyIm2Zd3QynrURK+2WDmz0oDQ81J
E8YNmUFQMEXltMhZSrBoPUpd0HCZBlTXhgptVaZfip/1cGCgXRlFdqtPNMvtCgbxCqTg5f6FhtY8
+EvIVFqtiJRBxsDHnENol0X2ub9SYzk40YqkGf8B1x7r2WzfGJ56LMF96qvjnIIx4e8OqF1CwAjH
57bS1iNeX3B6bdGz98CprzpMm8Xf8p3mOSjH9WnwD3VU+mSsfpqptZpyr7HPYVokgqZRr+aeyCam
4d6q6pKW5LY+yQuaCgk0BurD+cYjPJWNlzipjKJfXZnMIrEniLBOeRKpQrM5S6sN8x6s8p64wR8C
xl7kzI1MN/AObtzO+F7G3kwtpkMJdmHmAOrzwwV5G7Xq8dys3V4inciIeN+1nBhU7q2C4E2htOv1
3dVTKQdryeQISyNL/fqO8rpS97OwVFL9cWrR/5jM2Botab1Kmc+gHyXhvqUbuU3O/gXgOqXacjfd
5uj0IiriJ4u3aeasx9PC+l5f8xcI1WkMtioz2EvW8jbSWbHIVj/Q6A82bRypdO6qDNRdgZ28+WyS
WbO7R/ipQBem21VGfPxB9Z0+QZgF5Xlic26FcvIrAkhhlx7HJpy1s3prEqRX6jtLX/YWLqQFEKmf
vDcupb8pfKJ4kiVVL3Zzp+katnXjTdUuk03nuAA0kVUbiwQB3/7ASeWrYB2G+GLlUigcA9e0JqXU
g/pzFiXsz68jBKxYsv6bljjWvlw3nFv/asr+oqoP5GljnWT1EwQE9Tg9HvdRMQ8G+GAxTwlfUdub
xDBPJ/Jco+uXfW8L/yOfD9xXJV5S7C89JhOuMhqCSgCPctzlRVuRLJlc18SONh4SsOB37YNPAWBa
dzqAD8fq01Jp8PU3mrn6kBN50xxKxGgWxbeApReV8KMZeD7ljHKIRP5ZY6o6zsXCuHx0uU98/42j
VmAAEhoqxBL95AqcWWHVZ3H6CxkUIkDau5Po+Mtblf91QuWTRByfzsYquCuzYCySXHhRsok79Vyx
wxZ8TaPKE2VdCU9Fky3ez6fWCEzGaucV3Ns/GvyS0QOAQY9QFmL1UPFPYG6CzBmBNB0CbNA8q8zs
ozh4KsjkQHWoeyKB/WZB5dNGuAdazQ6RKJ25NUwODlw/l8QM8edA7lkp/0hbpwkUQvtW0QJfcD3T
KAjPqE74L1pzi2fxg2bihmYnMqTbaZ6YFGL3q3KvnnXwkTWWSGLqXyQemIjjDABalbfO6TTpfI8E
3eF/bg+QeQ9qTQA3wqa5TaktVnnBDhsVbEFvcyTqixviPU6c/4oKHSZTCTrVp25ygT5fm0ROaYXU
KAHBl0kqnnv8piKnvHiHfMSIzENcrzB02mzDtJbx1Ma+Y5P4s6dEsyuZevGRwWB5Ugn23Ofwgr3B
UtWpm3tcswhoIL2W58H0b/hM2oiXY3uNbEu+HA1kTNYxCX6CATbmA1kWjpg77Up+O3wW1U7v8mR2
Y/G9yw5qkVVNRTaqFqnPWxM14NlFhMR7AReOhfIV2TpnHUCvCt0EoqBGOWLWYge1M4nNNE/5nlxU
Ugv2zebI1JRc6MvcnQWyimDhz61cnizNtlRAV91u6cg5g1JfaplL/IXNGcg8tLU5FIxU4DOvvnl9
oKDU4YphSPjqMf9cx/9K0VCzpFfXFdmezvLlgkCnPboDGIcXNaL1FLuUaNlRXL+Us7JTzq2jpoW9
EY0HE8O9Xxl4Zrcq5yRiSUpuBAsk8lVvrlg4d0KhkJbdU2Bmp/wmWMuKhM3Nr8CFf3hE86NldNlG
wt+Oz3cN7+TOM40KAxB38JYU9UelIlu4lCU+SyxZePOUNnKiNM3xpvT1WbhBru74/H3q0rBg8laY
R5l5PXYT+QoAKBfQbdBTHdShX3f9iSGfabNakfMZBixE3hnmMi/QxtTS1wz4Le69k4NQpoJwuLDx
TqMdS/QSmDwuveNDB/BwqVT4+0ehvxZ3ZqptF0ipBDNj0kLnf1hi4i5ki8JVzP/Z3CCn7DXG+lXa
sOuZIohfu9IDHPFTZzJIV6SIS6bqvgeLnNxWq7FgiQvr3k+JMBThvA0JRa34/5GltZEfooY+i15t
1RYvGhdhepeB3KpeU5wNeWbUq6v8iKHTkIerTZR4J7PC6LIA5W/q7mw0IIm8IfmnIP/20L3NgSIC
hxPhhcmCoom2x81GhmGqygbPNv+eVf2DKq5S8hjdEKCl7SFPP3PH/2ZEZAXLdV9HOcinXCtQHB9q
IHzA/VMxWg3dmyD5oz49OwC7Idk8rCu9TWa3qaLhr5/OGw3pOR2P4u/ynl91QqYUtxAuwDcY97w4
ucU6RksQxzemF+EqmcYdf+GgA/binhs8r5qUXSsKpqfCY+QJnFaD35raUp9WLFrx+wVZHGrNN1PY
GX16J8I5Mdm431966kta6MctQbjH7xlWeCxqZzGiYq52O9Z0cMUaJAVnW5oWFGTyv+lrg7pUAcc6
ggyTZkFAuKDiefnJN/08NepMkEUkF2zYhWNIuP4H9WcMBTTqZDewo0M15Y1wzOLY+Gi4w+6malCI
2u+CrVZ5NCnJULgtDME26DDQ8QrrKilD0PoGYMfBVLU31o1nSPdw9FAoUEW7gj+pL7Q7Wq3mSqv6
W1KiHBSJQSc8pTK/b5j8lp2wcKeVlLMMsKpQE/OY1a2dqgBb/2VUaDo1pXZ7ugWQS4+GaK2GDIns
OUptJ8i4naHjNhTp0PtaF2VyHdqAfsRh4V8qBTQuqXhGgGbqtY5Ff0F78AVdWH0W2uPJu9lfQQMa
ScenHbOwnwcCpVVtnDlylr/OzEgoMDvSH03eNkqoyacr9cNQutpRHbuT4k2TCb6qdN280j25qLQu
/ExvGBFA+Y8cmzo9ZffMbTNdwTVu/QmoTgVAS4xsWGkCxOLGLbn1z9hurHW09zFx+KsAMqIkYlrN
Q8ix0cpfTQ7kIuMcW2jx5AFnL3VEtLUaLBfP+Y+ApTlE1+ThddiaYQWk/906ugD8Utdr3z5kdt0b
LBWVYEZe4mpNN1DHBlQoNNIPX3+05AaDg5FLrTMvb7iK8byx8EKLRZvuUo7Bd/pzGC8/YL/mfP/W
aqVzojHuhfSEDx9M+KiU6qi3d0r+DsROSNaewy5jd00lOMoKpBgvjXdXibgHDhvUHudobcuJKJ5g
xx/RpnApXlTK3P2NF4RJaIu/x1CeeC/A+UT/82I+9nQsWXnF7V4c94mp+MLnsshb2wFqamJY15DT
edAgs4eG1n8eQOKLJZbI8Zlr5FlMPknmlOIcDCGRbPcQgVktOk6YzT3sbZ/g4CPMoEDDFAAHRm3x
1YwJ5ng7cAXmPpWFqRKSm1nv8OYsZbNCXzE5RxcbHZD7VL/lYdr4CgmXYOwaBOh9GrLgnCgROfvX
+UzELN/Xh9dlCiEoNOP9aA3qSg8hJ9b0Tg2A1ZtwNt6OVU8a9YIUPbQHtf5XRPw4hdKBom90LINY
6pIMg6+dcgW0twr+61omM95UqOK6c+Gc/X4ETNllLIxBvoP84pOuhHLjaL6vYPd2g/f3K4axxTVd
YgruqqpE2enrZ5+rC9cluSKi0ZLW3ulmyG8gKj6xmbPUhqwajVcXeOrxiyxlKzjg6fRpOoWcFTcZ
m9u+TZIupSyrf9x8J+1pZJEYrcwQ15igMVzwpepb7VD4viBlAJKnWAGLPw+pAe3FHXWLwlG+s8RB
PQ/BKZ6vC1XHuDKVEzcUNd/zzaz8KyORjyP8v4SzeY7Wz8ayjO9zhHUbPySm8RA+tULH/T8dO4LE
l2hfh+BP79JOCElcVr8thG8opXXo40ebQz3luS0x3m6gX0pKxCJot7Z5HPFDspjoTTQO1YJUpQpZ
fo5BMgTB7WFxH++rMAAK/Wh1hJcnp4w1Yj+igOhPEvA4QRVny2foc0mHOH7WcXsUH2UZ/51c12QI
Roh8KsLE7tNdYS0b0/yKxuvwZDpFwzu3S5Ztp+ckvU5ET06nsqSdTO//bVYjDp67fuVVCPD5RCw+
nTQ07AQWwKeCacZ1SunkOIC/t2see2gykWVy55XsN/1WmMY9i+y6QVacTxDvmF6D5ul8eG2v42mk
UymUAeXGevIPcIdqRE3CgTfH3JqZ1TrgJ3FXnNvGvYFNJMowAv0/c8xb2sZlocsETdqzwiLrqiqK
SXo2dHC3gHzSKVzSZSHzXe8VXaeG8mgAaq7QneHY1RAzMz0GSNu16uyQoSMoMFL7/wm6PAfyrb/2
XhX3BMUJcwziEzTHTvtOjwuSKGqIjtsOf0EZQ98FUQ71ZqzUVnK2Pt7V3yvNxKMAf5Bioq5/2QXv
cLRWl1tAi+Wy8Vuwy20pmUbnUn7jLYxvIv6ZpI8d08INq+4ApDuryqxecdR0K+p7cZKiOSRr6uXZ
dfdU1G4Zd6LDmEKK8g65j+bJtZt+Nu9Z+sWhsUALVxDgL6QRSJWvaUNldRzG7dAXSAO3jBuVGLjH
mwXhV20WR42X8alID8GTEXcSIunlq+SVxb5LrzznYzg2LHQx73quDhAYLuzqBWQC5zNRZ5BSz5Lq
6XpiU+9jjPHms7gMtR3Uf891f9PO8qsuFYmiooil5Zyn6XMWgIdxLaulPLdPCmbfxyB6ZbAxSfag
ouvds3XLCqEpwxDkzrZBf8OQO4rf7n5hc7dwxkKE5WV4Z/EnTUFn2TUoqSi2s5zARsX0QkoYV5xQ
PrOIuET8+Q3Vrq2CRwgkuiQjq0xJtAmoJoiQdF14Wis9iCcoME7j2a4srg0CmOPEucjC8yPzoWUo
W4d172DAG+pNj7qbBFQK76iYsKaDUXdvhvD+1x5GF9jw+g+iTWTerHGVmZDh7YIPG5pEIJdqIA5P
ijjz5p+ALpCQXA4JUeIy1fIbs0XBInRtD1bTANqEISqoSBDplNAKhzb/J1/ws9r7IX5URhSlxR2P
MTxYmTaej3gNpp9PsJz4zaAP/9rW3TEKaKhU/nyn5SkkDBREV/11llVQG2QPdeFKthSxjWPkUv0x
DvCxJUO6LSa0B/6dNqou2oW9a2gTstnl5/JHho6r4+5+OJrk8uVKcoJ2LQYMxVxWlwUZaJVyhfoW
za6EqPbZSmlOTNFlRxQWdSyb5wgknLEBt9f84ka14rgrNhq1466S5NdrsgjOMWSGOuqSbxscjPSc
U9C1u6pzSNYaU7OXCV8UtSKmfE+BXNvVu3sFmaLLo0FXEo5AnTonSP64tkw4/m/uEk4oNvK3itKW
3MeNnvSvrUujzd6JF6+pwIz2iPWFAStCEDwOx9XdMnfEwwRjbAnJjaCQA6fQvyBx6Y6Fe8yxD4DP
bffyOaEBk2HVnZ3J67SvN0XKpSlq7u++0RmajncoQ8wYYtkS6bGRsy0/i1pxtWK59kkMQtO2VZTM
nl2SnA4xgnZvgLJhZpOuY7j5W/uEoYsJW5OE84GF6YBLm6gGthWJJ7VUyBJ6M2sd/j+6aM7ZmeXW
YV/SsfilQ3Npvfp7OWfVjb1Jn5CQXLhPkxp1SqMLiLFP9Lm8AZcpBlhLDmLXjXDbmknnm+M8fmtq
k3PWLDnRJXBxHSOmksCzpxzXBWNhlyDv1cPWdjKUodiiotJMs/Wu4ySirWZNG9CAcdOK43XXIyn1
tWSARh8C0ggTbI6yBDm8wEgeZvbQTZ2OwiXg6gxO8MmxYn/f58uhHN2+qlDOBSCc2lugIceNc5TV
iOkFE3bcnpK23LsMcA2/PB2S95xtKsS8OxYX3gMSu1uXYUegICkDkH9eqHXIsdWgWdl2Z001CDIX
KFxWynxCNZSsUXiWF0MrN5sud6gyiSBMsbJSlUH5ZvYz2xZ97GdQR4ftonCmEkEsrbjZ0/Xh1dun
t5HIb1RT+AjcHxa0VAUI8dA0KOyCAzOR9CRMl2DOQwRiyx/Xyo46sio9yFDPCQm5wzf8mgN/m7qR
zEXUb4+NC8ghNfrcrxQVAYXXJv6Prm5RGWrGtAB8fZAkqv7qXS2Ls7ZUJB5iKmFv4STbHdLN044y
gkgrUIllQAIvh/TnBpTqcIeqBcKId0mbBlZaPXH0/wYrlP/c4h4e/54PCTYZvrGormQhFOWKRN1m
PkIn45nXyplpQQGxHoA8JXxG/aANeMaJXO9a2E1IWzBLJkJz0T/3cuzqyLY56rboz6kl1nPQ5FPR
ifNzNMMNI/PSz4YHtT3niRNVWGACX9UUElEnc7Wcs6wq5ctyYTxdSNo1ZY4cCXRLKKYYbFfRwD/r
EE/xDL1FNT8RnUhjPShjQ/Hbpe4HqBXEkQNAcUJjCGVdFk5PMA9irnZnSg+sELSWQTDp5Wzmx0vA
jXvdIolRKIak9UNb3VP00cFBmlBgEwdjYQHlA38rZGSkuoMakHGjRdK1KZhpcL9OK/ZWrvf1AJpZ
+QEDy8/KP2qEQE+pMglimAX/0cjNyYxxdwd2+rH/c1P5uboiyoAjv/YarTJ82dHdwtIoK0F9s+At
VMPdMtkQiYiSk5dsyYI3HilEkHB+KUo46nXQgF2uEojxX1eGbyhd1qGFxbb2CPD8SR1kDYTpuLqJ
E+iX4LiFkjLN5dQODuBO3wBaDkfxzaGK07XN7JVkRNMiwb9G7XUX3+sRVVKai6d+TBL2rdyGfSVT
r+F4bOs3ezHBy8E9WVGghdmV+ZD02LsBHeXRTgeuwZxQsvizsV11WDPN0IJ0SETt6BN+WHv+tICj
8N7/D/3DGgo8a1D7UP8zlSgHV6WYDJs9uNpZtXELMFrvz3SYnvx+HPyIAb+EyWF4fHgFAKEcMJ5j
IMsR+6OF/ZG50YAAf7M9J+qYXHgDiCA0IkRorcPrXT7S4r8Oq+D51rG+tv4A6seKACHfRKK6TSy0
UIgTPYuHHAFr9BVag48ZmrQWfAAThI1/5jjjeNuee+bIEo/Px9TD9NJO1QmBzx4uAk5kSo66guxE
EPIa1Sv7YRj4os7+89x+VJc/mnfhDefzU33YmPB4Gi7w0n5h5Mv5l1OLA1M67/8ApqAo572BTmzO
7dcJuWPZ6BUxPytF5Fzp/02JiFFWiQrmBP6a2z0EaEaRD6CSNSjsNZJtI3N68+2KVwUCM+WuuaAX
S87ou5QqQ0KwTGZ3SLPDILrvOsAEGkF7Bts/2o6EREYLpFlc7DSJymrhCkHIrmKWPrdrL27BfoZq
GxxiM7ReZRqVDu928yoQiDnVyHOZgqOzkiR8fNcl0jkGTnZKdAmnYk33VsdcPOHWRgPFdUEL+bz7
fUmRW62Dcoy5HPoVBAFgeWJ3PpcUR5bWC25rxAl2ImVi7GXgw0bVGlBqlTGzJ2P1yg4hGtTwdGxu
ks4xHsi2XaC6Xt/ggNn7lECm4ga4FZgjEzRZ4N/wkm+tMOKaSi64SCkljKK0e0038jFvM4x1DE9T
9ekBuPhtAKi1vT0z6JryWFjgS9ff7x8TD12P4JTzhDl/oGtTgeikQnB3vLE3n/JZZq85Ix3PawJn
6iNb5V31eJv05P37wyD+qevhALHb+gwQS5ULcR8BLT+eVP3N2VyvItS0RIP3xfjwATyIcPjM67V0
PSmoHxG3yPSC73Xk7pboVFLnTOJQ10QKNsj2WBm6wcr4FPk+lmmLBL2ndtutzLC4uy/W61uGRV1Y
ZxAqoVtrNaAr0wFgoMYEl/vpxQA9btbQBSyNW5CK3J6RJ/V4E3aHrni8WTCYOK7WWP5k70M6IyEC
NSgLIWVYSl3j8BuykvPJVsO7tBA2xgSP1BfbWFb4B3lljzQxRINCSiAqdr3pqOo/iupClPIC4GOy
ikYSrtLpCAz1tOSUpIFievMB12Ikjmi/7hlx9qKDtKcWeREE+a9TNBzOw3U27XnddT7obwqkLWMy
kii11TrqmAJSXkBVoVMbWS047DuLMY6vbXjD898IrwLz4dSHGzsp4eDHifxnSfgnmRYImgExCam4
B7JsQNSiN+9UU2hnBogUkfj3hiOO57xojxEmEy7yf8uV+et7R/mg42vN+1PnqHPKp/6HymXIl6CX
yIis80jKBduZ0S08eYHyIhtGnP6kkIFTCuK3xKkNCVH7xqq6Yc2hfiALyQWrOrDn4fxVutq2bQTc
5prgVR2cHf+OyfTHjOqAoLpAd2R5s5cyMBKL8Y8WmrIUWZHs4HH6+VVzG2OIybGYaF5ahGRMuH9s
EIoJOtFVLZfIrnk2E0VQ8IjagdUrfclwetgC35/96UFTpUl/XuLgcWqOUjRSzDwLWclSsZnXYZEK
BfOYqRY3z3++pK7XbOET77+5e29xrh/NKroFrXXaeupIlXSQjP/3RoKK7Qnr0iZUym5SyGQxn7A4
F2BN6qRuBcgN84yyCGtEnZ3Epgfr2TybmCarpi/SfSKXkdbDuYkTh/CBLZaPRRyPhsYn9JrhpMh7
co8dGwXa37PXWIzGaFY+d0AQsGdJgwUB4faARXTk09U5W4dTcnpkFp4bbKeC4FoXsOuwAU1B+2mx
3EPZlxgwvfH3/zTLCniuMK+iNWvYMTY5cbM87dRaBSHUPam77AQ0th16TDtSD1xmkFqbZWtzsuuA
2ebOzkY2c5RDtuPpNmEqZU2uq/mDb8RMAa5T8wC2kUth/sVf5+uC0R5ubjbd8AL47jmVwfrG/qwd
7fWxd5J+IsR6EQxUGey6j23xfPGfc1Hqgvz4NIZrmCB/iBr+Qbp9MKJvRELu86ckxxzH3RXDc3Rk
ezjux17aTFk5qJoPwHTu4pmqbN3PdXD/tUx9d/G9S3lM872msC/p7vFjChue5QOcLPmcQ2FGmKIK
r8YueSV10dlvG8VOhytG297zNKnOursoh7GSJvqE6FPScse7PuBoBmqvyv5dG1p8cbcAlmTcj4EI
ahvZZPpRbjOgwlwlbFEXmHoKvig0fFIueLfnobizKLmgAWyICJ75jt/gRhmlWU0It/xZ5yCSetLZ
C1r8Jqq+iVyfeTbYUyi/D5MQXv7t+EHcWP/PktpCq87QlcUFEq6rhDm+E61Quv5bz7VydO+X3LMo
3SayZIAHOj4fYVP4Uv/KnhHLn6R4thlfd5onoKbMwUJWPpTijr0m3dtz6tBhnFy1qVJnyjkZbePm
jxgprp+H163c/BQ2YRLNrDzmAAyMUwgGD4rUX1Kf3/JQQLwMatmHrqXf9FlY7Esv980i1R2O165J
XWr79x3PQuQkpcdIuXt1h6XbrDEASYTCy9zQof9zes6Y3eleHb0MmF1+HD8Ng/7ndiRKVU2e2nGT
gweMM36r9LXol1YM8bi2nJ5WZPh6cfqcrHRHX6lt5nbAQrsAHtgvCK8AudZ6yOVXD+0AoXEQSTQJ
SoGAdxh2SMTZ61no/ATODR2KK7JQ4+j1DIz70+xC1MQ8L0JWEZVXXIG1vJtinC5J/Jck4TZmtS60
ThKdG+MfCQz51TNebDbP7qKVM+PcD9oAt3vTpMrzQE2zTZyhpibxZaALfwwqIBzwKGvmNi4QuUnw
178Qp89uzwDIvCxPY92aeV9OFgQBftZlUNI5/k/EaOtdXj4MZNMp+EQQh37Jsp9iSSyJItQ6Xoyl
0HrQDWdmphFz/92n9VzIAPs/4OEBQzOq8OOjHmkgWdYvhaUsqfpz2GIzrl8BueLMV1b9P8sU3VtP
flTlKxY6L0B/wMSVcbifCDjNMXabfqfOmRfd1WFV7SZlgTVIBcHLd0gQsRuL9Mya7dNMkzocU/Xe
KvolVoesmpuazOhc9+4WhwFqpXTjnImMA67wIz3SsfH4de4j3VQbxsUhd1Sp9CngsHt81pmo0cSg
KVljIelCdFUhqDfjE0di08G0sfOYQqz77vazQxbTdWRI2JZGX98ey8HDuw9KXv9s5MVKlEzZY3vA
mc3Fb4qfCXQSCn3M57TUn63s6oVx44goVs5tluxB+XHGGw5/16/I1RrVi11MIFWMrpyONJb/DuQp
ODrx8HBmoxm5ydST3lHA6t7QqC4ielIO/o3hUxkTQ22mQVV/FblYSHlDkVVcud7bCqGy0VzsM2JX
4TdNrHQQrqg/rQ15nG2GL6GgO7iqZBoNjXJWDupStjrdvyDHevLalFe7xMFaMTwvLAC3hR4VBp4y
mon6fIZXnsdJwJSupofG1ulp8suAu44s94704wJ3nJI/wIIocmHPBZLVQj6foMBL5qCppzWLrnXv
Zx8gKgjWuxbiEcGlenuO2SdDntj8w1VYsMpPaB1ZSt0a6pMk2t17/GD1WtETsYb/1BzsMza9g7w5
47/5jfNYre6MPfLjoJefPB3rWnM9SL/9AwqJZnsV++vaPbzE/ElTbPwGzfEx4mq/fgfKOeVfoqJN
JBaLiLt08iHNkwO2mro8RshP8A2xrwQZ9/c/2xNVJ3VrDA4dPwWk3WUSbD++UkgXjbPqCkhrc3jm
QR+qLmo7BlMAMR+klTXQQDRXnYbTJI3Br4XGbcwvtc1jjhPfZsx64SOrRqv4xtW1ANS5x/aP3Uay
GaYXaMwkFfH+SROoMj5ZL22BXCwRFUaAI4l5N/JjCqhotlamnE/lZSMEow567AJMd2fmNhiRINeW
2emKs3OYJWLrz/NABkvL5Rd5+x8qVREnPwuCd24C3CepFRNAElXV8Cf6YfX3PDFGA0Jn0M0kYCcE
0NSqUbnlzZermFT3d9JrzIjH6p1qCjnZCdON7ksahTQwDpxqmhROgCdFXS//uUGD5SFVOyrx/W82
anXJulEarnc/TMljOnvSBj3YtVnBAodR6NNWkCx1xl+1aEU6k0rYpuGU4/iBdaf79p6FLyyp4dZL
SIUAz4/XGc4qVJINWRyCokVmBZN2l9ihR5A4zMqIP/5J50rjtlRcH4D8CSJ8oYaEzDZxWShKhJKL
5EP0w9rnuFB2qfHmqEp725ywHgv7Sq2DyuNe/EWhcUCcD1YFEg7TDAHcEd70bnWXv4EaWIRXhrSN
x/qezADxP9TvWxN6ysfJni8046Dk2X3EzudhY7WJNpds08dVp3BmgmMHs5qyhKzd1pALN1YGQlTt
fvzah8vc7jhl4LmVdinXI9Vp32IrpjtwlosnJhBkSPr3ssrYwRD7iEQM6Aiu2oXIO14ghBzTxSrO
5/55Cj38P4viyt1oV4nqEIK2F3pc2amY78ao8FQmfcgvEZw1mJdnnPVml47mMXDxim8v6qFBC2Ah
qjc+OvAZs5E9nmWUCIbyx7ZdImWWEeC2vtm9DeGzDijgirfoSzjG/ddk7IClhHdYpGnpblLfYftx
E0Tg1g5R0Ua7wiwIxVoy6dNRv523nj5zl1IEXXQZEtbI/zsa33W9YSClOA+5h77FSZbeeEYSmjy0
NVFq3V2k7jfWxj5LdnVxIGqgLXUA/YVEmMiP3ePpN8ipaGN9iD5KYHLZ7fByz7gwQBPiLzpjhv9G
5t9lzdoWmivwhaz+5kG4biTnAVqFfMuyJDtDhhEFnCLZS4DZMhXsUR3PceXGWFzwrDvkZn9QWeHX
a31fiz2g6t/U0vk7f0QeTECqLhNMDjixTp4qFNEFsMyaB7i4l7Quu57nDGbemaDP+bumgt/oD/lB
nyXsXZV9yEhdnX1M2fTM4ajgHSIIZWVUV7cI+Z1tg7MpRyui4nWDco7siaGE1ybgNUgWcSnByXyN
U8NWQC/MyD/WE2VYBWWvlxL2yuPqQJhVkc0MDMghSHCaY+8iCgqEsl23V7RsjRIDKXhf+u+sl6+3
E9seRDAUD6jqzG7j1CgxT7Rbp53jX9kjY41b/5yaQXmvG4qVpgHpkprkIoa/AvkB6JsqJ7e63mCR
DbRS+RuW3w3asrK5TklzkQt61C3+wXrTxuF7feV8KvntYpX0LACTEneeIksVt8mGoHXbkh2fnJgf
jGXhAqRDyk5TUFj2vvgZqYy5s4oslNLKuqOOLCaZUANHUr9sG/7YGVL0Qzz3/zkurc3bgSye9Lx9
rvs5zOU2+nizroWSE7D9Iu7jmMIcpwI+kokRg5sMgtP1frMYuSwqrYMG1h3/kFzeRgPs1IozBFw0
hncfjUiuFlpIU0a3bsnG7ESuszA8FDKy0EgZTPw89KOPDetgWyNuGKnaKJrrvwzPTC4c/kdTP26/
KVnefGY1gIk+yw0TBaeJ5SsL84vU/nAlWI7ZtbUGkiMxzLTXJSUYICmOlhzxurv5t7zUl+Mh6L2o
929RwFc9lzYtL7fQ75zP66k8+Q9W6dbWh9gHyfT2tWVepBP8PFtaGt8JRdGBJ7cBLQm4hHtLFTgo
C+MeJdgUT3Nq2yz86ppyb4H/K5v4ZZafodczjBn4bdfHQQlTYMxgpMK4nyP7MZU0YbNYJd+3z7z1
G7CYJUlaMP5/mGADsVqi/+uwc4ct7EZwhNobH9hVsVsWGETM6QaV6SNzKteouPqBZkVt1sDzom8t
d+ml7WWqljlwcJsKGcFo1FdcK/ZDIs4z5WcSHhEd4Zc9PRLM580xOVH5iWGqkfIGkq10658kypdg
AW/61tTQ9Kw1sHbSUJ4LLWUv23LKYE6o9pVPS7SyQtRTPJ+77fNj0LR16R6l4iLpFHXvbI9x2sZb
imsOJhnQT5b7zt/fHT8UJo5CKMyMhZqwx9A1fMy11C439k+7NthLP6m3uAkDgG/4or/goCNo6mlu
A5bYhyK1MdsBpUl8ErWYdYaHsgZaU6luFkx6SKgqq592KCkVdZd++aacYh+wV+vwAp3d1W7Sg97b
hxIL5/Sh2A4rqrOTy3RMeY++yOauuAFJyY0De0Ds+pZN3l54+EvXyvU5CbtAWQ79yX9qnyhw/WTz
FTC2QYJEsN+vQoGt3mI5SDEwL4kxEGQP983ctPlSmCZRB4v0roLSaQ7ZokWD0A/AbZBHtBgtAxx8
Ofz6pV8Wjx/TLl1S6NDTx/KlBnIiu3aJRsAbQpl4tlpDhjbQalR7Zpc+X3ax16OVISG4ggyinYLy
gTzOeTlZle3CGjv0cGrDAMlS8gfHkgN29wd0yzJ1pVVvnn7bZij+dbwSWCuNMW7C8usIRehp4tpe
F2eTQhElC0oYqTxnUB5Zbl96fCFtz19+mv2lKW9fOrxkhF5UFUdCL3v8pRhQMub7qCa6aRJEpVrM
DNEQpZAA1Ddwjf0CwMa+j01rlE0e2zx1gRE//bl92jhj+mqKMClI77S3X60A4RXNSvcL/PzALUem
L8XKssRi5FMhyWYtsZvpP3RXkcYYuqm2M62QT046IL6rqrYczx2CWgqAYGowspnO6IE9F8zBeERn
9j5oKs8rpwbhfKk6IX77XKFKqHFmV22uv5lvbICCh2jUD8eElxEA/eOk6U07bqPt4KA+Ij2CkfFr
IqE3L8yw+DsdkaWcMAmzldWb0l0YsxWSAeAD2U/4nNqrGk+y8B49NiNTeBdaeB8zEDeabzIK/7yq
JyCR3kPyqiM5k3+KddmFNNax0yTl+6Dl4IQQV+0BOU6fIdYTk/cuvXfwyVYV7pe8rpkpvtSdvDlH
NfB8IX926QFkicQHNFjjWvRZxatwSYqoCAs2IJK8LcjaqqBwt6UrbpFUkEWnVFunMEjv7tlDd5GZ
D/rKrVCU4i1PZ/YOKdLI6Z1w3gcDq0w3th1KOjVtvXIv0ry50WrnuDqwBmRRfNhiOHsl/FrO834Z
m2NoxfZLDnfuh/YNQOB/dkfRxIqYdy7BSSmLxs/gYNQTLpFC3Y5yypVgMRJ5pZ9eg5/unrV/f2H5
b8UkrigWuTHFfcsxAdxLymjt8N2/DbS+F+4sfek9jwzGLDFU4IhbsG4CeOTVZWJYPFNBseGNrgLv
y9d+vk9A7go1N+bdA4zmTPFLnXdeXHyeJqxHkbbM6weRbgDzEZvH44sPu2jo92cZXCH1mw6tIZPb
6w6pjTKsB2J9f70OGPYm9GIi/0X6WcCk0ut50fKXZKqs2CPMXqnyeRWJM0GVJ549vv1F1OXOqvwv
zi+YRevTVYebxByOAnhIhcjsJDyWAEnhRLIAtsxSRRD2vcp0q342DWd1U1kn+18/EeDneJQsqPPS
+3R1zYUpTXhVkwwWQSmMgzFPQD98NnpjI/Mp/auV3eDpaan6WkYjwfsTzcQQCGS1tyG84pD4itRU
+2u6F7f6FHsMcdQfow2BKHqq4LDiEeHogsuhfIEP1yu4HZshU2642d++m4Nmwbm1jPFgfR+7a9l3
u9ZWLyz/LYqj7rTRBkSUfjTxAdiE/9EDVs7cKcNz3F5F4vKae2rlVi7eIuSbB+PMQ7EVuOoj0z8s
I6OY0DJvkt9CO9+vfP6hYI5OaAYXkaeRSTLCEUQpITuax7V6nqMfO8Qtk65z68UIeAwsoE2JiuhZ
HVPIZB8Jw2a/MY64D7r3QbFnIUgDnZnEr5HWr8xo7+8+VgNXFY54bt0Kxk7r+qlgPwTm8KVrD8+F
HF41OSZrEyHHjXfD35L0m/0AFFS2T5WZP/a+/EyDCu0bz/rQOvNQPFEk1itbdCFPS40Ysp8OtRtd
jRRR8CF3ASjziCdoqwTiFeYVIzI0CGeBQ4T8uRAHbKS+Jy6HE4BWdK0X8soz+t/S7lmkqvqtnZUf
68GTHPo+I9/HyBmLdfflBoqBNQa9ovSRzdKpX+j3THR/+LPlAux1d8SFMeCtJhnX9ZaXqTDtTxKG
yjtyNcW07nV5SELYD5ZxHpwbpGAg9Kt7wWC4oFS81XoD5WI2TTbEhBsW4R6F6o0od3vPbsWctfeI
I5zBH9yhe8E1cjiQvaBJ/ECLnDfqW01lX1LYMjJxVygYvLQ5GT9jmv0ftt4xpHNPZFuwLj5Oy8VN
BDbF5U1GAv8fFpp97FRGoYUAT4OvMPWtBsg5p6QelfqUE66/WQuiKfmSdwYRLElkjLAyWg77GDAp
eK8686l1CT74mNZsqcJUptErkBiCL+cNYZHWbwAARX2ltE5Sz4P5+0lzdDIlFZkubk5ta9VIjQQe
sucbLcLpyHn6fVa0ik6Sxd67/lu4uiWWgr3mS3fce1n4gDFuNPux14j7WWPWQxPWKpAdrrvj6+Gb
zDYc4UX9lbmOFPPj1KDOmXS09TTa5aq8dP72u/kIkosfUNJBTyoKji7gKa1TKaAySxzuQgpzLTCO
Yh0wW7o59iJ3OBom+Tl/uOESKpluZQRDRCdz6N4jVzkSb+11COgdb2rFKHghkwjAQ5YmjLI5+JKR
jMCXnwVXwzntZI1PzTznP6lE1cjWuPE+STd+sOpnjUkfg1UQV+Ut27PhC8uagVshCLP1lscIBLbF
34iAJBh0LbNE1DqVofMspZihNs1jyRNrvxjeSPUNp4zALwmUSPMuZjPWW5oV02nf2MaVM6ESrp8o
P24VbclV3XhRRyAdAi0eI94NlV6WGJprEbWswVewZHmy/foHhzbwMbzeSUnpUWVNFyunMFphqX+5
2mxpIBRIb+aSYdPYNpd8tBUMoIGgtha4AWzXNqm/IDLHO6AE9DL12MZVXD9wXNH1wyhgDkPUaiE6
WR84IiUIy7mCVVrf3ZXzUXXcntQmemkCgOuOcIEqtadQhOv77UOsLOrMPV4cn9F25PD65m0QZoPs
0gqZKODMIxe/hCw7RAym9FmT2zH6RRc/li1yhIkXLxxbtYZl1zkoVI6SeWGCwrvwDoBFhAdLTYME
FRjDh5q1/kFU5gNTWpQu9tRsr2IN1B/MYZ18U4VWih3eh6HHJLHVovNUfcHtxcQtKNakN8KQw6qo
sKb5NVDFgb4aiGlrtE7IwSy8qM2ylUG2BjKmsIaSTx72UAWauNl4Z9z/QQYLX1QERa/rVPebWsVj
9urfe1Gp4C+57u9Bdhm87yEWvCtIA1Ca2z0oyaqNP26cZ1KWuio+jLIvnIDgHIhs4cyde9VoU580
5K9xzWg6Dxig23hwRusJN0tL4uci8ODc2grZoYb5G6JvWxRcC0k8GhNhKPO+6QCjNXe3Rfx8ER87
E8S15enspnEwCvq6HmqMxUMoAFlJcVNw9rfdJfoOBb8xF3ZhnM9uAHGdv8Rs4LIQZbQ7lIltme+P
7RXLHUkiG/bqGGuC7kp4MTtYCl1NK/iaX5zDpZoXBw+SA0PlVTqA4TIu7gqdXnLJeb4WcgaQvkuF
8bdEQL+IIGxVtWEcUej8VOogJ8ZPK7JLG0V8rSl5rvhLU8X5o1zogup+wiahkGQhzkg3obHLOJhL
M/fFf3VE/JmvJPbkLOnsX2XO6f/F0t8uh/+914VEDIu6cUHlZ52tAzoa4teMJSFifvchNBqqZfH/
Jla99e0ZoED0gEuWUpEp200tLYrZBfkNSxZFVA4r2HP+L5M1BQ+d/uDagETdaXtnWjcNyGEzMSdY
Hhwy2fUd9BvbBTxiEOwAy1dI2dFPUfWrkRosSO09p+LZ/bEjHABxIj6XD0NdZq0b0Z0Q62FIQXD9
IGq2pK2T7nvYu5kOfQiVc6pdMR2vhu9/GtBXrzMINRpsGOyzEbNXW1psVNIykF5II5/wQWkIIOAF
2GSCsrALfp5a6WFckOyJ0SvlhQNIb6qnsdC4MkAby408fMlyVIm8oKhDthqqWcL+EOWHYd7eHea+
PAXYf+6yZH1d37Qb4MpGfErGh/HSqUTzjrgDgU5A1Bv8DW/nmhuCW1LjuEce+ey/pQcQnuIwhWJK
YjkDdRTwqYXX6gCgIyBSzdNJnxFF8bod5K0gflIQ1dFOAF4ysV4LfYNiWkTMx7zR1h2jSEgNWfDk
pF+UhGoFW9V7USZ52miUs1vHsQNb2SrnV/MZCbWwoG824FO0bokcsmmrMJWXS6fE3neKhFkfo5KJ
VN7CexDrerDANfAVFsdlnb/3Uns439YgTv5hX8SRKqCdPG2kOdPE4OBwG1nXXkd1F7ecP/uek4D/
2Ww8X2UxaYNrPbJ1+h1zNInQuML35aTohT+6nNIFQzotqbaG8H+diGbkmpsNvgto3DQT/7/4zh/e
HRKD/WxxiMR6Q3q7DL3290nv603X6dKBlknWY58O+7osGzjv8Y9AZ6XWHelfdb1TwnpnLv8FzBTB
TIx2wuztnOZsl15uMPslQwYrDWuNwER6gAiOCO6vBwsEDvnzYmQlzRrVSApXLVDDTbrDGWA1K0jO
myIodzXfeVDlWyrwXTlW8lYuiYE9TcW8PA7kjkopzs0r800j3giuOcCj6tiPSNZpmdPc1yrw+lSw
3B0xX1bQ8W4f+KOk8iDqcVqlSogbddcgXcqNkjZvXiNEYXIvDagZivYWp+d7oFXWJoNfIohQRrX5
OCa3dgYX/+9ke4HdzU1QlciR97WF5FRMKkV5hhR3qLKp0He0OkKyUjTJ9D03A1n0MlYLRJGSkENi
FEOSwEYfOvhLQEDe0CpBQunGWwrLWhJ67LmW6DwlTZ1AYU058adHK26aaqv8l+AHl2EppjYh+Xbc
JtlQjZFrwlZDw+olRRoS546uXav+0KSBP2pT+Pd5HbR72nxi5m1Rd4V4FCQn0evadAcucclPAofk
ohFNpd1o9xP/7XRlwm6W/fFu7KGaRBV8lGMUzHEPUHaQcfqh9spg1MfBFi1mRyW3MHKFu4cfyW8M
UTUVi5R1UyiKnULkOemnGJh/lazcbCuGA+uB3dqSLDUrAh05l2KnY0VXrJDjW66OQC+0mUndx+1+
wAKVCFdv0gb/JuD1hS++paeDeNKy0llyqLsmYzGCPqRqfGs9sE6O0QXI9HPYB0SQ6OIn+B/C+hDw
IKPGUsRRm1pVC0ayIRiD3dWEXbEgETLWmKwGNdGRLvxvMZoOjcGnVlsm8xjpGu2/re3qhHZX6uPt
QuBKo7IsgFhwDDOLoHVWQql0NfQ0Bjyu8vTjNBtYXHrXGuW5RYnzy870CL54liP877suRmfZ5qkW
Zh1byiJ76LeXy61I8q9nYHj2wCMAvTPyBvLm4yPPPbXucYDbVaAZlKDqkl4QKO29S3b2bNUstDB+
uSANSmeTsNxioOxBtTO+I1sQUdBiuJwaQGZ7NT4p7/K/2PQKSxmpWSxcVpdoxQuFlMrof4Cn14cr
7CA7uBu1D3sd7+XiBg4XPbAZn01TtBIkkeMExz4JWfKFGzaSH+KKNC1M5cnn40TnBPNfObQFjDMr
WQuRotBg0g/1mKREf+IUxUmQrkHLku99ZpdNyeqIKhNXS11Ey/7RS4+GXoB5tuFJWBhaNjonzPaO
OhIE/rr8oZ6diuTIn7XetULUqFCRacb7bhPr8GPKfgpF9ZtCCFmeut9c1Il1WSq2PsFrbprgrnv/
sp4uzQJMOIaCGpwkBgAczPpCY0+wzEHRmGMdIhMguYQ7dtYg0E5ZPvUKz+WRWFYUmnVylmSpMVCN
pgjxFKIACD1x+oLD4Ed4osVuhK4LvtthjWdDszrW2+mxl+EnjXYmyBgd56gV8vijWy4FmZ6hnfVz
57Kh7uM2h4BQZleWcvnwncCSffXGl0B+T7jIWk6DBe5hdnB9Z3C6gMFhgVy5nEjdLrP4ibQXukEC
qP7nthUonI1RlLuQtnpzTTo7lXywfgcSJrOChQ80QGYAq5EjFhIDe54NO1ihgPHGeKGvt4qdqdAH
hHjGbGUJq35qnbUb37fPxpreaMKM1yD927sfgzOdnuYHAgxIvwEazfx5ETdVrhOCxLjWpAE011iD
zdqzJyaRciZXyUxSG4+QUoCyD08ATph/h6UYGG7R+UnuMHfARUJ8Tod/mMSwkURa9ZU/KL5SMpb/
eke5A9Pn12tJ//YpbtFvMaFtrIVQUdf2pHjbgOXbCJMj0Sc2hNCmAQcNvKH4Hp7XNJkqVQOQ30yd
oDrK3cXij1hG7GH/p5HfWApXj1cuIz3a4vTZal0i7JysbamCLX09bm3DDhno2WHrkjahu6gKFrs8
l+IL0G4z2csgRmSWo61uaHhWStup5VctnK4l0rP1tCNOPTyUEv2QsveJwcNbLam7jvI4kEzblS8C
HKMX74dWuIZQo5olme4Vtcc9OWo7CqMWpW269VxJQxAtDmZttZbEHqyN5fJ0gBhy2htm13uxNrGe
z7rvNEn4x0xg3sF3Pi2LUTRY8xFTQGgiORdtXSfr8k7HaC2IwyDWa+L6Sm9JlkT4RnhFKG0QUXc3
u7sCi9Qp2/4+whpAvsFHrbctEHVMcAAaSmWEPAaZ3KIz2kruR+BgipCivHhK0hX4X1QT3jE2HPtY
6n71fhLjMu/pfYSqmkXwcsxloMCXKNxCAg+iJUHzgR0e8f/oByL2s3XBoM3Xow3dS9THqedi5p2F
eIGlc1amo42SySTAG0uUKbVVSSFeMD/a6lztuy9x6UVJQl58Ei1L9RSAmefNPnKDrtdS1M+VvwJN
yA/sXbpvNodkYpqfCIfspVQSjxXUEYLY81XAn9v8dT8NExxtBM2dsjRv5hoG43xbT0YwXw5OC+EW
zrLPhv5IcB/EnXrpvTurp8aKzH6AS2gl9x7uE6RF5mK2fAn9JrvHt4xJ0C30vzmzdenTT9w5wqD4
8E3FU8QAgoeL7wNE+DC+4zIZDS/uPuKX0DWBrInFVRcbJaUsp5IXRFU2kPg9Zte6EHtMZMh2b0pS
p4ni5x9w6VpqOaYsiq1wCJDKZiOpVgcuT72Fg21rayXMzJrtwZbUBv90cfRUybJXw77eAcfrOQYZ
fZrJO6dym1DIbsf2VJlXGsZHf9+toqAz8tZ7afPNMvelcnVVaIpnq9qDEOzb+InHJF0F8GfkcN6d
e77V5HX/jPdG1nMoCGHNob0IKGfy9NMg5wVpX6oXkZ4mZwyuBi2x9OXFv85bgzcdSrhZSrrznaG+
ct12oCflKz7OSzwYGYgBmDF9nRvLZgb5/rWDd+a0Bs18NlNSJX7aCTBCYSNWZms57DIUO7uZyP0R
OfFKnhm3MChkst+1lR/galT8R/5DuDbHJy1UCWNFFtK0bayroX5uLqMgWlsJrL1Hehgrvl+eNbIZ
spb6hvEuPXKtBzWc48+BYjhNS7RvPr2VBgP397mHPo7YDiCYHopbOahA2ZPF2niMZ6SjVSWGVmCa
4HmBcgRBN0KcZ5UX2xu6cYg/cLf5e01g7aTw8Wg3ec49QG780M+6iQu3SXj5VqySI2QQ7nlb9QCT
Tq5E3ZHeBo6WAa4aH5/6urtPJNUbQgJ4gNNthFi5f2F3wx650/d1k731/1GOKsRaNXaUrMc4Ifov
GX5sKVZvdpGB+uN8iNokiLIWCo5JpqVkFoWNbaalNvuRJz23To/ORuLb04XHjruGQBo6kTFEIZpA
vzsd2VS/OyXI3hCho2Hwdke8yM5+9DfExdEXFSSI0zxOAmNiuHtkINwmWrBMgvNR2rHSQzoiyuhD
leEdZkR6RnFt9LsdjUiigLCu5QkOVzA88ZFOot+GuaNmOmdv+MKd0ld/kU2hG8w0ghLnt/D9CrRF
vIRFOgxalldZj+JRMlad0hP9j/G8fFH+uTyjrQbN7U7mSD/CPql+a4Xd8ADcQolqOi4uFaYbwTJ4
jcrzovrCW2GEhyt4vS8OOwBtbUAM2zmO6XJ9lpxIw3HavV+81rcxjGrYyGvBZlqDj63JOjoXsm1E
uAgFtHpCbx+eXId3jEwPUXkIZPcN5MX+MbYxkq/ws+NQRkMBhDpT1oFmbJ0mD7SytEmW6fvrx5vo
8B1klW1rIHVks1rDM8+yGVtJ5HTjiaV6FspBatOWJhblhm3OmWmkjto3Gtb4pFCF4G+uYISDQwJ3
XCSVRKOf4l5Y9TSSV6e+NCGMXxvYQeyo2UOGEMpl1m62ZRU/wrm/Ys6n4tpz7X3iEmfi5jfr8cnw
sZpZB63GcXZPKpx2ZJ5EwpSJ7V+A3ivy5yR1+aKy+xY1ZfGoxAtOqo7BG8KOJ7wuijQHwfod3hhg
6r/afrhaj07QSQWL2BftdNuTSnmYrKexyRjNZkEvUiDBsV4qFMvRW5jnyY2nHtgUz0NTdbpvWRLo
sDSHyMI6h+/8wQRSFi2FutRwYNH+wbbcjIBT3gE3Imm4DoTWZJX3o4+6v6JH+l9xB2Ow30EKwiyL
NuHNREO5P1lXtufN0gH60ZDmckqpjlTFf+IkKhw+rEkHNQlstpWT8fEZDcXiQCiA6KfjUP881Hh8
HUlDqEoLbrDMassWUFMecsjR1OO7nqedNAy3sEu3+YsCmqbe9y8zvDJ2iKoLnpoFzg6mPQvwEsVf
l0Zpt3FaPWLHnGAgxpU3G74rHBuA6DQxt0sPIv58pqyH6OhM0PiPLcGpjpLLJJJwFF0oNbx61ZOk
E6iakdRr+x/odkGuCFUj0kPzLQMpbrlMZVmpqA34tRIVcVsXhCRVnhye3lDRnhUzg0+n85bK7i0q
ogEZRQ6J4uh19p9OW1aTyeeZ8SkkzqCMVeGjmcFCqvcf3q1uL6sGUGdb24v/EM86ckUIn+xM+XPN
V/QdVBd8ZwC9GZ+b4wgbE34xljNyBQt103E9WoKpW29PGNcVT6WrHpFMUbtJWXvZ65q1FPgwMQ+n
LzLzaE/qx3Gh34sQKgLQjkUHIYS39wUgVFsvrmm1ktGepL6F5tqEO3ZaVDaGml8TUAWHX7xdyO+S
vR/Y3kYyKm9WkAQYkOhaDmuQBr/dFQiEFkIs4XDCOxzU2COm0vTcsuDtCMC3OA4MXe3vuzaXN1Hk
DbS0mbbzzS0uieF7j06jws8HsP89f4YMazmckxzReroSkkrcL+Sbe4Lngj7djemz94MxI6t28DTG
5cz0q8ctAPEAdabOgNlUyTMgr+3YHPASEZTgcYoIySA+PwE5Mjyx77WKMOt5XXqO5nr+/0A4N6kX
RFqlLa4Kars7Knc8cIIY0G6uWgHB5X/nCRd/p59O+hH87E2KqxD2BZKaD6EYgp+WkQTqcTxjHQof
zdQ+iG2CP9N20WhRAfU+dDWt6DJ9pdidCLPxLq0c2XSTYOEFaODzufXHxaoVzZaAu6FHGU/DK+cV
JvlejJunIDNVViI8iGW5OS16bAkNMHowguqyHdxnsaQl2Aq3aGVFT8cv287KNlFh+wkiQMJHowsB
b6yw0tlDzZMwOfym52f8U6vPh/PIl9Rns3G7cBedK1STHNs2+G1LAF94PqNRJUciddXL5To07HaY
hstHxaE6YlPtf2Xj9utbanLykfUEp/QTMc6sbAu7sKUhcg/MGADc72uSt7vhLf44S7g2UXkZgY5G
dPsGyKwuwtOa+DE7bxXBZIp4lGbizpEXOoIcJRA1Xsy0jPK53FaEhK27V120S8ucO3Xoce5YxFyw
F/jQ3cGXIPloMvQmMH4/FfG6tkjP/s+sPl4tkWGzNIGnKFobzhwQtjegsCUdgs7l7t44JxMi2lVP
HM9Q8lT/rexhgYkA7t3OMTRCpXjIXk1TTG2rcUtZCQqi7JBX0d8Zf4/2VnpOeuuQo9/z/3nsSWVk
+CzaJIJKcy/BO2+V5jLXEqoA8NEtLcF0/G64UX+1r+mifn+bLemxOJvIdQ7pgefQ/PEzNVFZnXHW
D7VOsz9iFvr37COX8sT/bdWU4Pqy0CISzHuvAb9DI16DIZ409+inMXQUkNKrC4HG89fspP9G0NTk
E1jaFqgFKigtFZaABeg+mIH3knw7ZLkujIL/MX+DXmxz7DdCBF2RynB7URqD7ULacps7sCABQY8n
diXXKrjjAyi2psT1Db8s4R0ovbHIQQmuZCMgLPiaqag6mDSGGXlpUz56y4Imdpo30nn52LqRWzZA
/l2fTOYfo4JIABpnFZzN33nzwDyRrVpuAarvl9CIxGBdJOFo0eQJ65KuDv3d5Q8eQ7ef0EdjJkSs
/pF5kSUveTW2lagL9H5Q+C9gFrg3uOIw4G6fdfPHfVEzBNLzcJYfcTF7FOl/2++nvUxXXSNvSy92
2ZaOxRb8+DP6Wrc5s8X9Yz0RbveliJeXklUpHzB8mx9Egu8NfzDl4m6Kr881rz8W3kS04HyUVFhi
4VobiK5VrVLbjUBMf2Rbm37krQ+2/yrqHWdV8wZR2wdDqjbpiRtzNTcfWnCegJlSaqdYywYDNqe9
xwB0anZfxuPrO/ehUXmKpn6XhJ+UD05hYuePBp1ljiYl8QMP1VXk1c93ZTtahfh42ksYCW2N4RNA
Iq2kcmK+iopaBf7rs5KIqjzy0QyJ3eSHY1lM1LdFIdvdYp9uMC/V2JKGQAxB/l5NJbzxlla8dakD
5RRwPMA8LycvOFSHxHl130LrWh8jEh1VzPA6pVSj3AE+jZQ7jI+cmdPloXsjj8rG9UwEUNWWd+wb
w7R8pYp0UTbpA5ApKRJQhtdKjz0A+p1sy/v5LgRCTpU9s8QpPjzrbE5rs3tlgUjz2BlXju2BSoY3
443+z9V2oQ5lHaQaDB3JZKYH5h2GOYh2+y8v69JE5KAqbtuStdBjytmy1QZOnDMJJ8bn9VJbiWOJ
VlD7jY57RAfkbsTYVpo88VQQN6bVlESfvJbLYA1yzAY83VvfRtDxnK8VtpoW2eOFnLF+dlKtgfPe
qjVQ+pb1LvD8HB/3DbRADJQxoNjeEYCMZV3Sb45Bti84xQcSeZyZHYLKROaJ5IygES2iV8+lpz83
2mLXaNUKM2400GmQ/gowvIyewkVxIUXkWQjGVaNTW18ZgW5qM35xBy+AvRfBJveyEqqF3gXCDUTc
J0P2eopjUp6XUPl19Wsa0j6jjN/DLlWK9NJ+0E0vnL8tHeLcHB8pWf8QLVroYPmHWd7IJU2HJ9X3
tGQ9PpFAcv7LeVUtrwL1/9JqbhgcaHjA8iOZcWkRUjzQKt/qFe1mvPw4UJqcqYkEsbpT18ruCZL4
ZSs5C//W0k1YIpn0In9axXPaNpRY2UMT+OH12eqb32CrhpBR/E8DZaxh4DPtB/Jl4/niIrV7H8qH
mrjo+1/onCl7XH00OIk947KY7JRgDrMnKY6JsVOhj16gWLGy5W/4J7FxPnxlRhtjpxtTn0iMrC7H
EJGE3oxD5Mgz/mFjWiNf7+jzkRZXCaZ46kK/V0grcnwRXJDjOBMaaak+epGeSsa+QDpoTDJvGutb
c2VUUq6ZiPWSUANUjQI7jwVxh0h/OqhH8M9nKXYnWYHe5pBtezNrdqdV8uexRe77nJWOyxuuLIto
06cVX2TmNeJhR078UGvotmF2prjwhnuMnPyHP6DXBXQslJZUEGERjWyeM5Gp3Wk7W2jp66WecGch
fWpDB7pPs/mBuseOVCPCgOtW/rRbXNlgm6jRGYfW84fvW8J0WSuv0zYhh8YMQklqDL4ZGbxRWS/8
vLTrl6U5GEBu+v8LbxS+X2qwix4oi7oiFmpgAAZQw9Qz1aacOk1RFoIf2Wd4xTltITTz6BzFVqGN
L0k9+7Skx/ayHrYIXewdD9z7hVa/14dKdcd9GjsCxSXRjJ9BV3MofLWBm0rDGZ5Xi8Oy3LfSbG1R
0MbnuCP8qHLn/j7W4uVVDUNoCVN66V1OOZWPEvEIeZWWpcHlwJoFekKZF/cMUq0a+LWdB/3rMAk+
pvTMrqgNT+43FVf9VeYBfaA7F6oVCW3ZRVQGE6wXnaOoEHg4TYDybKxpKYiQUqMF7UwSsDdD619E
9xkDKGWLjYFzRXXUOqPi/FggDMTdLi9gmGS+2c8LLsn7Ykjkzp1xoSv8Kw8ivm1jKarScoR58ryu
FOB9iF8pDbB0+3u3W89zjyLFg82JMf6Sl/WL+GByiY5LIDOIP0Y0jE8x2Y5pWVkBk0gJe02fXtGh
kEUj0L++8p47/2r6KVBsTaDW2Xx6thd9oy7dIpGZcBsNeDWW0xdQtzjues1wk2g9L8gfh+e7wh66
paWQjtwfKjO2SbzQjmvmxX0zAvJEQX8WNmZ5vtB2nb4Z6n48b5yBtlsBsLc4tlOh0BJs0G8WLpnh
8Q81tRABj5ZoYjbCGc38xUcQPMY39gF1XBtnGECy+lrWlEnrxZJrWlwB/dK5Np+aQ8wN8Ma1s1It
D7aHXz++T7kzLsT3uBYLT+Z36wQ0FrsnSVKAzI3/0qhMecHrMxp8S+n4lJlR1gNLufB/Z9nwNh13
/NbNpJLorEzWMk6j2tRh1itUulh/AeL/hCJlcqa3AZ+Zbkkp8ovw5BmGPQ+2wZwADNBYluI01kOF
Zb4ocpca7n0SwrapFm8NXOvmgooktomw3EbjZjbAUaTnNqqp8A6t2LNYfNShjmTfLSEUkW7brWlD
/qP/sXPPK+m0B6T/UmJLj6EwsapZr24yRYW6mzf7wtL9JQ93yLo0A6osOtBhp4ardSyzCgv6xYTL
qI4nYOzRsiJGkghPpXeuMJFuatH56zDUMQCckqmdF9P9c/3ujxrMvaJj036kHVos8/86aF0P+hHj
z8byWcX4azyHlWVA+QkFs1sxMQLxX5UJzA43FXfuwtAC/FzuuocnSUcKfp/nQBdq7tTcoHN6IqJs
qucoswwnqd6iDcQKqD79tA65vEBSGQp+Blg9t+djDl8AtBC8IJpy2c3hIleG8vMbmDvsJyXQcr4C
Xf74yIbTZremp67/iJ91KOJgfpYy4wQf8vWjrWZYP5rjH1DxA+guBZ6wt7I0+j5ZD822gOBZ6w7C
1HUId20aBDU0Pkm7Nqz05gYI2Gps8+vGsfbcuGFj1yP3BmHw/rGAg65c0QSVTSekmMPSD+FlD8j9
JQFG40w/5coftPYHMTIzOXqDZZ249vKn9JlRbFrzd18mCEMisQP7SBjGJ9syZ6GJyzimEvM8h7WN
8/cWTDRmLqqNmj/w7aoG/Ng+/403osYev2MDkoWZ7QvyQlRE5aUGIm1XHE13zTlZCTs8/nBV9Zth
YidnrSr1Nl1ZzsZTtJNptlOEjSk/pQtEkFdYlxQHsbGEOT6HW8/1DrfQ59uNgi3UKRG8SawWN0cS
6N0HY2kH8hCBKQFJ35bNQQHCHXrQFWtMrYIX5z4n1s0MheeRoMaN/I5+bg38OKVefRgdnmXTTlib
giYChV6jNJuIlbEIrFZY75k/uff8pSNdqGzvpdZsBcU04zElgGN3kzoXYmmgiZVqZv8yZ+NyK8HA
mPTtmvA4NzefxRnRlzVavWgK5Zgb+5btWqJ6aYxrx+NSUsLTjOhuN38BApiNsYtfPfD8DLU5dY4E
lrvawn05roSi+dTUJfiZ4CTftd2w7fvw9gJkO3X3nsIIQB3+e+6rPmhNtlmBnQS1SBflOWLxRlzw
kq01Ft6wZwHRwWbLgRKksDRLynXunvPEsA0yPZvJr2hBm0HLrxvA6D9hiV0KS9iqfkgmqdWjFHct
oVARMbKuht7B3cPcruKK+hRquyUmP1D5P+fJ/GuEQMYz7xvOviYLEI2lgcv0BZtm6cu3SA3ba/e+
AO3aKRJxsXs8h+0uiRONep7IBFAOAnXfKmwVCAZcXZcwlE3HVTyK8E20R9caSy9aGQZcrRoik44z
8z/hqD7nJOgF9XaVayTH+6HWviY9flMsSb7LI3WsHmJcJ45IKaid53HDtulKHHgk3R6xw6UkhV3P
FqLKT4Lfhs2CWlIqrd8P3sgNZRpZs6nIUUk6zcc3I/NEV8Mpi4B3TN8yQ55+cMl1RwSR/CikVPWG
OIrZyBMjNTe4esQr41ay6Iq/crqPilGE7PWQBqceZ4NOWpLRJlqZOJbFS8vFk6TEcojGAZWqPNsr
KQQuQtfWW2GPWQIEaavhqhuUOBJt5IboKughIjWZNYaWjPV+0XWCHF/u52LEKEWz62re5gfYPWuM
V6ICdhIZylQw8MVkJ0A3GDSgLE6TIAUSOpy0nSwDzy5cVPfpKAWP8+FuMz6qlCwtSXzJU0d2h7x3
dSVpkWOKfefnXi7UBLqfnRVpswA+SFhmFyD68RoSXcqbOHhKbxnWzY29v/gcnREiKrqyaEzPYka5
F2+9ueOlc6f9mP5KFHPaP2HuDlbOfDlGzrNKom4zF2v5TtBV91I+OWwhocVy2xwPhLm7srkMEcdW
bL3OQiR2SeUNLWMOfQpNP+Kfl+EO+aKuT5gzW0tuQ8aFchpOjt6e1N/rJCs+FBTemhPAn/Vk+fyb
reg/gpXkhfFeZUECR1uhd4pQqlufFyRZ22TrfiFtjEOmULy3Ey9CXC+RW38eBcEo055+wl43VFiv
aajbeTjjbnm0xbJUbUgcFGctN9YRAjr7q6LgKrXuJ7uydJrxsluw4hQWYoqldjfbi4IqhNfCxrx7
gg++mma1lBOTx4LuEuBHhRdVjAFZvbkxMyhwVBTOIxqi2Ge19XuYbstY9XXkf/mF7nF556wlvDpF
0q4GixkIKDwgyI6nVhvDM7/YBBFgtM6pV+FfonKWxOCPtMI8HYctAcSe7CXXmQoHiMqMfNFNxe0/
P8pKhRP0i2zAJIZpXZKCaJeC2kn0OSkYV9xe8wlWl2jql2ABCulnJIMjXQ+YpETJ4KXh0HfiCnQK
QGBzvEX+Ulk8TP9QzlgC7bqNKlzHK3Z4rwkDb6mbkN5urNVJgTQKWsmH5AeKFSU0qrARkNG+GPdv
+gP5bwPppAlwLheiHXhDUY2kCtH3Jvn1+iV9ixh5+ySpTM1rA2aiKbeYEfAa+t10fuvu1fE7YnNj
r5/qiCiNgxVYIWM0yG5S+/jSoa/8fljUIX5dARVR3IfuiCayURxIRgtEhEYTu+MM0oYxLEhXdXIx
RlrZ8nAt44ftVkQsK9uAze2Eai2uuXeJ56dQXvWa3zJKxnxuBi+nwFxGV7b+VWvgjftJqeK/uCAo
makwgj+AcuF19vnF6d7h+dXu6duKK8SalXcGy2u2CX2c4CAv91RWi09TiHQPg6F5J9OxunXRpf8h
llpsPjAgBhQwK2AIZ4CgsdnL3UEjD0Tpr8FfJRUjv0YNedJb9V48BOwfVbkSF3I6Nhx8KP76zJjT
WAPl7JSPK1VrluwG8ttCh4h10y8737SUSotKjrvidMrteTo3TUzlyLyOiGqm+V/sdoBHrLKFBcfK
klwwKRwC4tD9/PZce0TPHqjyKtIhDNaOx974a5FjqYsd2lH6DuygtNDhqXLKXI3eZV1xXWe4csYU
umxcwnn4TofExFtC3AUrxbDPSoB2RACkrZYd61NMsVCbUEVrsEfPcpsEj70v4tUzfIVQTN6HI0J/
1THcwJ6vp3ig6u4TkRniI2OJx14wK+s6EYGYY/P6MT96FZDA0Yf6z63taFZtzWz5noFkiOOq31R2
f1mu6tsUKqrjttdudYdszyitK9lfy5mAtP8kIoL1ZoG53B1pGOg7qYXLBIAxSzZDd8uE2y6dbT0N
0I1U8efCD/Pi1hAkQidiTXsreCh+VRIXJ3Gw89DSgvNcFkpSyFy+6rTQg1YsEaG/eahHGiI0J7nR
NRIjxZjp17Z1p14xTWYIvQ0LcL3H6ZH5FgEhxdzJW/3+5FwISWe7MAOK+zYooj6CkDOKFrsCx3jX
GOHMWdkcICKUtpRuMb1a4gG71/9ng0G2u5234Ik1DQg4mCEZwQDiq/aDgjwAVji901APG56TMGtH
aQfL5rtjrEVhceK7GL+4VzdZRMidC505wyzd8Cpy08XZAS37uZ/jRZDpnD8H+mtlB3D2etazTkW2
irMpRnVADH5ncZLpZ075NnExkNBhz9rAQfzxreWP0uGB9JS3YgJLwEdw+2+f39TkWjtd8O4jpaSk
Cj8mepUrPYR+90F/Yi9Sbw1LOzXiRlOQ9IUH7oHwXOOXvkps2HLg/T2Z83oq3Xs9PDHpj5qXgq8K
cv6oA9n+qmpxb64txCBcAAJfF7HjBKRhGhRa/s9P74P8ulXQs3srU8jh9NbjCjZrLYJlrP4bNG4i
j0OSOpYd5fxNgLbxN/+oj9Rdd7az34F0ncZMCduYRdOU/96q2F0huUPto13kPUWg+4z9F2H0Alsa
9RwFOaBh3MOZeLa5HtXIHlMPCJrIP9XF0e34TsdCgUtnEWygtpxX2EPujyGvExVWDOb/Hqz4CHUg
p3udSF4C7EPyKES4PV61ihkvAcV53Ujx1iBKUuWJpakfhSD+ZeoCmydCPrcg35j885gV9j9I9DkW
rXNBUq7yhP75vBdu8VPJ3n8XM94VsWTzFSv+x+lIYs2EvbAYmXHgP7t43u50VuortMNt2a56Oe+n
CWUs5YYQFmksQLxjEpBntlqyDRB0JKUIsKZFZ2zOud10V2y0zdljgBYhBMaoJ+5teFfDldDuP6bJ
JA64SjWrRCkLydKcz2sIYrtslrSz6ME4530Q8KYf7RWPnlqFfVipDrXOpNifZtyNUfPzvFwgtufW
6sfTH3YLqVO2SADb+IPJ76f1UiGoMyy7NzSCJS+qo16yph1RDa1xgQp7LhQr9X9YXKKmxbWVrOiI
6iW91lRZUQtIhL9CtduMbXOLYfa+lxzNoXBPX4jAYcGn1E734s4zuIKllC5vcdkG070SSpsRmGii
i+DiPj/LBA73G3V12M80qXEDdvBgJvQDmWiDo1UnD/6YMCPSdYarpjhbOLKgIdkQWYf7d46KIcHx
AcPVEazlCZ1eeBYlJRSz8komjzb7tDZudm35hjtP3sWOM1GPRrBGYNgvaB6PgSfQ4XhrEGkW48QF
hNvgCQDWQv9Fjsip3IGzsGNv/fRmyhkCWA0XkyCAcBwVgg4IYN0+ZnG9SHhXHEMM9TvryChKEqdB
BAUs26e9/7uD1b29j7KY2bZz2H2Rle2Ks3REUxUPMUCsiFfw/tllHGNpC7NqD+MOHkUYYci1sUX3
UsIQ8UgmtXIl//nzg98oM8k1S9cyvkSAPLHi1EegEI9hB45qAsqe1nIHyDMfALIowc8/36Z1LIkM
sQZhg1Ylm69SXuby72vJibn4iTx0WcUIzLTBSpbY1Y/geQA1se/Cnexl7yyVWRC/+yDdwFud6k+M
3AFMOL27s9o6WE3IcoFjhr5ZzJ1ySlB9lMXK5iY9FAdQU1Bw1/oueDYod6kB4a6Rbz/7aZrnSNxD
pkh/GNjmdiE1Quvf9IST1CqV4rSO71lMLHOEMiv930XHRUKQpPhXM3VTTPl1PMLcZgxfKj+jFfoI
yRQCvlL5c0VD5/piNmS2jjGxyBfLXyW05RxLyZ2H2x76vMtKduP7T88dkJNS+zYq2Kxjcmad2q99
lh6slE2ZmtbRRN3jtrHgYPZhkUzz2S+HIRXBOYSc1VTUUMg1B/OtGETnTv+0qmcgnp8Zr61CYoDO
mwiIOQISKJks5qj8sjUmra5iNm33eu4i6q6ryOGYZcqK3geupf0KCj9ZguyfYKvKK3328c6p1w0I
G4uWLsHUwcfAvtss7sg6DbkjeoXnzH+/64Dpe3hCPFIEcemCVIw6Kl6X+5wVKNlFyM8G3VzWuWTo
9lfR1Fk8zRXPM4g7RhWjAOG2F3DRTNkrfe4QRHB0wtE8zgVAtVj0YeXVhQxg+r+Nhk+3cMi1LCch
7SYx2npo0iDIKCdlVMVAvCmbBB2/V8BCjax7IimDuo4rEmI40DZv44ZdAPrQAFjb1isonnU6fGx/
bCQpCup5z6F6dG3Q08OFTzPBjSF63K13En8szgBj4kG90IniMd0AL9FIhfJ7j+QMluXo+bo7fq2i
lReAbXKDJwq2Frw/mIKR7qE2iEJvVkCUAS+6qFpJSYLKxG6Cm7RtaPrMUz38OL5lAkMce3LKqmU7
grPNKSQepSGnRuyeZCLV9LaRZGdrO6fNNCNrtuy3cufgBvIFf660meCcrDyD4wY1SHO3NHs6U1kF
SaD30pxJF5mHQkx8FwZI/vceVFEdguDhpUHU2uY19uLriV9TpasWrg0Lt7O3StHbYa8vP2dJWLEw
zLZalNIswBhzVUIRs87dhM2wPHEQ0EluGGuMiPuToOGnstgslr5vySUUoc4UdLe1t8F4m8nkRLGc
opOWDS9/cY9qAmW5x5/23epy+qKaJLKkBYpHrbcYTLDGq2JDgrXHi2Y46C0IeDTriXuCGiuRefIW
itXbrSFtIDK/bvaJkh6C/L2gKQX/poW3SBayRvJwKFD/joIGjwsiAFMp6gXTn77EDc7lVK6BhP2q
8PosDOkRPJGuEE1ZwMFGTbehST0v6QQFSVxQYHIV7SIvs+jbw6NTfk8YT8kT/pZ08qoCs+sUNldi
CCdV/20AT8rdQv4xQPTdWS1mLDrP5Z5MItS3psv+IiwK2fGQzoBh7r0B5DtJO7m3f7I4kUVLGdtV
hfd8IU1WW4r6UEm0cJLvkVQCe1a+Rc4mawynOaqZxD10al1OiVoAphUvsBgRadTvEiyu3X1jXf1V
w5wXJ3kU2N+3dwYGwzNM6kv3FecrCD1bMoUqW2aK+eQpPCHtFBnVSp8cDiY5hfabvWrrSFJdqnCP
TzP11wr52XA5odVDZ67Vko0ymbEGyzXUwmu7yqt26/kjgTpLApCIjvChIaS0B7H++g1pJU5S0RbA
g2o7xvmi1L099JH7gQisJpJ0sJ2C9clBQOWm62+tL03aEgpZh2/cGh4mc8s5zbemmK79e9Q84b3q
/l/1sfwnqd571OKZfFmEBFaRo2yBnz8L/TXUaLFMDwUwDlL0rhmQlUnRwe8JAF8NvAyG8TciFHfV
G/Ji3Vbmby19O0ScTs+7SpABZbXcp2CYkzhZ8HMaay4c7Hw7P74CRFsL8IK7H0y/La+GYNCEOj5n
YDF7fzsXob+d1/eAuFmj8WImel+vOvZ3D7bQp3S14u9JARkN+zheyVHxyWON6RGYkgLLFGQyzIx3
RgyB+5qqe6X/ZVQh7euXasmrLrNCj10Zm3WFgR85zq8bSbnNjxCAvdTVZTHgPaTX2+6ANRIZIm0i
kZXWGelCfnglTkMx8T70VlOeejGVIhl4PkuCGrBNb50CZTOI+iulC8nXc0zEEUcOVXaLiRzY2gZj
uISll44lvziXgdjkByAC0IsLNmLMnQwNSlPeQOppvCWGz9PxCVzWKq8k1/uPd0N0Gjsa0NqNdJsB
ACGm8x3Iw1ryzdalvLJowTGthPBaiXsrjuNY83WnM2Vd7G//n1UlyKXjE3WPDCrqLYFmf4OhuCs5
ZU85QaLTF2fO0/6DR8mpHZ8w9ErUFEXFpyXbWloIkUPyOBrscRWhP3kw5piGSL/OkRYBuzNkEanv
vDtKSUBeahWCZ0H+5sKIi9AEVfTh4yEFFAdk7Rzl1b/6sY9InTSLLRB4uVXOWPpOhUwCYM2LlKog
o2YDa3TrZX+aZFVnohYS4HCJmWy75mI/4GbSjeGcVA4KxNi+2lfQMeO9eyrgQe5ka1YJilvo1F8o
Ci4smzuZ7YMQmRvQ/RZ9wWDn366UJIPEGJs8CHoexIiwZFOycEk1R9ClNVzvxgl6sUWPVJNfRNPH
8/PalOWRAt99ePtTzXxmKEWz6CdcB7X2ZJIvGg/nXaHKEkopvCNWKJv/GWAWSVYMcEnYtL/45Rna
EBRb+CrD7jqxf5VM7nl5wCrcRuM1x5BLqHrTCvgBBgcG4QpGsgWegmcaUsazARQnVAlMg6+t7lh2
0JHpqM2/mSe2n5T6iZWAaiyDxKnqfoEpbln0+MxR799LvsRQ2tA5XpJ23TqDLCzsgkRzJUCAMKqV
gyusNZe9vtSA+c+H25tPi7xxZHGSBUlmF88A2gZFr5ZtBANcIzb9QbzJGTn890MIGAMaFeOIDWum
vtz1j7yBIMTKrnSuQXTUV+DckRPXLzGjwpvE5QkVCc2h2gzl6saDHYbOu3KrS/uHpcRETIMpguCf
rd5faSROQ8JliXckWAEf9hBJkYi+eoV77i8tKjYZpM+q2y2Mw3Ypmk4mGWEDaOWoe16Xoc3AZOo9
YG9ZmbsZEtFCrikwlO+FDVdc0zWUpfyl8kC9XBWuHIiQR5IyqKY3+LA7+Np61eRE340UFfJ+u//J
D81zFzLZzUlL/FCiVx67ICVi2jagykh3bT5QfpTzmOCEyzB2MlNgYS76tG+VSd6s5APAUJwJ+al9
jPblC7gZ7VI8XZmtXSqXFHujX+BF6D4zc62CP5k8QFlHoaSNgsVCrbp8sQgF0lx3+qiF3p+Lfnt7
gps9mbmnK/cE69yn6BGjy141yxi1XmUZMvH1VfKEsScG9+/On29WuxB/D71vvwKUP/NbPgF4V+5E
7yrIyIbdsPuaAA1y7HPMO3DDBeaxsMu+u6NvIGQgbUrY2ygKDjXL1HqQENGu/Z5tHRY+DZ2Lg15p
3w73vsYe5NVd9MQoQ+0YVg9adyBdL4w2yzbGByQLVloJ9Xi1KPTU833/YOmts4aKSwxq4JzHmJNW
wr+okFDgE5BChZgQPCkC0pbZj2xwv8yb2XV1AK0CBlaqg/H5lYGLrKV3bOJQt8fmIZil4IzG3VgF
AUsxaVSOl7Ju2CSus4w6X/r9AawfGAQcbiisIgatcr/4krO6UYluw8KTFvbUCMzYvA2HAdMTjPEL
qBYNF6Rn+78vJmLOdisug5eVeVo7coW7TZctyzIVuLtmeZtIb85Aud9YM5CL+J0Mlq2mQ6hjFYdC
gQn+/okQpUyWnKCUVhTyDkglX9PxIaMDVUtutOWheXTbhdNUCAW6NxbV5GE+izyYKRLyOBssybBY
Lm1/wOxAjra8WpB5lXj/XvzJcddpjBiJQYPQCIxIWULdRDJ4Wplbo6Y19qujzEZ+sJwUPeKR3fSQ
s99reOL87+4WviHiofOeI2Z/gfUt9T15VI1XLqWJ0xf22BSLFw66t/uNbbuxHSIzlvUzY640HGfc
ky/DPeG/pMbUS3vhskF6GboQFcZpyqbN0G+uaQx2hdVvVcdWoMJkcmeB+K1xA1B13EErC+0moNlH
UWATMHoG0lj9rN2kXV/zlCGqgL3UR6G41dFR6C/8ifwcxXCCXM7JenoO4l/2tl+FwC4v+Z/xd/yM
G42Tb3kiW9qUwV/QQ5jRLxbGinuWDBX0FzgVS8DUOIATchCc4uxHCP0RGIqEHu8EDVa2iWNjVaXY
rbIsfmUK976BgnDMzjd53kYv2uMwZ04cf7oL2uhqSYIRBC9/jgc/3h5q0BqMg3W/ovYqWR8SiP7t
znxLqXmtylYcnsJvPHGoAhZpklajg8dJ9IeEdoebCj3p43xH6rqpFwQb42dCKppCjcIA702cNQ1x
xcL/y/cZC5vuo0LIneKHQoNpfLCPFzuRwE0rloJ6EbiKYfNPL/esbvCtb94kw0ZkVZtZlblXkD8V
AaMW+AotHUg9k/fyQsZs1g/GiFQmUHv9WtGcszPT8fK7RRVplKSWdF/EVmaIQAnToHXPF9mGdIn8
qU6edJPv6W52CaQFVNzbyubvobIxWNOmWaG0tyTxFE1GW8r8sfp6mK3xzDkX7VVsDxe8D5zRRbzS
KAku0qsb1Qt0RqdoEoicMiQp59q+iGYfkBypUpwU97CZQaq3MIPCmxJlCNvsx7/ZY5P+7brcfGpt
ov0NBj4j2MF/vHZ06FvDT+m+ZfxpR665PdtcLKOtEiIHoM69XuU0IFDQVCho2FjOIa9zggOpGSBe
bnI1tLguMbWAhqL3iyOjsCOi8HM/nlah5XBjvXz7owL31Iwkn7ewXoKgY6eD1Kqy8NW208ZXB/o0
4LbBq8US5yv9I9yMMehfHqtGHbw6tjWFGIwA/wUjVN4dGRIIUGIyvljtmR9dCEBd2438clnEaKs0
9EbNIuahf83/4SZsOeLmYf/bX8LQIINaJCq/NdmLZIy7m/eTOyPMKIrb51j9UE4gHdeiVNHXFCxq
g+eCizU4/Bz/ZfnNIcpemH9BqDbQLSZWenPJBYVPrYi8kH9vhWJ2KxlGTxtDChcb61Hr24dz9aHq
riP4aSNgfy/7dVFkyw3xOjWp4vAI4JZwRnVCrQMStrzrOQR2tJEXfcEEQ8d9pf+oCjaakYs3OXtb
/9vISad+ORFfHIgVudbASbiKbbM1/O5+H+CyTrbA29RdPUh7PabXKP+/YY2Gv4ZTOSks7+3Sodk8
DZ674/a30SkCOrMJOLC0aLqFjbOHolUbDeCm50MzYkcw8iAzVYDlOcvJo3bSzK2zK8KJyb+1VMHo
p74baT8UcFxohv0vyREIxxs3sE8P8a8JiwNR3k12imR/1opXMk4L09xy3r7ZiDmMAN+L2Vcn6Cd6
vXc/aBy7QNkOqkPF9y+qYoIWfj0D4c9Wb+0hj2VD8ePH3HEhp7qD+77hpZ5sbCgLP0OzUoOF9BDT
HjJVJF22D8HyJehE+W9et8qA56GZkTy6eTvpnrciunKuu2AXFSvuwzXQiebO4ANCmGd9oc4kvav6
xpskhotKviFqVgcVpdrcKJLz52U2e9IuNsQug+xa31kr+X7wbwiMO8W18T4XqmHHacNZzSC0mNIX
MyEJtHnxh74BHZ7zIcK75PnP2pAks8gPPNh5jRWxg1Y5mJyDmobtanzQjMoHylprJkJrHqRek56B
2EHFzJTBAcGnMYiYBzdu3+IeN8Axb0kVDPRyoX1C4ieCblIoHg38VrvsmueyjbpGN7KJP84X7XsX
1sI9pOJaPZ/g6IfCmnirXeTVvX7OJ/Dx/0UQsNmaJk9CDktckWEQFNXWHfnezvScSifzSJDoUNG/
ZW4cyLlT4BHWIYKNevKwmhcryPnVxbrRdUOAK9uLiBP2/7LHtRFC8nHFgIXR0ahW7OdoeVYytxgx
xYCLv7BxfPLAc6KGqO3tsKk/alf3y0H5M9Rwj3t4EvdIhbd7Ik86+njVqvCgKIVgXrFI9HNFFDIa
Fe8QydgC0sQNDlT5nqvZEdOzjUfs9IPh5Ev2QKEubyygUTiQWpY+qYMolSzynN7iZEyRl5U1w1Os
pRAOVj2WTsPODzj+7Ce/PnI3E5ZNzI1N2cNDlXi9imPP38zcpj2Djd1SIhlMvfrgpC6OMFojg2Q2
9vR/yPjfW+Qs73j8IciqIiOXAaeKTMuD+wuFPOVP0gVWHSEB3gdAmCBj7ydJAHgFi9m33kSDuyZb
zMeL6vh+hUg4MnGVYGe9kqrTty5TxyCuCCPnSpD+n9uyvv5eibh9XKWpMSiucrxLaF3/ThlWV4OZ
BUfTn/adZWCDNUil5tws3+U6w/daFdCpIV+VztFfMI2Bii08/tJ5N9AhElie5Eo+x2R6SQJ31Kfm
nN604luCRAYKxlg+DXwxduScPfVqalkstv6Y0RvV4478uT8HFv8YMQ9oryVSwkCwe0YKSe51eQA5
u+WeELlXzzFgys568QEN/peB5eil78aL/4ZHk5l07WCKmvG934B6a1S7eWkmQ7DPIYpKsIMhvlGy
3GVNxMiADIceaV95Or2d3ZShZUM3BapKN7mQHP2XtLj3sLM5n6qorMTV8msBreAzT+7jcVFhHJHF
VHPs15izrJtRaycc7uaLrP+57NDWEq/WGOT2B2qS9x6ZTHFvbMZcpDyOD78YEiBxBxZMtMNmMr15
Rk/HVEQk3AF8yZJap8UUs+gNPY900qlgA4yKMc1HwLhWd1fVASbeQemQA7ltCLIFsLoIGrrQSWR3
4BSRk+qpilhd6ESIfkTYGqWmqsU1/Vze/7IM2HyLS33hcPaHhvgzxicVjKLaAYl9sUHCEhAhoSZA
to2reo/FsxOxbgTEKQR/S5hR7gn91Ir4fY6NUjDV44nJbWqbQoqPiP3Sh7cpMOMQu2TjbAD0kPoI
1JSydImpLgFeSHiXM3GYwC7c3HItyqwgpOBLjneGGfZXm+0EOkziRGjGO4c1SNROpnertx4NubTy
v3eLDthufgF5URAtncoQMD6jO8t+PD5PxWrQJZDdSgu4DXk8VpBlSf8ZdlePVciHLGd5veUg2VnK
xn4xvLwnkJWVms6n6aQLJoYj8+IRzORAXWj7pD4fYE+byynfFmveHGudq3HAyZovhHcFl+lgQKI0
lWRW+DNxSEhnkQ3wiWHkGzAsnG7/1sxWHcTq5KVq0LONGnYtxJnbGKSBmr+gZ8JRBA88VZnJUDzS
dZmf/SMhkhPFD4oSKFDyyMgNw9do9x2VtGJZYKNfpLLn2pqzvsrOvLVI+i0oOETXxqXpyBOuqCO/
r432fGPL3MtZK/ZW9YU3snhJltIIMHsCvjZP2IicJFAXRH876CPxUgTaA1PVm6RzhJeCJzxQqdZc
47Xw9ptFIZsxfC1GbCOHuh6HJUQYnKbzIUVH4TeDVO81K5WQQaDNLOqb4cIygKaNB/U2sBa3Oul+
c0UPUgwfLJsJpIHOIltzF8kUZ0WtuCmiVpXkiSGiQAYHxZDOC+uXtb2D0ZQoJLTpPJHet1lUbMq/
tsskZIphDkb3h+rT7RNcz/GFzwmnfNoNuQc1c2fGWbjzVfz37IWyIb68u5ivlGHdti0fCwkaDuWb
IpzMmXoPwmywrLHJeGGYB0XT97WzcBZNKa1rP6VNp13VhtGWSkjPz86pJbcSXXEBMlBWxfAOb9Bm
zNL3ocss4KVYjznJqAEqjaHR9/A18KiT92Cn2nJEoRuqTbkurG6S7alQ3SEkSTxPH4QLyhK5G2on
6V/40HVyp/iXZGINMULWkWd6kOTgja3oZ2QY4+wqnhxEOD6ltjaJFbcqll9xyzHd4ctQrZZf6bFN
KVzPl0aSG/mT3fdYL7Vvjbe+wYAExu6lZHXKywvO+1VIY+UDHdYjJfulASMfKC72yXmX+6kdBpgL
euc/3kBdlZ3O7wI6zmLxCg2vXPeuou0lUewvCAL5bF1XtfFzAWz4I0B24Z4tJok+dlbhJqQFVOnF
jrQ6OBYqdY8m1G3mko81gnullJMa4DX/FeBC0XPcj2LA/G+GWZWHTABW+mss2kfGZZm8w3O9Njts
YLQf19ueI+BQm47zOy5WL+VegczEgw24LvZXJ8yuQ4Cn42uQl3KZBExp7XzosfgcayFdPirhwJnp
vDMkYR9v8exoWOY7rPwkhczNN+AEF34KUeDafJsc8FaLCEvSw03VgHCouJTKebRdffTFZ/NLvhkB
UfmfdX3K4Vyf+79tDeopysyzXBlRobtDRhH3lMqgJUqhvAh75483mDcfZsfci10JR395eYBYYfvu
PfIk1OVx3Q58fkTncrNbv+L25HNzMy02MVb+Hw5Wqj5QSjudyEfgDyr+OvazA8z51i920L+3fX6T
1IQUTj/VvDuZE3FG1AKnR1uoiN+EjM9ce1n+pigI3yKOsjqPtPh5V1mG2xkM3ga0Mp9A1CCz8zDG
JIFjYguMvYJv/87l2voArvCEBlcZ1sDGRwpHYl2k9lzPM+nMzRbTfTBuQ1uYrHBJTEThMqAxCUna
ZO0SiNpZwxQBHP5D4YkrX2HKvk2j+37BYzOqR6QFZLUFuBurwziY00rra5tiKPrSJhODa4k0V1el
OvfC+dghUEc3e1yvfRM4l8k8m1yNmFrPZ+eTTV2x3KH9weARZOBGvVxaXG7+WoQiqt7qZ19G7Dy/
9UysWkUy37pvVTLYFScumtwhwhsGo+dm0GvVeu8/3H7PZneL+Uyvg6HDsqOjqqREpZjpzgLpkBwY
xRLIEBwwsxV6Cj15kQdsoYwW9J3h+nYYaP2OqkufCp/zCI+pmOeJYstYD5b+6/77ZnOu/lYpXWJ0
xbeD5t7lF7487O3deZgwtXdkO9t8OkzTM3PEfrD4yqMc8GAQiZuScQdyTuEgQKehiJzJA8fOUUfy
YljJQq6dWJugdpmye7pxvv39DrtfB87eChGBEKv4azSHJ5+LdC0Qsaiz+JnUZKdJDmfBXghuEDXN
P/xH4MNpV2mJQO0cns/WGHnAG2eMMyXNqJCPzt7fcHrYDxoW4P7nFDejUeKxpONQ3usCNzWoXJyU
BgCvqLPKgjqwyTjdqoGXDC3aZxV5qjAo/y2uzyKrqC3G0siiqkkpEt7jzrHdcFqnl5Qa1rXNLcrW
OQETJsFUBv6Nbl+pfg5w1rThF65FXxstA3WDwkdz8o2vQRVF56AInwDAN9sKxcmwlOueOryk0jXv
ut3KT8P+diuGZOIas2xrKH43sWytIWwmrUKuWOsXZ01EfpJseuaK3RTOsqsPKWjWz4mkJkLpeAvw
NZtnxt4RanFywKZ7o7du5u5smHvRjmOD16KDwR7IVejYiEFZCbdK3iMsvO/luXGcrCczfXY9amwF
bmajexIKeIxuplDj0skZVJYozKNvHK6XI7XFGCIcd+R6zLqBvEMO3+J5mZVhGKmHnOxZ1stxNS3h
Z3XPGNzzFZHZa27TEYmSz3h64KhENGxKUjTwAqsIHEobBl30jC7wZJEBqHmsqkY5MgDWZVFHKXhL
UUFjhd08y7QWabqrDGT7CDQn4bgf+8f/QB81/3lfe3ff6bvsiY0aMprhpM+l8y4GiSKUOCsgtNhS
sHiCo1b0myVF0dsnsvDZHyhtLg57OpXUveP5gmxUFEgHjS986LHEuaQsQeS7kQ4abBXAua9pZNNb
ue1NijhMbiRnVyrCJXMorkP+Ajl4pU4UzO8yX95cokIJ+qM87ARdlG6+Ym34eHM2Z6JZsiVC/O2k
1fHQbqRklwJ3OVVz+VONaN2ihi7/aPnek5pdLXbYPgtrRuCSSz8Xzch4NX6yO+f5w9Z/XyEc2bU2
gW1qEW6GqEuYAI7PlRgygvfLhcnnVIep/5QM8rsqniyNJb4xje0YsZLTDrYIbR0xs+/BcO+hHoHQ
5D56P7NDtR9GwxCaT4s/UXd63spV4C4FCLynbAIQBRRAHzDoGxEYejxaSR3onsA2BO31bY6CiDjA
LCaApUwp/gmj12aa/m5eiv+wVMHIeqkfuycApkRe40FtkTAdbdbHBnQmsJlJHU1gv8BSx4DI7pgg
1CNqUAz8vxsde9j3PqZJvU2WPpraMnbn3nL+cH6QhEB1INx8HUADIoLDNnfR2FG7wzjHAph0BLJu
gA3kk7sk5kKVms+ACuSewCdRgqJ8UC8PFgjwcmczhkWgBWZUkOlGEnHIZEUI2A6S/IPuHkeMtk0L
wTVih7PN5y1Je4ETCOxBH+E5E8O5kOfoSsosJzybV7DPVbBe9FwWvAgM/BmogU/3w3eUUircuiiw
YKfu89DwxqVCGOra09Bug4F6lf3M4k4BcLIaAya/Jh7Tdf01vZrIc+npjgRvx4yAEiIt4DlHx7Sd
qaWvrHJ9nVb6d/Ul6O34oIbkVMqIgzb+UgAurV5tP6bgOrsPUuy7mi1KBHW3wUBc9cuE4887R09K
xCwSJesiUqw3QitGM5CnEkPcZy8jQtzWwoGdUCbSofoJaiN19KeTW7kxLVYWbwUIyfY768awICmx
ExHbgBGHCHin4cvpB4iVHLC+4YqInlnXu4kT/PCNhRNrlKRpCdMd+Epvlfvp+fLpnxTq0Zkv3TqT
sO2Nc2q1CgI5quWp2LX5ZePj1mWDGwjHdO27q1bAGI8mC6GqK+kpRRgRBccC6ARF2vhJmnz83bJv
fIqlHj/GV8BeEhPFh+yZP6tQPZrU34Y9uJ0UBRZQhLcq+Y/FRLaJrNhHfZ8p4UjkNTquzOfFHENs
nmS+mpsfe82tJZPP6utK0ziiK6lAT1dPvc/uzlAuMLfW0LQSmKRmOvLgf1v0/VP7ySa9CQo2/qdC
9uU+Y1tSfhwaEK/pc1xWtE1aPiVDeBLaCurw9QLRYWf3J3jjy+QXb8QU9h5wEtJjT4YWqX8BBXod
d8cIxYM6NQURn9/IGxNmB0kIxzDrZP+H9WVh5i0wFBAjSZsT4YtHm1tQH7q1ahupNFRDJckYg8Fn
83KknJ9KzmptN/qkh3iXsU15k8PZaJkCBuwNNtFXLpBEJyovAAUEy3FXsicWbRef81QnrSfcJra4
PU5wE4A7ZxEIIhA7osYjkg9wA6GDoi0qB5Q2EJh+q4UGXRxh6JsWI4JvvF/A+93mav53LcraN386
W2iwoKY0OrPtpm4fcoSmiVQeW8Mr1rwXT3BFLv+bII7wLwt8aDoL9WCyfX9Q0viliv1gPbAca99+
GYfDFYCy4sZMSC3K7QVrk1ddvyOqVYjFFxPknDAeB/kmBDlWi+yD5hWh0gVz75dIY3Z2DIT9+C3p
DhOeWR0eIdeoiKxxPAZgL3hGrPkZgnWuYvQpVqgEY4lAhrwOmqz+xxkEpMtpjLUpy1TpPnd7WSnx
9aTfOWErv3UqGBbR9qHk6BMZyY8+pWNRm5W0Lvtn3erUmgW7E96eDqFKp6bkqAs/cK7SrbL+7cER
EnKqdSdtTMQvUJSDgD1Jvvd+t55l0YP4L7BkSiPtkM29PNmNcgBzG5b+XdbgAZVEmFvVTj5vW3Zm
6Z4NX4KsnbNJoQTCHH0Vt/CpYJhk/oi93/hOWecJzpOREKRSm6isfHlWNBctOA3LR8IgQmeiWkvK
RdzUMdndBbqjF/v4Ds8903uXSW8Q8lObPEbWzOFqqgyKDAzvQire1K8F0iBlWhFE1YwwxDw9Q33l
d72OiFaNtFf2KO67hjQcYoq7dMVpIbsoWSDZJq8+YItcJSPj+dZdiCP2DRAkMrQnE6h0KJpnvKXw
iJgHqFP+N6IKV4dQrYUmn97t5gBRED2vr2tXROZx+LZuTl98Uv7uXTDfi0hg67X5SHgamsFuS0vK
pK1edQ+wzqKIYe+6ATHHbNMZ6HoMwVIAJNexHOHF4xcR30daTQRJZyUv4PdwUmwLK19uJ5g0RyJv
wh94IEo8/PueXACEfNE3M6t2sni8MEWDJKN+rBnziXz0FmPZsGDXtFdlF+Ji2cf4qYxu4kGo5CHa
I+PGtukrF4gvTyF4+C5f6bP5X4x9zFg5WUuCu6TQ6bPh9kdbjtCFA7Bi3oCDurWBJS4c56YSCPFs
jYO/StUNwf0YGEZlCx5bWJoxIlZilzuo5SEtYSnmXhqPx5JhWhe3xKj5nZVBtg6gaus4KsLjEFc+
Vd787tXBfcR5zwVQ9EpeFRynBh2GWDCIlVFDYqQ8la6/eyhjtRQVKxTqTmF637GeQ3b5KUrao8VB
ZHf+YFsx4OG+hI2APWctNiR+KgOxJQiT2TWAnzo2YosQ8eg35R3Q+p0J0UJAGaNnmuYw97/f2qGv
dYGSI3entnbSYrAjbaAKFGTovPY6WwGTGa2AAgsSNCwdnnCLav0jA97bmazXF7IMM9xnLTb2CYBj
rBwTuIrcwki7E8djM/kzRBtjZ6U5pWxl6+UyOw3yoE0u3nmRKDJyA29ERpEQDSG3JQy3+BffvZIV
uiAhqRivrHnl21219KhvQoe40AHcFay8GLxJ9O+xlLyKHfmh/IT2xRoYY3Uunk3sRg1WTeDOVE3L
NNFM9+LY+43Myik8jRHG12Ot3UKYf/4tm2LqxKBcFyqjNB3oyRkEaYK70M7RI1bAh3kV/4HEiCwU
7fzh+9YUPSm7bk+5v2McbAoq4T6nFfSVFdz6vCvz6fOia29Bpcav7J3tosg4iGud8v+wr0pOiEOk
6rpiFlU+/A7nEtcAEkxaHVNrSE2TSTbupZSo7WgTuZnno+K7yDMNrwOBL1/xLgXxo8Yo/6lyeQwb
W3InrkwV2JKhDTDP4shH787x8ivIo9ZwHSYv3DVtYYKQopR90xzHeEOamMJ/7ThIky0iNadgLo8J
5khu8lpqgH++JbGKGGkAVBAxCwqrxQLTZK36UXDmDcCd/sN7jrZ/j8QIqE9cvCnqPqXEeXDQpNYx
b0zGNTQNw87UaaoHaQ8wGH73FXlUE3qoADDtnBIImogdEe9utoXCJM1Cr1v2JP62f4zACgBZ9C/B
2FrB3jzH2aotZUaEp9gRTQLznVKTqxYR/4aS+4sMt/OLdgpAt5bLscjn7bmh2sQwvC0mf9Xx0Fq3
wYPkIo2XpdgUDb9a3yEa9Orj09p5APauVil+yaWeV+JTVx7mIfsNJM6tuBy0MGW0gvlmFDblGi5V
MNAuoOnwLYGLY7cThKVaRIfmo7D2CNzSXxsDSm6m3QmXYpYRKwDLVnxJZRcXlAj/OspX8Ps2wf52
REPJ51ni+t9DjqFyapvrgFxOChUytMfqQHhnXjWlt8AReuujsRPlvpoWwqwYk91VULRgaG12Jm0B
4QeNx0OIa9C7Vk77q9zWe1T0BpDxzg7FnLEHHLH0XYr0kTjBzIY84MATXb8UyaDFnXBm/AWodeMz
LRwv1OzdTZabxW4LFF+NOLvBRAgFh0NJFqTquHPDIeEHVvjuPhcWH6U3JPOu1swAZo/9C57AZXXF
loMMxakEYJwVdkkVIiGIejLIni4cbtYUlatYXrUt4yZxrZUFHXE6GBiiaBTZpi/EMnCrGJ1+oJAU
6tMgdhBovpA0sPX5ZqalOlCpyGZA1jHoYzqu0wMor/yr9ANUKaMbVHkoVGz1+HUQNlmmkMOG+4D3
i3jUSdR0KNw+8Un0nA+YAjQhIR29BgAUXyWDF35mZB7U+/VDBmX2ZXJZ5NkGvbHrRtGJFwM8FrhW
P3o9SV3lSq7Rj63gLnemoP+QhXrReuEAZbvdQNTtQw6G3gXwU7fKjOhYnzw7VeT4xHdoApJ7V6j1
VyOxRyUPhbWEVRofEGd2ICY+Gb/WzbdviB9EyoXbqKHp5grK7g+b2jmRlKeJVnQJCNocR0UcYOZr
OYHEh/e3fb3ZkgsD5Va93/i85nhn3XxGNM+hVWLLnwQ36tKRIMXlmf6gxc9G837WpDxA2iNpYhwP
daeU+ppclNe+vNEWsHTSUAnp7oJJG3Swr/yJ27/ZtTqTOTRonJwP2J9zXJ8PDwiZLigxMxLNkSDH
Y+5uooVpITLqCVm+Nn5805szypr0n5JlYwOJfDhjT7q8xa7+Rh6dA3bWpFRaC5eHndvkYB0SMl/8
NjxtdAmn8qyi6pxgiVqKdWrYpALbggEvdGE60DESbOIcB6uUjvnWB0+DmJUFDxqPxjH+zocjN5pt
jPhSmbO5zxcoktuDwLYPoYs+qx0hIGEl6hoG0HMKs+cGZfJQdVtor8LXgPxtpqfmBvJV/H+Mfrr5
+pSHp0m0Hv5op1gVXiXIiVZ19qYdnlxgg5PuaXzpysnESYXZGj0wmEd8Yr2YCIHrJu+eKuwYCGDP
o0wVApjGEEDhbMdTG1+ah+IPt9ZWhWT69wXQHqUaMlS9zhm5DCF2OSjP/aztbbxqULwBxgqR+lgX
f8us3V6UojERJpdAaKd41yXnK38Z5Oo5tOPHWUq5Jo+OYZwW258AzxoB5HslJJjybJgIRMI5reIL
q3tX1tIsAjgZWP4XoZoAYb2RmXMGrZiS2xCRu0mqAXDGMNpvrHzOU/xZtoMOJ60hiqC8wlCZHCZP
VjaFJtLE1ezKPHC89JSlddXVU0zfgvNBXQLahRAzuW20pGHmP1qxwOdFPYjIU2RczzjGuAEkrBqF
EwgsQcttRAjhcWwgmFEESZp275dvGWA2mLqSYvMdNjsFOJYzIQxu7U+w8DTWF55LSpxQRimqBt+c
2UOFdY4AYXpRaAb/d+lxFlF3uAOctG6kKJ5JPyAVfI8ZQrE/oBMYQtZIT3UPcqErvNUfH0yza46H
XFcEyUJeTkE4TzvpXQuOt+HnitADJg23uL13N+KpZ0zDSxzKX3pVMKuJRqIlxbb2Oc3u1uvPxf/J
XpGoy+PHAxA9OhtD8WD0X2HBrU+1r8+A/yIIQgjo75/F73RXCPbBBd+YOiHYBLhrY4x0LOHhoRdb
xqrasYoHiNLhXDebSB7ERC045AlgPNP6Jd928Ztb8E1UwDZ9HuK4uoFlaznwFHBcopD0Vk12Fhxz
y3ku3z1AB72bptD4zYJVZZO8HDBnQrpniPxaHwV70aJJHsILyw6BpECXNc72V6PNUKta+fqTrssh
I47tlNuaJalDJcCTavDdQ2lNtyomARXjO8B492Fx/gRHvdiPU2Y5vMj5kjJRhcCkZCL/YLyx6J/l
DMoEYcSgkv8rYppbWgLaS3u8PbQOAMUak/Tixxsx3tiFt6n4K4OlTyGjv2fStFnhoBx9o96iRjqP
KcayGcRCfNUxRomP2OGmxaDOX9fMlIiias/VWhg7jwodUwFcw8RrLOTR2woC6+F3lcZ1F9ysK4ix
6r+YJY2PjK+c+8v5NrToeoC6v9rW2HiOORESLAbWzR+ZdzjGr3ymjwtlhHJFKMzdt2BLRlPOqWFV
Z1evTSm8zIR96x7WFlHjuijYxarFGflDJTnj51r+ajMcH8YQySlSGpzq7qEOyM7Bh8CrIwuE46ZF
wNDXcNek3NWZORq9GB/C/EYIHnoPXAtgUt3He7dlEaej9qrj2NexjctJ+6dLfHEe7V1PiExyiS1e
iZQYeTMYJrqA94rAqgQz3iDGk/+HjXg1oYtK7aAY7kyQbxCOHjXTueQb4ZXb2w0Ny0loPc/U3K2O
8zzAs2CrrQu0NocaP/LdI91xs/R4dsRLHNTbwrfs98GNf3vrK5ooFcM1aoXuGBZJkpXp/AQh7rV3
jCkpmmywjZxKROa7b3dgtxcWYxNiwEc9wp3CX+j33YdmLou/zFmDe981/P3tJgpD9Zz6Ql2A+2rj
wl1fV52qP3XjeWhhRctPtq3jaQZLKlNZpngbKOBDLPHqgPwF81wGEE4tzRXWBtcpHpHdgfcDwPGQ
W3ocK+NW4korpkwxkYuY5dmCyzLFLM2tEUrB1MFZzacbATQW38V5BSIj4eKdOJaReD5dZr9U/tew
QV8DcRh+tD2vPAkffZW65iEw9AhKv1lKnnXL6twdEzybrwG3cAVBu/3cNVGj7/dJRiLR8wkPr0+n
D3vELYhHxDYNb23Snfhsnk0+dZwD4UFc8uKG8gonQkfmwbbHbmutbkgzctN8rn4aoMv6J5E/1fSU
MukcRbaFnHxSPU+sbklR0yc7oBQcWWnFQ+2UNlV4vc8GEE2nb5nFkzcPLGt1ZOZI4UZs2he+eLuF
bx7XbiPFvEk3MlJjIhM/IP403BS3U3BuYlT1iVgXATJPwmvKaUXWhzcgTIjs4XaFutbJcfsktmZf
YUApMe1jmnzdy9IErvfBISaTvrd7H5PqK1OrUr6vbQGt+Bh06WiBNfO3dLRZ/FSBzgQcwcjjC7SF
jsk6FbW9oEbXoWN5lwTEq0Bc1zl3+OIVOuUdaRWZuJPLzbasdJ8n1SErrv5vK5XwmtXtw/taoWZ+
l6n1l8uF9t1XAREk96g3tgRqcI+lR0mdm34QoJIgepWj3qUFjaDdnMrJIug5j/tlNwOuYGpdTtXm
nknuR4YmHMretKtwPlnI1Ijcfu4Fn6ivNmLjdRRDY6VWNcMpATOPgUuDCyepO4EUdF/+dn0KPu8q
KBtYYqCT6QXpsCYXagnei3SXc0iC3GBPsqYaCHMy9+u+llrsE34LB7l5YauC2mvJE8Xei9SxgYB4
Fdj2nMfCLfQJ3voznd8G9RSTcEFE0Wrb5j3Ytg+8UHR1deLk5z8VWsRStsRpQucN7Z3VeEiCc9gT
vaFTIU/DB/u33JdFE5NsMTmWVcDxP+yUZ/hUj68JCuYw7WdjfwTeAPAltuaNwyvkwq5SbjR1sHJg
9F5aJHCzVjgBcpWy4bBltbRf5C9q7zlF9jFBwfiRSUCo2xk1Y00zs1m8o2NjzBCocsaXcUTpm3oD
sntRChY0MYwtZx7GKTj1TI2+q1sgLnqO3QPbjwi17bKhLhKPbZ+BJBfsBgHgG5UB5/Zut/xfHUN1
CDPLiGFLHPSsPJjHT28cQCaMtjCHYgMPVLAO8fwio7D8ypehs6aBnIk9HV7I9XqCrFltt4/7Heo2
VSZ70ev78QASJ7DbVJ2H0lRtK+g99jfumi2j3KHyvMbvUPe0E6J/ZKCpNCyDOx0QL9A3wOfCDNF+
rPy0oEgi5OafrwKAjYlguit8f0FvVfPrhot379WmEmuToapKpzCOYlrs+E3YL1Nhoib5c7Pgt8hO
WbPMabdhG8+T7V2rpgQmaFG4GHQxpMUdJJtPSmJQVyj+xSSlxk50BUVSmq0b8tqN7gC+hZ9oS+vP
y+QSJrRB+CLJMhjEUboGmARL4OVi6KnfP+NgJ/sPSrOqMxebN1mHwr0tCvuxHynxv2vM7c0gD1Vb
L7PVp8jpRkL6OdWGpqNQj+wPRvuJn6P1DTaPFOdEO3j5JaF2S7NKrt3Jv4LLevjCiYiqSLVdaOfh
ZzC/StbLZiRKYB50GH9lWAwgk1uiGmLaUExSPyzAOvnx3hIc1PPRZ5GMZFoPML7MuM2aX4Gi5gE6
D4WdBQMc2nlwE6xNuc9TPXj4HX24t1S8musciSsMvmQ0fza/WM1MCjYLpOA7soG5tRR6yBg4T7XY
Wq42SBVuMJ4NzZYxYGayg85gGQHyT+dY5UGavZELK7ZvmKmheOY0rRbe5CCnASoLN98FqvaT4Rqq
n/x0RYBhDR3f7faPn/LbS50L83nvari3EYJkvJ9U6X84iLYxgbdyJ+T/AJOH6YLUlayiNFMdSDxT
3VEVbRGNG7bLxSSCNB8gPd14OYalf9oUPpFEVjd/kuKdSBd6SIGJWHuLzaCVtrdibqQNuWEQ/bkR
tuJo1bGzvPjmw0uUyEfipOdfgId74QhuDikFqq9UJDbWHpIhThd0at3FNW3L3k9FN8jbLJRefpUU
05w4McXNoa8EBijJDmJj/fsdCqh1ik/QNP5fb/tvqHz+Gy8+otB/JQyltO+TyxV7ZijKxuIaY08L
fvZyxHIkRO8lKTlkCgBpNhq8rVZG54LXUBg/Ff5YKH+MDsSR7n/7YdDaULn5+K635SlGYQE1aaXX
WRYrpmWhaeOXF6etORwWzNoAcn8sFk6TH9BThS57PjMpo68w5dHlXEX3M63sc/BVqHVyEndFrXHO
o0tIlCVopBorFFFTwnirRfxjwsVtZ8be+6O1fpzCiTSskAN9/fAONqjf0sAuG/zwal2eToeKu3Nt
dN7syyLhgP7QTv8u6x1h6KyYMuQHl103wn8rDQVSrfUy79HYE3qtXi0zWKb7xUHKG9DI92BitSst
12VeolDR6sPDw6IKrhbDd3mdcoKH4GjF8k5mAIQA81Iifd2dxBe+v5Howlu/MSdOW0hJR1Z3qV8+
6M5h3yUz0/hc53oKIx0T1xu5kIq2e9CGuGk6ozR6OxDZEXqXu9kPPpi8uxT86C6FG2PPoLgWimdj
8SkBCEd22KSz4t2SmEiH0yXlaYFXYFKixYXJ5yGiBckf+REK9GvYoZy8ig4H2T6eT+NJn0ObWJxH
98y2FTcLdRNiVn+tKCpubkTtHQaPRGDoAMHMEoDUMbYqnvSGe5qr84/Qx2H/bb7rSdAANByY2P+V
6Ago4slKKVM7qIv2c5PPRifv7KeGmTH9Xg0Y8KN4/dzMGaRMauii3qJgmy2ERwSJCVooZ2njhUOn
TlOQLncPZAUfzyz3CBOwKifSad9Xu78IYtkwVjDd8eyHEzKnYeCTb/sfSsRvs1lB8j/lE6aaepbZ
dytPEz65QMBI6HYcXOWdF17ciP5GK8e5wNv34QKDZ3qXRfyYuBc3u0/i/ztWk6yK/fouJWzOiwMf
aozXDQA5eqhu3oMhhj7Re30ZNAGbWDeuPrw/RV6WlVdsjwWnWkNgXmitlcYO9NX/UBYZiCcT9uAG
GzNv32ADWkl04Pa5UfZjUSKw+No5vxQn6sCDnWHbRIV6c5+gkNwRi9CyOT9/mZA3iB+lp1SUKeA+
GGbBTnLJrCmBNmiU0lMKjEwXI7VqoLKOUhuB/N+McLvM/YbXtS/5K2qHO+IqrIh5QM2Gc38yRyEG
HedUiZ2Y1u0R/kKxWFdLsGx2ufKk5Ost2M1bdxJwIW/2jXW7dgFW150yiGsDh8x0IJTCN8DxGn9l
+PYGa5de+R2Vx0ShxXqCQfxG8KRVYO7TWeugXYPm5c/p8BXpZDmzReQv/e4XPFWhCVEaPEZRYtKs
2dDXoJuDYpmnZmon1DjJozFJTvuqhoGTyd/Ky3F22JS0B1HBQIu8y5Jrfu0izYFSQAal/GXPNoKk
fPRVWMuh6xaXzogoR5JbY4OgeAflu/h+swsbat3pqFAJRZjS67ck9Q9M5zGWYpniUZrnoQo2j7ec
1/6TkM8LMut1nENoxuvWpiWI0x9SEkQucYbhuJ3yYash5Dvhr7Yy0jt/COJMLEhB4sbZksshiZDE
ERfrEExtFhEUrKZhkjio/k14zPgUprKHZj8nCxIY8yf+ZCISziomMpHXy3W7sk7OpaaH3SUERP3u
wJpsrdiqa8gjs2fSxrqmNJusFpBDhpL3LZ0YbGTu13bCBIkZuRVX1JaIa+mkXwSkN8Ay8Y5OJhZF
H8ZxMNpWWhSTUQWYijNiZi7YMci4sxEHqnNG7l5lSoOiz2mFhLQkNi0XXm259Y50QUVR82uwp68k
SyQNynv0OQ0QsgTy5b5NM4ZcJCOObtlQU0bGMo2ZexHc9Rf377+I9B+6dTfd3MhGkbUOs+JCWk/G
IfaKsg627kFnI9KbgF5WJA9hay10cJEQUhJ5/VjE1ndA0vXlalqb8ghowLt2SLP6PMslO1cmLFsl
G5sbK52tg1p/Iu9CQ25ebhnPITY2HxxpYAmHjRtrlUEfYJIL357JkHK9peURIcD9FouN5l088RA7
zMh60EYD5gxtj/hiX3+O/pamdWy94bMR9Vqd1LoXU6jJTjanXFr/g44+7uO9ha7U+MWz8Xx+3SLw
Yv0MAHhkZrrSr5rRpiftXOuqHvdu+lr4SThS8N1wGq5rWNsynkHvPkom8qviHlgOUDTChGmtlxl7
VHTCqeIpmhN6a+Qj0+Y+cJAuf4L+98NSq2AzMR7wuoUjvfeRcwdtbtslgD/VRvXP/zvJ/YPNZqgn
rI2hpvB/ozMepV+HrIDzyrpokwATADxki9XdKHI3Tesh0MxQMm1/4wt/jv684fAzITs0CzMp+J7E
CGsGbmAmBnwjkivhNozJnybdTCf7wyLIreAmhvoAschYRwt10RSmQ17IAbM44ECGdEsSz0Aa0V7g
qy5nEOTuBhqrSDUgKvBKHMPfpQBwMTmS58jD4/LEqUknx/TYDlPIJ7xVCS6iewzxvzcZ7k1S4lkx
MFxPL8orWeWqR9Ik/klpYLT7DLo3PQlXmyRngKCRZQsukVhDHhhRPXFAg6WO2YsWxpBTdTENg9l6
EiDPhqA0b6gxkLDrvjcRgUE7KjrGU9d8Cp2t//rkftBaI7oUqyd4RmMyTL1AjuAVrFqTQrk2cqzv
40el/bKcWOFSOhxZ7fEoNNTKo1HXwVnNvyM5fqeEzbYWasMmqshGJ2t75UH2x++UZymz9pW5Tn/B
MwRqNLLh98VIdWJBlWn9amBeT2HLJ4xDfykYR1OG2p5QdYmumYnNK7shNpR+LB9wJwFDuAaWfH5b
STdZ80Km1fbr00ldc2Z46VoCUaJ0jidrWKDnKQJH8c6VnMsDoAFuEK0bc1tcmQxBnArM/i01adX7
Xg4gC/TemRnrEaXkgvySLawMBb5q4CVi7Qd30YAk+iGjAlT7iVvhhAzST3qp/zoh2KUFCxCrWuen
4Ury3BIWq9JoRc20qJBMTiYBhcJzOqZrOC4KCZyMnWjJO1bU8KfNn4yzionynSc/NW/Ybsd05/T6
Vtc+pNTAJi39XKTA6F9OO7VGVavSJB1T2QOkt/WEVG3+WMVeGgAfBg18waBydgqptzGhS18xScii
GemqSb3zA3bHdcN2gwo2WTd5Mnwb/C/BQSL+U1t66VzGBPNgQ3FRXFg+gLlZtndSft0BjxC98JXe
XgNOcL91b9mh+nw/b6LY0Ip6py909a6jyBY1PpXEoVDajQrWU+Ez2xCf8/v69SDctfjZJc3Ghyyi
97L10+l3Ic84pJ2TaD1Jd/doXAXhJI8vLMgGl/TH4upr6JekjZPNjyL7hz2euQ6dc9+D9FWW0/Bv
jzql9eB38sdl2+XFScnmJu9YYcgLufR74+1r45e3p8bVp8Xu+TbiUk9+r+cO7azUzuE0WppX6cbe
2S/58HFW0e4Qb5ofUYoP+VDE5rY61fsfcd1YHRbl5+2LD/leHqu2XNE6frHKCWzMC6GUkxX0rXUS
oA0WOF9yJUZg0lSMyCbTaGOeQI85dEhLRpcfm63SiEpyLzFCbBRr7jBfoTLWfUagmkOXoX3OMhoV
1prBd+ebfgvT0NTlEegKxI6OgpPhn1XwahrFKIHhN486Hltt3+teDlkhGN8fu1GagtoOSdJe9Vai
GUa/4Jz85l9v4dYPpuLcQ+I28qqs+CubfN3rL8Gz1/h4f2fmHD8SUxjV9z9oM/Ki8jjTQ3EcGRcx
wonHprRzqWEUkTI2iCoi/bBKrZqkcLYYRZsVslPJDrh2sycc/0GfEhY5wVmZiDov2Gr6j1UCjhAz
+sH5/zhTenCbNRtivbK5oruxNAuFTj0NS+OhSjiFp6QqumLQ2ySTVLZr0LnHSbYjj7XWrt9ulDFV
NyYFPA26Pmx6Y8r44poHwvZISgc4uNcjKS4EvWPGD6rfIH1Bt70FGpW/hksDhTxxyJwvfktyGXJd
nWpP6Yrc4+vIlkuoNZ4y10pCNa1iPAah8XjBom6sTasjRaOIdYFcYPRhXZCK1QQNkuVmYUiNnM+p
wwtCxGz3rX4ihwC0iSC7tIrxmvsqAnfrQD/fJii9itJcgQR5IY89sG5SYJb+hM8UsfhchJDwafG8
vLzlSDZKy6/N0kqNXCvcl2rd0ncGPCphcwZyQt6zsN6AOJiqlY3s8pxo8xx0zO2BD6wRZ7bBurQM
H3EmPVOimkKg5PSRJVOSL64N/6rymyJUB2ZsrqG8RWXowWQ/WIkwxWiJaHwXhsTZjQMcdjiMXobC
nzOugxxULFUEudqyD46crQrzqVStQJQ7eV5ybtKKen3uZhtSVcGGshLgAvWM+uh0tC2roibVr63N
tN/1D6TK+IBy3k1DHzrCgqXkPQY1ClWeU0rPFwZOScLlj1k8wiwpAj9EAXqDvlmQ+zz/ipoElovf
XAccWW7Z+J9S2JmNYUhHkFoNZnO345AU79L2crSYArg2ZmcQzWiV1s1NbYFtVDQTsQUhIXAhe8bJ
C1kAdBV/zgHQJCLJo+7h5B1nuZRUEiedpQvmKJqF37/l/rsYsgoogAz4S1kJhT2FO+EQMoF2vDQK
yc66/REWrTRoKPtOscy8PNPvzBS/EsrsLRL8KI51W1NY9pwLp3nmmfShuMKtwNpqra/bL3ojC00f
EWr+UfR6kL+QAVJe4m0RXKpJyFH2xdZECen4H4TiLw/UCvaMrkiQmKvYQ0Uy+52iY337ILwG8qwB
po9QEaJRhUfHBXlD0v4v/dYSHl+ClpEQZdQkWg9S4JTRR8ECY7qnUBqq3rFd5RjNMWlexAdXUPqA
7eZiCj+tkOW85aiC8jddFNYbyDIf6eOcT03+FGIqw3x89fWS7VP/9PmmcCg6QW4EGbCH7dYVXC64
L1izV80THAQt8FwbNyNy67Q2dUV5/VnzyEg9eL2jqykLp/pIdd6ziLgtkIVjYxDRa1myt9BbepQU
f3Alue8YyCCrbOhMHB4BYKrfNFzOhhGTPO2a0qESjHYW+RXf3GelWUGUvjq0jiTtJW6AY6kdMrYw
PNzg54tWaTO+Ms+FtyUObGd23PWKSqYO4Oi2TWFpwkVGI2RwgoYebIaBRBBHBtWOZvMy/RyjTok0
E07HIGEhVR4jPYHt1t8Q6VDKJ6Tm09VOZqu2N6P97qoA1IOo9rWOw0FKkOC70Zn3SKHvwRskyE65
2WCdm1A8gjeNWp/Rzp6lMxlWRjDwlEFCaXHEgKw9ZINVIia3TnfEInQf0UeCMwX6ybbnEF9a5lLe
cmHDR//Ot6a1VznJ00wOIgMWP7PhvliK3OJ6790MiyczmIizX2ri082NrczdpJf9z6WxCqKcfmZT
PHwrejWn4z+1u/1pyL4xkvxgQ/u5BGUFZi/GYTxjSJiIimewVGtsJtSIlAChxyQbSHRIDjuGIXJv
xbmorHe1hpA+JGfdRlKM0oI2VjqB58Xs9rNQ7MuYjOIwojvjyvZCJzn868w0BZ+tNW6HKm5FrQGb
O2HPaWFYoJ3XVHMDSwwrgsgFtKCvaD0c90CGCUzinQSkR+KRRGSxZ5cRQtBtowOCDt1hXVdkF/x8
bAuikGKGCRvvId1OFHj4TN0MynxouGr3nNSFDxd7/BTmxZyQ9ZLMm9A78AC3th0eRMISWWrE7m6e
Lk7eStWRxj8vOSKAOL1l13hp3YdKhSb0UygrpYD/ZxXqo3EjY5CCZ0OZcpa5GMpIVQORO4Oj+50p
kYMtaruxnKO6TRuyXbnDNm+sNK/jVqFwkj6WCSO8yaX4xm0Gm7wZN4ibtbjU9Ff4fEx3CT5ecrwP
G6QsNL14/nbSSSrR/z4GQHTCIE7wSo9HUN3vG7+g6hbfAhCt+1PT0S/rhdAJyLgRtoOUzvLYFm6i
tar/QZBqo8nNKHWPCIxh89fVdC2bMn2TzwriRv8z6SgzpFN0WBV4Lu9uYqk61RXYVrSRzVqV94Zq
BBb9QftiNbwc0K0qk7qWNmHitaICHX+CKaGBF3TYdtQ4UrU0T3yeRF/qucipzXOQsFiolXQ7RLIS
XnJazlc+Rjzhr/UzETcP1hjNUIsjuvjDvcmGO5O7DjtiGQ3ut5UIkZYM5tUrzGQlJEkgAZckyLuG
vSQuDAyhWw1Tq6FHODSdQcGSzKul5M7xRA+GTvkpiGXtpiIupzd+4kCFcOzdpMgEeEvl9k2hCJdN
CTklSKlF0EkPnS+xTaqHWKLyODpfsxRucqmw/B/bMjot5hn/47GL4ckTSQbsVLeZIenhHm3efzP+
oAI+CyTnoeeqWXVO/BifOgxtzmJmpVnbV01Vfj26YoD+jDYTblOj/GHZPuXyYSp1mZKSmoVAv1l9
hV9m223yuXVR/2t3TqoSFY7jMQRsyYR3MOV9TFPl87JZwiHPNnQNv7ZXSHYzdPIQrrlyRfzt0M2o
IHBlAIlb+pC6kmDEmqzTbDaJmkZoU+l//fgKdNmgBLGD7cNCC3i6i1E9S290a7S0rtJ6USfaTo60
HCeX24ED4hg6A6HlIYHrd/eha+Ta9/JnGV1eVQB/t1kOlJbNNQVrreu+8UcdQX7HHZrA3Jwp4YoL
VymKfxuAc6poDPVYp1y5k6vsPnRjowv4yf44mQffkq6cWFkDo6oDtAjdKSPiMV9GXuDiKgQt1tbD
gmotDUHbZ8+rj7Ou1c9pa1+v6dcds8Ir7IVgGrHqcOBTPHnQIh9lpPYfmvxIgem6gJLdwvMWjJjL
rJIE3El8GYMjtVufO1rwRazF65xUtOeMfASavDEjLCcboISkveTY2WHROmiOr7SSE5Q/2PK0V3zC
LLCVHXfVOuxcAWNRZy5PJRKTpueC+i3qV496DcjkEK4ozSdHdd8oNQJtKYF1DQC+l2eX6t0jHf1B
LD5k0xQP5BReW9+j1oQOIMtS/178+BQPz8d/jBlZSlLy634zj1OCTBoyydOzLHy5zZ0EYhADOWkE
YTNZy4FygJRwAlJOwh3gHW+ACz9aolvhbXeKHA8etsF+tKm35S8fl8I4fgtVqLj8vyVKiczOjCg7
gD/T3JIVcnOuznAdPVsrYiX1GtPwph/2Yr4z1odJ7Szo0Hki7gye2IXMsEyqkjW1EWnYY8VuCgWB
MS8HIJZns2MgjDA++k8mPYw/zadbFK62YX/0oMvwt7w8APw06dDKekMopa0nhG+BCxJWBLR1xkQc
Syip72LpBMhQDOofanWcW46wnt3sna95jQ+wRCTtF+YQKFMva/augDxlpscu5FW6WCghoBKaRxlh
fuJtcZM1iIB8x2/24krvZcpZsTknZN88tcDnab1kLLwEpRofT0ui/nrud/VmhLPn+jolZmJK5pPp
cGmLlbwk82+FcP01Oc2RUcy36Hz5uh6jlYW74ygqgQ/DEhiMGpSAum98QLa3p8ifjhG12OoPBewS
Ti/P9moG6alhimMCnnXcLYRf3TL99ElaX0jR12Pxn4dYBpum9jbJ3iXlEDr2dHsLqqooTXPvIfTr
eTlAmV/MWmJg90t7mp0+S1YdpTgdAnvEWXrqlqbBaGwgtkHhRAuSpOE2nlWfyKrS5n79RX0trQlm
9hWXyIYOTeTo5wju06yTETYskOAa2qQVKTjaqDkhQW/6kUHEEghLjiOQI5VcoAiz/uhubV56nhrO
DoyH9ZwswY89pksYTVTvurWjJHH5Me4XnzL9bu5ud1hAZ5tB5IkmAqYLMY6P5TughqU0SQpUHiOq
+sx72mwWovqhPt9rvvSNbyRxol6ZdxEtSxBFJZhzetb31QG+raHx7TR3Tf+jay1RseohJ7P760u5
j9pYsPgKGaZ2czllJWHV/TZz7YCFSFtEgkKdcIl5+umbJEscWivzu94aLSzZ3B7tiJQ7ZfALX6XB
2LUdULn13ua3sGx+HLvF8zr+YuA91Hr/92wmhkElkGRacvz0/8Z0BQ7U3ciXZtlBdg4Me2N/bzSH
Je1GVczaKuZsrEI9rkqIIyyBnFSQ1X51RtXuzUd3P98o+cxjNCWS+aGNgrPcAA+qYDpoRtMhaZwq
BE3jKDir0RbJjStKIYE4uzvBI9thXj4N3k451yYlpEFfVQQPoqQ/R9W5U/etAZPYS182VNwYh1eA
vaDMo2FNJExUECyT71dsVm4UpnWxXVDD1xjKgKC1MYlb/xqHmrp69YiUrDCt5fVmulCE591v4WqC
RP1YzP0UeBzWXJPncdnzx9Kv1qHBbfj3u3OyrFGxOZmEeGxOddCybOlwA3XMqozBRkQXolzFB03Z
9UiTt50JeTIIe+U7+bhcP/PLx/oG+W2AIeMDt/nItFnFkHUK/YTWg0OCKTikPJdVFwGQnfDpL0XW
557yciksyCBCJch4HlJykCntDWol2KuBNfOd5ljIwEtIJHJyueUSrevuRkhMn1Br3SFGj/hK5k6D
XHZEILbGtSgPZI1BC+Zg6pVboRmV8Tw9CP1aNTPnm3j7y8SSRXoTN4lOH9dt7iNYn48J5kS/5LYC
tbNVZqu2P0Sw7qHUNLIEoWVs6oigh86XgHKjkMYvtpAk6E7gdH6XRBSagTz518IJTsAoU6jDnvmr
XYon4VJiPJhWqL9WR+mS+W7DPKS0d6IVZOZhs7L/harStwjgKGGQEJBxUPitnmTDHCYrOtfM6pP4
D+1VEBN+zW8VlgZ1tRp5ju9YnUrLYzxktw2fD0yBKQicMHlVHjoNpWe4jBk1Gc1z7IBUN7z3K5AG
knsOTO1PFieArUfTReJ5vwIZLa8Omv1LGTXi+S/eJFiAktNQu0cQxwSwj2XRozmb9pWKQIdgUpGa
dLG5sfUSh73G74sGaSwcmKeatOW7znabL7Y32eeECCutv6Z4PQfChnlQ8VGhpV8CBOGf9gonv+iD
NisWEpw7OnBPMIGuxyr3Y4jsoIOzX/FV8X7699AkO6YzmerjJfIoyebEhzOb2NOzPl6Y6k1DudYu
z8Y8VM5IBv0a5QQm1amscvUq9CN+HTaVqJb6Ts+kBdedtb7o3bMuiwMtm+BfMceQI4Uz1asewoAz
iFClCPFeEApk8jtGnRW+Ha7DBiDJOvIt4G1fIRW5Cw8XrEJc7pwTvnn7BzXCJ/3ky4wBVovT+ZFB
uUjfXXAn/02xmVDJzWnW0bJrQJhoAFH7AHwKGYJX/4cXKVywStiZRRHsmGhHqwOn2+csSa8Ynhxu
hwqTzD3R1F3Tyw8VPGDQ8BSW7S1HcmWOAqs5P2LpvMAIPBmecdmPzjNPZMZjEy9wBbWHyvmpTNvz
M8JF4/28OQ+3dppOoFYjF+k/T79zsqV+/5nA2Xi/TlXbtIuBFYqeZtIXGZbwIUua5uYBUzrfNeCt
w4NupvWJ6dyLbt0X2MMq2ifCLW1S3sMBjYli4r3E7hSODJLnSLFLPsOZdJjVzG/e8OaO2E97rdnC
sLumQ5VMeb93HF21xa5PRLK1GMW6SUUv/legKBDHx2MwGfH0eyzckR+VyGnn+a3E4tBRgd2HAFnu
VjzcYZuwrWvhIGjE9cO86q15TWeUYugyf3MUaMqcl3vgcb4Q6OhpTqcEJEh473DXIlLjQWZxb+Xo
0SuBF0BDGWTwUSCBRciGGhL+FX1oO8RdRjFlejV5ol0dOBRFBN9XAX1PQnZK7eok1AompxVZHd0P
/k61nV0nxI/ZcmMKvbZ5fGsDw2ntjeiUTq3rQciJSHxuZcw4HMDyLCnYqk1meSE487jOJmJ/aVkX
6YNMobgnUqPakglejOHMuC10EAfh8rsx+HMTmmI2h9jkG4QLsZKIOR1n2U9ZGweD/V/pUVqMvE8P
6xchksHUCGgHE/7F1w+3v1ksvq2CKXt4mcsQifrec/FKofCoTFDDZm9Iq3GcnQtTPOvRyTpvwZBk
QxBQmFdKWgSDROW7z5G9mR4HhhCZucfsAuL1lW4kSE4AY9AGEVYwjcQC/KsaB1fHtYbIvJzbii4W
p81QYUejWn3GtYg7h2oyI7Rd7hFCqpQ5XR6X4jDi7C54ritBEMS0rvWPLnNdDEo1q+rVsbCy+ASC
qa9wNMqLmhELH3FTlYTXH0C3D27PyUxozgQF7MzaliJru/m7CIYjVRuh5FgUgjJFVTGs3gaw1u3L
ylW52FQOtn60huzwSsFhWRNPDoJoVWTxpjeU+v4yafnFgjEIZgplBijY474dIUDsMvs01i8fiCgl
Zw6PiodCp/gK3mCyDI0gHK/TeHjjbFqdztxccQwjI2JYEWOIIvRY061DsvvaXyByIhlwyD65i2BM
VGlKgRtsOF1yEe7e3PrQy8wG5PYTQk/mXlbyJD+RamFzMh4xPdl5lK263juWHhDe56fl6w6sMBB8
VM8uZhKgcAI8jEri1vnsfxI//+lA1HZE4KC2ShaMPwzqIpmuoTdm8zOtAd96qqA852hkRlWmTEwg
S5qt9m401uM4rAU3reIO8Suhzm22ngJyXzeEyyILjlKC6XQyVO9IZ7LgzJzqbyKBEzzRu1VctiJf
02SW8UNGWlgh9OFhkgtTm+mjeRY2thzd+47zdf5YQJ1ySQ2qef7KkM2BilqEsZjqkrF1u5Ck5wXP
L5TGDBud/mPlPKAVIYo9OETjDiSU45ZV83CjF0kVAp9e2qZNQC+5yOs10rzj4Trb8nZvQABIW3z8
qVE21+hlDgbv9kY5UQuH+lDBmKpOnZL50I7VbAMGiuEM5jGoAlGU0sez6/h7nvGj8Y0aL8Ehmnwq
6wSckJJIjl5jehXn8jLgjejav8QoRvmVgqkr1rYDmu7n/Bhq8oEqSTDNb8L4W8ZUwahb3cH37uAY
g5azQmGD09Q4OZ+gz6U/IAJn77++qWemG1lPdkXkcUwJQHVFXQGlUKIcUABuCEPmVmLo4CtbQe/D
Sa8rPHSzeEQ+EDL5OLKKposjzpUw1UVR/ma7tdcNUXKZTF+DcFekkwoubffFS5+bZqxL0SHoM7KI
stVlqjwRDq+nB7pYnHCHUoUggybbirKnHxog0Ru3xNbzXxFIp0NN/jkFTvCJCFDAqIfBQvIjIX8j
kDiBiepJlR1tNhc4GSMRa/WQRrml78C6MAg1y1K+6+qxw3x83Y4DJglPdEZ6ZLI3Mb5fThTZhjej
he6RaegUgqV8lXi2KJgOO08uMDvgxkbrMnwIFpd4vobtWZ5vvkOA3fh5auXP6C3+b2kruWnHvGdp
MVqo/QsYf+5yNSEWFphK3KQg0lhku5krJ1K+LXtU6mH4rwGmRUB0wSGk1IvosoM3ijpUUTturpap
Fg3GM35ZNnMpYaEtcfV40mp/XPUI31Z4YvNf9eGfhVM4KB93/NGszdIEw6kYeZdKnoY+oF3fnr+R
Hq26oiSXJmKK6kt1kV9XIm6hXMFH4dKuEl9oeymJrSHcJhk99rsxxq2DgdPusIocRtVvWZtqBQ8d
WYsku4BMwgTmYx92eGh+W3FZcJC1KooYvZlsFWeJv0AkLcZ2wsVB4k1h4w3oC2uwTWqmglfHweyS
kKfebTxL6dkzSoIwgyacxSlxbdqnpx/zmjBtDoU3R/2286xyQbdYvP9t6acGNxmjkiz1SZLIR9te
PcyIO/GRcI3MHnaiVMVon3nr7W+GABmQ3C6ueIK/MLtloLkXiTpHVxwa3Jg7B4Q9dtuK88XbGYmU
0lB7Es3oHd3kQ3i0mqUHkccpEoo+I07jBXMKyS15PmeanLyuZC27tpsxawM/v0CzVjlYMQsjNU0P
KHoEYz9QUbZmy8TmkvkLeUfy3cmQg4tOrnxkOpl9wqUQR9lFPHOGM6DWtGepYTg1iNaxwafuN4S6
ZTYusH2nbUp5YqAYVDfmGc5Uf+VPWu3WJK+GZQEGf2281zmR65u6Ky59vs/gGyuLOY8+OyYFhidA
HXGAuLXZhfvHRLWBW/R8JL7firq69VNyygyPhqBlwBOFpB9m4X8nPdmaSx6Bp/upsepyF0vFfsBh
nJca7l46Cf7rh0YmXmqhkLogf2Xq8XTZdJXAzxHfluy5Ha+M6H/mKk/bLni4Li7n3mjY4vBHdHFV
PeAp/sOCumCMDpQF8pOFl8cFcRRL65lo8axZkeewPjR2ft/t4ujOSqQFJQ4JIqihJT34AzSqWeTz
ASGoHrHHt/+YaM3CU8nzgz0qsDj0d6Uy/GN2J75eP2gLbSBvEeNiweh2xyjA10sjospWYaqcqBz8
JWpIbK7Wrv6Bj3s2ulgfSvIgudFT9i47ZwLChttMO8daauxt6nV0fxs+R+mSKkS9yv4YAVrhmqAS
qOvZKsEqhBmD4/qePCKM9bMv72yXIMS8SoahET5L8HhN7EDqVlmsWsxucCmeljPSB5sqtxN3E4Ig
Fx8Fs7kWMlLB45VRIZWn+qoLezaoKP8cNREG9kf74+EVMbLX/rcPcxdG6PCAcXbFPfDwlRXJ1cgR
1hxLhS1XrK7xfyf520rwBZ0pYlvgv38T+PBBYB6nloSEJaxg7xR4x2jtdnmyLZLfi6MS55gI9a4o
p5ngscSeMP6xZ4N9tuZa3XfU5RyUoq8fK2OZeCWA3f6Qq7KAZ/KqSLqqpp+EMKwviV/buuRNA61z
rThFCdwokGdPAs6iIji3Pw48CfAxoXpeHwVyTdxfFy4q5OlK0SWcStJzKV2+hkTLbtYVbeh6c1pd
E89ujFKbvqHNZSf4buUWdEh6QLJ72FzTOaWs2q0YAAgVBFDuMZK+McUWwCdrGQrDf1RFSRA3K14J
f2+kkVVQhsjONs9LbIAjGKPivUSRyq1HN5/pwrgoWx4L53G75d0vjOTZaYaNYjz/dHiAa/bxbWHu
HZMgjzixeoRt9WL2uvFrPY65LifMCIXyrRaETRnCAKVVuNUlNdfkQKPWNgpma89E8NzkOErWW+Aw
zLegFU4dmQx58aqw3eEq6vTzdX5e560dpboiXIlFkrJE+sCfB+wMoJKnHA2hHQPENnmAGeYQYrXu
JH5vFXwCUPAcBn785TykJ5n8Mkk4ix9hswj8eKrRMe1tY40taq7zBuHqP3FvTQxt5J+BnGFUUVtF
yRSuNq6IkT1zNnmB9t83nNYIjTZT9GpYaZzg3LaLX1tldZDxwMQnEnjdzYr977omi8veyrcyOwuh
1K/cPTW8ydjMQcZO4KFBtQpbnG8LJr2e3vC0hCWqmk0eHRAN7HAoVJgoaw0kSy6l54vNrAgYeX7R
6zo3SVCvcJEa+516YKm1kvH5I5j9PijhI838Py7bn1HQkePH4vjH/sMdVRBJZ76gyLp5ZrBGtufQ
8p9vItJC4fGiz4gAjnCj2rZCLcH8GbfNt+Uy0/xLh5jB1o+lv1MogMDCo0NklNAo0bPFqm5vE5KA
+RXnMRbUOcBeW09lfzMvvyjoKJmreOYjWrUC6kIXqFk9Zf22cDS+yRpgi18dD5bkxnPsPle8zG40
XbNt0Uj6PrIS8fLbzPlvL3t1eHI1zDsXc6Dks19FD4r27A0P5iL8m2z0E90HTTxYTBcmlOI9v3gO
lAYVCBEhBpV2I0dPnMnkwwLU0CS3xF88LdLBg3vhrlCW3aIUmaZ3e2Z+OB4+sXcOZ7/DWUVOcWPO
QsIu7SjLKG0yaw0UnzaPHGvwtFfvngP8FQrlx+pSanHryhrkekcKDLBwvuDCUk2ROsUJy8ZsxAhP
cw/Hsg1ZoCdBq0NKd/V6DKodL6ekQT7vJLUnUiN9SRfW/Un0fhiyJOCAjC5QMX1Z0VUBOA/J8LiN
x8PcTfmMWfkKS0I90hhy87sODvfbRpukf0D2LBtm61OJndf6lWYtjzGtFrt7Um/CufCwOZzXCbP6
ysfjWCCNYU+52se/eQL7hpH7V/W1lvpHMkbLiDXU68iZb1mRlopskBXYer7+o9nhJeWWIH82e2D/
EbcqPA8jtIzdpkg0Ip/BarqDLObfQdye3LHo7p8sY/VDNSXqcxKEkSgZfA8Nvn62Hzxy3j8ExDLs
HstZM+p+6j5ZpHPXNOTQHQHdJaHINAa7X2BogUlDDu02eIIIOarQn+cpwAIrT89+M4HGHPDNW+v+
6/AsJeyYj87KN8yTXCyzK7BE5GVOPmhrp9CeCe0WC6BAftBk4tRg693zPNCg4GPa00+iDPFoxZuV
kM/9V5M7JouRAjlEZo22Pi1Cb6uwwHfAWR/goAJZzOclnthmrCbDwJcSTdNyqUed/4LD+eKqgJhN
AGBjj+t+KMB+aVUYJxSJCthZBVBbd6LP4oQqi5HnTJp7freMeacJ4uDj9cQsIPdUa33HnyfBzlyr
sn+P9ZixjzAtoFNfCi1ErJ0DVtjPPHk6p7CzJgWARtaTnHkMRwmottjL/pBXVD6401q5kG1Kln0q
vmzlIN2U+5J8VYesVWJZC9W6ojIVHbK7BFCjf7pnnz83zUGRfuw3LXxK2Ze1EMinQvvwxl5R5LLJ
YcvPUijhJjyiSPWR9rUUdnE8u4VD3c7RUgdlV6a6Wloj6jjiiGLNNAWEd4wqkeWMk53bZqKkLZcm
1J+6Zdu/qVVu1gZ2WuV8PqTB662czvsolPY8mle4h6ncPlWdGVz2hWJntzgRl6mXDDIqezPvhQLI
jSzk2x92tTltGgq2W1JRGd8fKl6VSYR6MdK+jFbj3zfVtKsz/ghI7AubbndQ8jf6ZUQsDwzaEVQ0
gZiNiijXTWL8/lPHhFNtSQlTJCJrs9Td9WIDwycOceTKBwAfsAVl5jZLLVuG+YIun9X+hnpChsB3
OAsn6oemF3H3reM1V+aGt36o7kFbzAKt9nuScY7bmvF9s9V4PL2AxZZ5GprMQuzfp+kTwT3eIqtz
3ueU3Emz7jZSJoZvPacaAGu1i0d2EgwfP6XnHYL9A8BKyJIuBggE3RwIhDvIRqyDJu3xa+WZU3yN
n7QEZe5dL5CMloYRGDzhXoarLNZB16NJI0qUFqEatV6MWI3p7sWGnju7h+AKW5AaZlLn0L6hP9je
IaJvQRgviKTeZNktnmrg3u1UZSI8tWQMvjwgv85hPy3voYuADAvJaO0tgMGe2yqYVNkAtWWDJmwd
Z323DWb+JrGPl5UpWWpmoZhg+dPKiV8/QR3VkpxPhBa/cqeexOBxrlf6X3FmAkx+OLsU2vYuQHAX
hcS9/jGOwQYdFfPNls/Emd6Ui1juUgzmEkb66VTscHMDrejpIQvUU5Q+QmcXqm17PQ3ut42fwooT
cXdA/RThRqLiDastuCGq+5sVNt9R62iVEEyQHvG8RhFJ8DIkt1DvcIRH3OJVge/x3WGmDDjD0IEs
ECjTIhxCNHXmN7d35sdSHp8UhnV3E8t7d/6vPn/agy9JYiOLs9B2al0hYy8GYEc902NskzkGN0zA
JiDLcucYVAKZnjgICblB/B/AQ/fIwHP+Eh4CawjrtNGoM69mMfm55xJCMzzTLHPb9bEzXwt2Tnqf
u65flC3RVtjxBVDsHZIB00aYW1jeoXRnVy1mRpWc/Q6MSv2prsCKj5i4tULKD00gdvaOgVwD6nyx
Vmclf5n0vdIUvu75ubwMSKixDTb8bHlE1lc5cZ53MsrClmk7qTSKUlCuiw0sM318Ei4VWFTMkoLX
y9ALMZ2HgVXglXm5TEbSiQskdOMCuIzA9OEpdhvfeeWfK/HF5GM+THs+MbJib03zwgbYcTJJFqAG
pFkUswHpb11g8AcBGWQNi96nEwkMtq9XkEGhXZbtUyudfnaADzpJdR882I/xJ2/t+ShiKNzL4F0J
lAmniOlpvU7IJtA7JCH23ycIJuvejg0d4BJEudAzJd/oFnuXWn82uZY45iFCFJGXHny+PSYOo5Qs
64ZmVdyFkwFLAEuXTA9WCbKfL7qxkCWB9E7gKj+yXmCFnM91tWzZRJPKIk6wLnMVdPgHcl+O5Q7S
fbPHT6YpNnxNVpOaGSrus6M671elpf3o7nNtqEcvl3GjBmQRwQD0AHNkDZlxncO/oYCD2OGkY32z
Sy8vaGe1mjDBA7vkkyaPSICrzg/XKD5Fy1tSQLr391iAGRVsqnsYSksC2tdYJ0/f0aNzp9cAoJXE
Vuu0n4RN4siNlLH9TvflA8wbPDfOZgszv3HcecntuNcD4imTT9sa9Vvu0GcAFTs2HN6Ema9Ji1d1
jOEgiXf+mB2R8YVspHWI+AjCBM8LOZj9IynSFlIxVYFNGRHsJ80IY4VGk1eN4tL6YuAqv9sSV2hz
0t+MuoMEXA+Pa38/a0U4YXlUdiwTVBKWgNyNwU44cmKy1FLq9EtraANb75ffAl/Fc/AciRb2YHik
IevEM5sx8V7ctfv2a7N9KeqF3vj2yI75Di29qnoPX3DpGu77W4gIOjQ1SGcRzc7pICb8N2frmNbL
SBscVN5j4OuaOyMVlBMD4uBB+J4MHQMvY+rbXWDsvKcZDwmD+RWnoq1trMDnoPSVY0JCzHIF1TC9
cGKC/ayen01yj+KSlArhxNuTeT9Bj4XjsiQuRh4qRtd1VJVQES9/TIwINbGbTzfLVlK0cTOfOIfN
tGvN5SYCEqZf9LC9/55FnUUOQPlnUDByXZuzN3WGh0vYM2mhJFDELusn6lND81rn1Nv1EqE6hbFe
DsejoXb1vQHken3bbHYh0Z23ZSq7xdcehcnv5MUWULM6Q66yRN9N+CerrWUDZFkXj0RdGlNfS0Wc
ygbBcmc/oNsVeMftb8d2Ory+xsoe6Bv0ouPfx9POcrSfOWq7HfgXtBrTaf/eKtJmtKfGDv3UHCt9
HnwHxASuZKg1kpVWbM1nSZk6EZKoRnxOESLrcdJs6/8yOMUVndp3MXYmyUG7a21jtwk4xfyH4ASO
g3RdJvt8CemnI5imfazFJ2+dtUoRaYGNTn1yJY4lA1NWOsqItqxv8Fjp/JYe+pGkU0g0lerY6t/M
yPsmUMgiuJ7GTJ7GvTmz7HM5gYewjYCkvsaTHikID0RC1zOZe2Ceu2btI60KLGU/P7sEaiSayk8F
a9jfC2A49IFu3kZCWBf9ucUJg1d9FTPWjLT+jlGrAvbv+zxz4F267NcxUE/5o5CvLBLceq9sLRk0
GmEwP7BCYXVsin5/+aW28X6RFHfUmp7XruAiNxEkNxxQXXYbncOHXTJJ+2Eqaczn3zIBs50guuJ7
YaKe0SS2l3NzObYItvJbH8gMTKQ4o45CvzDJAUp2y7jMl88lh7si4DoYdLWwiD1S2Qx+Busfm2xn
DBd63Mp/x8tOyp0zmfaExn4ZuLjLgOvGDRu+DQymg81u+eE1Co7/G9OCP84LWHg7aHOZQBdju7yC
kIP4gOTIr20i0N1wm0NrbfXb84sK6WKy2yhBKqERXSqwULFhGI+R41CaPz6ySVL+ZjxeIB2iRbv4
Vk0MOmiP1jyt6pxY648u+AIwtVIedZhcaubrxkTrh9BkcJ/FcR5raS8Q7tl4SmvIkdt2B1ZtqDdK
B3BroFDtY6CN/yaC0Gtx8TRXgmK5hqc0gUwVbxY+uTMxXJvV1W8RD19WEFX6YtXRowuNLQ7WeP7R
P+A2MBca0rNEbz9liEV1TzJlmtAY42YhCWU2mBxXKrJxAD61uNMw0kexud2sPwYio5FDO8gklHKI
zaDHIQB8ZHg6eHjGDXQtjcHhJ2bPcZNyhryRofrVGtXdyBGkpI0wQnvijazuQfcHpHRObN6tfSkv
sCnAROIkMmRGV94M+nXT1Yu/ddMe/cew0F6DthJOe/vfy62oAynIwQU5nl9LilN6acYvfbRDORcn
6evvcW96WBoW60B10zAkpTAmDoDjQ3kgO+0qgeR//eEdjw6zzydSwpsY3zk/o4p09Z1YWzdt2ayu
5vuo5uzANxIL2JFQ8ESb6WxT+esEbYddVUrpwXs+ln1wHunpIq3fBwLL5tr0xiKkQJZPg1tQfmIX
DV5Ama0WZr4KMMzT2vGtjXDuK8p8i0K5Rk2GrzFEQmon3EGBx2wHHcT6kmBOp05DvhKTyKnhWEpe
j0B051AVfOX1eipA6U0rmx9jHxYDTCou0UdrX2E5f2C+09p3X9MX8GW+HxWMS13aduAAY1qjZ9Sc
DLVLuk3bRQZfphbLoLj2Faz0CSqto9zPx/REXmz8pGcG1hDE0u2GUt4bCTqD5AaU9BKMlo55LxdR
yUkxvxEB1fvQkYyqWyE+rItie5vaQDLYn8StKH5IZrZgTv3K2FhNRL9H3pqvhs2lcmEh7C1+9AuQ
9EhkK8SrBui5YfYm3N6VUEu5JsWnYxG4X3u9qR7waF4j2soArGGu+F64e0GknrA/ADJrVt2/FEXD
c5eHkmnIqElc/WgJSXqyNHqbKF9PyFYuTlH8MaDLgFKC1cP/DS5Pm7T3NfCxIThY8Yi/1d1sCdFB
KQokiEvBpiEvNkUEk4OcelyS4fzo2caEY7mV0I5B2h8dejBqkKhTmH8251Oo47CM/2Ikn/lTptWY
3HKJueiLkk4Lwh+Qe6d+xZL+Gy8ScLm4+FA2uY5jmref3O/2uYoRCMA5vR6uDmvZOwYKxAjw0CQL
AAfEvDN2ECZ6/faYJquT/DtqEP6xGW3TgpDTgS8AifcD388n2kxOid6N+FnVIvEz+BePkm/U/QGW
2Eq+Il/S9DOUIybd5rn7Y2go/bKn/B327b4MlbNFQ2d35DX2Otn/DfF7nWXTPOGH3GDo0cfzIeE9
b0Zi34OAZ0LtxpPOop4QVZAi0/LZolQ2Dq62eMtQDPI8AVZ/PyekaZx4A6DWeqxHTVWyPbRp6mbR
mX4QJjviixgm0f0DP3aZ6PpwqH9XrWYn3TcceWeldV7B0UCLLpKyY/yr8YEZcYt8p1Yl+mPt0cl8
031TYGEI1csgwOBTgYI6QSkE0GG0avWkIgNtjWtCc9dXArzb019vOweJIMGisBN0VLSHcRO8HImS
5pSCDeGj0UoJdsuxAyuQtzQDXlND4MQ+xbFPDBNJuD+lI7VbpB5LyERwk7+VWU3lttv2KzJrAx5Y
QZMuL2t3jY34KeoDqbYpH4+NLnFURe+nCDOfQUYiJHUXPij6ttPKQ3uuEIktOej/aVVmpou4HdFY
R28gTR2JnaFIrBYBCyb3W4qVnK3mZgjxYeiZYCsQrISU1zZ2cYTWsaVPTXWb+Db3ZRf3hosnRtlE
aVI+Oe19LmISvGz/LkUfBRCF1YOV9W+e9YHwPpLnH77M7+VsaZZOECYeiowFeZyoqKKzdSXcHhkP
QyMLwWITbvXP4h13l5rXAK7/+s6vaF1kvSkBoc454XELfi55oJu10iTpKPxOBGB23t2moiKMuR+m
X4xirFqx7cVVbGLa2nJGihiPctXJxYgXl1Nk81NJ5+OYlZUYo3Ah4bu+tnWXZYIdPuSRDEJ15uPw
nukR/d1eE34bg0E73EVITgwZpd3JC4VUip65XJjAg+AsuE8e3d8afw15qSxnALITVBAO4SVGZco7
cQewMTv6A4LybIijhO+BI/wNOsj54QGQ9U2C9GjePmFwRUv65lAgzwzbxqGIXKntgd9kLO4+Yd34
/ufbb6hJoACx2cvDSGPu2HReFdBwV0JpjKPrrRo3f1i6s8O9czhBmujGySLYjXydlAG4HskM14gc
3KjWsVXQM613bwZl+I9xomhaku14+Lv2QIHcl9wyJE9yVDqG6ZNWqzuYlnHICRZS8DBH8i1J2IJp
ew8HLmnSixKSatDH/bRAhxEM5wPZY6XanEFcoJLYTlyG16+oAP+8IjLvZx9kJKkhubOFrUcBRsD1
mSxLL0F1CP3/pUD6wwnqPynrB2eXz7wgnZZBBdvCBoCHy5Wu8fLWmq9PNkaRDHUTq7Ob6TaJOZJy
dI+NBt01DqN7Crk/LMWOhW/fIuwBJID03LjpM0C+37AHm+t+CKiwi5McmwSRzAbKHmn2ay0jB1EP
7nu9PAvFSKfDrGdUexz77S9+IJIARRukpGmpqHOnrIz0omeFjCuvNQoyqsAnhOtX6jaXcerlGEVI
LW3vKy4/weB7KcvIgvW9c9oyTyuZqbtaFOP3NFnmT+eUvQJzDb5ws5nLwvbk8ILLcKgLDVhkDQ9a
N57rzTMGxZCVAIz7FZFtLKyvymeubAuHn7J0iX3wFfFjfUHzbwvb74lKXXLKPz3wOARs8a34pwm3
POL+ROz2r7kTYSndXyYNwyNo8nzG6YgKWoKOGNke17XVw4LFYpmaUQ8PMF5mBMiSqybnK1aG5EGH
ZuIYY/sNbBpRkS92hCOnZI3vuLDxS7/rKZTShNVoffmGSC8m/kjBMJhP3R8GzeQMqx3jAdWeDMnx
AtoqHY7YXHNPOWgZu/HqzJ/x0Hn8p4qG0GELaCyDeTEfn9GMJ0qpTedYfHVkt3dArQGpDNFcxLFG
kYEqHzuw5zHHoU8Ww9ZnGKCoCKCrAlgdy76aJvMzh8lHPj9JHkbyyQzJwh9ZKtr0UvVN0sMaLV0y
Iltx0I/Hb8FlQeNUzgEBtITryUn3J0lvkTQtDQK5jTz+J35J3mMsTCJrSW8y3e2BMpv9Xg5gKEtY
kOhVv73U7osVSgPZtAKz9NbqVHsD6JpGiUxL3K2RtAnVDgBVa1PjnkLhUSG2N/rlnoI25GobkaT3
vqpgXGCf8RKZI4yPSCDFp42kt4c50CnboAgGtM4WXdFI3MQtsVL/XfbR1ijSQtHkKgXkeXXkCaSh
dClO4pFxjPPvMLe+hnj+QfbIlKHYVwD9ZfHyuFs/cZK+9aqP/VitVGxsFzxCDb3rSRrCaQRuDwtH
iGZBbNTdpe6OmF4I6mdubNf1EZkOSbg27pk9GtE8uOGI/yQVeS4lADcxSjSfH9w0vAJgvuD8S97I
PVUGSwpjm8wQqcIG6KUu6l8PN8FooTBUfpEcN7f4fOKOLSxtEfifMbCWT+SMYA9Rb64OxbdfhyRJ
hTWWRuyVwUJj9LQzYjLDnckkEZm6ZYLeaTQVHhh0nt4i8e7Mxn69wK/wYyq9LDZS7jeNCev3b4iw
xrvYZuAlRfwjfv5qVPzKvsZyPRvC9YKn99eITmjIEkUZPFf3jDV9qlLIcaGwzfdFjt6CMsAlOCqc
SJ9V2BU4YuIjIUV06dI8HdC7pi2pSmHcbWSzrwj7AsW8dRBbMf981ir/7Vlk4KHI7bOrdQIPIQl6
b47qkT75MnIqkyge9V5qiFuyUqW2/4BJEhezsiojYvsDFFFFGhJGV+lfKBf3yTgtSNhpQIieZXLF
P3OqCpyAbMmqmFBj5EJu99Pehlsh7ss9vJNHN1CoUbC00JNouUYU3P+YKGh6muP/HZeoxjhzSlaX
p9Kc6Hse9exbBX2cD25x9RIX3dryGFyKPv0pqGSDgKJHlo9/VibEh9bR0Cqas8mgWOgyaE9ChTeg
U7Mbmr+IwMceP7D0L4wNGN2CT4OLSan+ulpy4bvwll0QRq5RU7AWEC68F9REVYa4en5iaQzJnUUn
hp/PXp8JgPwbpPOOUuJK5D98B2yW+F9YB8o11UDF2jUGDXFssGFjR4CGRLBP7psdzsuc02a8rNoN
KhYZo3SXAiAtivmbqHQhI2XCRr020YYlA7DuxT3J5br5SxUxr+J3RSk6BS13yDKJkKy+VVEP28HR
51vjr04wZu/q6Ti1pyhkAe5+OM5FPEiDdm1+ME4eXSOSsBvfn2JtmvcZmPuETSBv/xEIxmtsdyar
GZ59P5fJHV6zcx9lGTMtDqyAt17aFui1z2ZxtoDjIO5ExYcc+1NIiTNEanz2xHr3gPurej6FS4mO
qALwN1dsNx1p1vxLepD1mzfqXHDFkJr1hojeSsNUkYsURRCrOV5IUEl5fXwKPsOrrv2QTwVaWEVQ
L1ftuSgQOzZ4bG7hVdvFbhkw1hWJKBuyP6zLgnd1dw0w6PwJhlBBCURckI8MJe5gl7b8aeTvQaa/
O94F5EvdNMZHeB++YgfNzcFpU+UpNqKvGgxTpB9gJYN/tmShWuxFKGXEaHyOzCVsYU7RizH8J8ep
tlh1tz+Nd1iEvs6rJx2PgutOHiR6jlVQ/70QcXesfLYbiWrbuejSwL6kwe4ANdels1N/D+zh7zTk
vNepVXc9/bQCBsWhcEdsZxqZkpXnuqVY0k2DlbqhGIdscJ37i0QGQwvoXmxEo2dHBbn+GLMrrgcR
aHIlZSTNPqiVE3algb1FkAkGhlDPv/JqenNXCwEQvCdMoesJfbWAQKNhAdW6ZJgK5IZrB36MVBNN
CSo8Y7DydZTAVsxONijDBtnRijMVJ5R1Fv3KsjLhj7wbjeX/TWlC6VtZmnyC5mg9oQuuVzjB4oSb
xp/uth+3c9qBYmTqcQYZtlnVlejPaKvHcgEhsth6GcP8U/wML9bktoFnSmh8epxnVfXN01aLgv0/
Q6TFzdZujob3UQEQ/q4k6UZfUABacfY/n11cMGwc7Et1m0k5jYcPXlF9R5lsVZQWwp8E4BE9Hd04
oZlgM+EuxpKw/MAeOD11HDKilbp9LNban9H8LRBxDAhsD9FIx7Yyl/l0bavGg8kh7ZHR8ohyyY80
f9PBYFnD7vwduwwSt/I/wU+EnJNAoCr1f/2Vcvcf7idiiZBzKWpSQ4jjLRl6/qBVrMpU0yPdEUcx
9Lsenl2JRt/zP3mxRLt01VpSS0TVGTV8AS0jW3i814KuVLvIS2PNWm871SMJC8zaQWQwZ0B7WsBV
7FiUVXRMttnzlq7KAjf3Gv3DeSfToQJzD7/yTn2rwYSlW2bOsob0cAOccW+kt1cyctMeugwXHNci
bIjc9wpBU9/eVs2hLkt6K6a8rEQl+8pQYHRAWC4gdcbL5BGUMx0RKk1nZMKl9RpgD9cSbVuBJqoZ
exhUCq1f7JUosuX+ZCuuOV+b0aWp7BJPwD3TJgWJVjI4Q5q4CLcoi09k2zAKw0W5srRqA7QcQA6U
otwfXOZUQ8RBtrkXZbIU923Iqm/NbRyGFwpud34YXaxQ0vIE/wnezeI1AmnTcz3NULJETWOZ+W8C
0b8wTsXcfeSfCJuu8UHMFnkpZP/sW5RmjqZrgtXo4TKkYt6w3/JcEfAoQNmS8BiZFMyeRce8QFiJ
ddGiH5VwTqizffR+x6bsWda1w8ep/RUXpbTNYfP7WxlIr4x/XOxULsPwrezXFz2Xrf+yi2+RAHH0
1FfjCzc8WoVBcBqsjAxrwM9IL/S+QKNqOHWUK/KdgJlEQ5N+0GUfs3SXQ9vxu/Tg07U9PhC7eJEI
JxKeyHBMUHnGU5tuy/wEFdPP5hzbb/cJNsMdN37iY/qtoxqKr0rpwq+NO7LXeCwAOT5e1Rmi3VFv
tVSGhXXtCyj9RxVqNp2+IUuTk80rM6H0ufH+x2knALwtdikwaKy4NwijlFzm8GBUjYt16uxAM0E4
c7FmsbIH3f5K7C7CwfwZ9FsSMB/+4HyowpomO/c0u+/ENgSiRXg9tF0aYC58MrMOIETY2l3Qfesk
vwOzaqIISDJ16QYOnEVZk8yemFN4ruLk5+CKL4fi1RY7qxjr408w1Z5MqlDQrcBlUcBwzg9xY59L
c19h8nLG6NAJhMoy57JC/ELHMihd6rcB4jct/JvBCJ92UwlPLNDGA33yRMkbWlatoK2dMz0+5F9G
SMonfjkU/AUDYBOGxImv8iuBsT+GdWLp+D8b5eLBsFJKesY/uttycbZGRDbHFTII/lxu8NL2hv8F
KarQYu5JkswfNIB9uWLgs+qQli4bMKhrO0yeEg2uCtOdGe2aT7WNaVXDM1FQlR0olqRuDb7926Ld
4u9/mJdKltr4nWna5uvBTaD9avNpNDwv0HBjDuFe/ucY/GBLZXMtq0cSKf8wxTlZZWzDWuaxPBBg
xKjfX4yObr2Z/hU4+xVy3XwsyODqyvEYKdKXWggXKz/8YMiT8wLpDCnGnCHN+X6urNY6Vmj0SXT5
OHdY7s0ZtYD+xuSLcauVknVWO68UWXuy/vmVnaw2XqHloqTtiD6Ui1ptDQuRBoIpAPSpQMXYio3E
/nskQoWOp0WsPErcjnHUnF6J39XJR2tNipD+gwmv41gIebZWgJKCe6Htx4xm/AjkD9e8RxKo0nYF
2P/Vo5aqdrLlF8QePOPLvxx5FZurj9Y6r0gqqSZcJWA7MvG2T5xFxJQJ/S/NVKYeBjJ4euX7onhn
1/UQ007qERNasWUa0jpRarYb5BKpO9DARqPuO7wpUyY4PtZglQqiLJ2th0DtgXrlpaKPOfJHZ5kZ
XNGQVTtyEyLCoi9rfWlJ3twQRFpY2W55QESRzr7mS0l3OWjedIhXwGMGToljVrKr9D69MfwI8X5k
Km6gU88begQry9GIntw75ppwNZOxUcHIsjvVWvkgdbboo5TMwWZPKfxcJQhzQlwrgRbffge60gR7
misajxYtZZZKQ9+esA4Q8eQ+FPzyid9fyEaStSV1r6LsPbhjWqkYt09e6nMuqn9gD8pS+hlEkpwX
Fl/uBq2Ipmm9F/aKaZ9VhI6lO1ursCDu1ueSEvbl9UM3bhlXWvNu6Lcl8JXrbFEBTwUu0olQRviF
9RKGmmrIco0wuYal32Rzkn+TtnSqbczt6V8QVERBxKuRiSlIX7/KoVTg55UEHnmdBKgg6i1G2cGX
w+7kUY0ZBy2Oxl3quL5NFmAjZyor6cR1EEFqO4MB9J1udVMdpuiFGMto+QeDTViSCkPn/mok+WT6
MBHoYVWICVKWZGVnGSVEFekGw/wwoW2hPHsbI+4y6d/9XWxU16DPVRy1ckJrLJeCSqUKxkiMPzVi
qnr23NS7me5XdYb/CX8PRXggMmkb16RsboZ0pQ54yITur0nd5oOwJOb/T/BjtAwNhWRd3ASloahi
S5Y09EDzrYrfxsdBSGLONBfZnJ/hV12ZF85IdMxolLQA76CMYRe1fTn883Sow2utnRvFO1v3idFe
OQAUQ56QcjMXtHugJ/rjXVv+U5VlDUNIgr5rRqkizgVVtvZpzP37WtLy0nr/+BlcMtaNa7HDWLpJ
E1D1PV5BUX0ZCyRY89WAa/x7SkZfiRhERC4D54lHo8pUTWjaUC7tK61LcXZpJGGQytsRJjEx6L8d
yNS7iovPgBQDfnpPOWMhCOsLtCMxQFp8+7ccfmORDuY+4l4jOmtYVwPQ5+0PUaDS9CNQ8sPRI5RX
gXI7g08P/UEGDwmWGw/dH8lYNbBDM7nrur1nVpeC/dYIjxdY3pkaacrI1jTgnRRlX5+TMN0LYJVT
E5V2DyTx0L1qBUOhkBCB9tdo+510DDkgFfnKW2YFIa2Ug9QN3i5SdoZF2wRiNTNf/t9vlnFYXcAE
4ItclxlMmP9LkaiEs7Kpuc+/T+aD91CQYZiLwXk2CJw1AF1NUPvJkU6ycqLU6Ckz8C32WS3e9NR/
loNJVkfzUzghQ5p+tiAtln1H1N75vfAO7i02AFaksNpAkMUXOxNlwDJStgUSyOO8RuG/x5uMbHrx
7nX4IRs/Wb3lZuO5dLFPSB0RNZbeGjvyY+5dT7IowJFwDPGrU22G4NYZGEuTt4kmnWnhq3RogtYz
cgkEygIkz8ZT9XIewAlWMKPlyuN3npjBoV4JgL17/ONcokejYkWK2Svxgt6rLfcn/KvGZfT0RSQK
2P7t74NaothP3KLIidIysdTeCur9fFxE3NAgvurYgFHqo91QG/g7xDingAIORxl+SGaHHTAmg0eT
hntQBBEzrIjCQzvgxayfRi91z+3DT6NVzUNs3OTxREbQVrVzgWR3b7rwX7vuX+kfz6lIahWQgj9v
/s/Wh/i/Nu2Xscb8f2bdfiJbh0dvwnYdYUVIeIHilU8fQV18Kvn2Ve99UhxWLCBJa/5BMtKie2w7
0AbWRHpky7w8tiqV3PnLYUgdGguaxJ3MjTQ4ow5a2XHnTWdFVvrAx8ODZmjhOmOyGBArzmpgJDQ6
/s5FQkihOJLudaLJgQC0SIpYJS1KsP9MlGrBWRtBhZg0AtOFVrdCVfX7bZOrNqnCAW2BeJlyLTvd
dQCwwsvW9/9FY328u9cdULrZBOulGxgf04YgqEdi87MeI2b3guCiitbiWYA7KsV38tGbeeIGk6ll
TZ37Iqc6NLPv+w3lfA+PxeQmUTekEm4R+oBTCdHNZPVtQl7AT2wSOaBuAyPKOxlvKk2CUDZ2sPmM
5r610jgOg94wzqzfjYWdNafzShdRiwwNWKx67b6C+JwL7YcOONIfukGzdCb92BstJ80FWEXUaBHq
QzfNG+Fx05p2dEglCblvndGdUYJetY7f8jCYoW5te3GJvyibItdoYOyBIcNBwMv1ISQO2DjRe0yh
XZFVjec+5zw5YA1GZedj7eCaJ5OpxrmHHmF5sqZBaqLy82AXxHRVlLToRWCEVmhP09810m5iboQG
9GSQM6du3YiOusLK5G55S7dUF+4rTpkIQAKoU6IvmtNKM7YNJ3v0WipE5k0xA1sx3jO2s30ayW2/
FT8n8llWKQYJS80JQndgRoptuxpn19YKt7/y5XS+888peKFRt8ueE7O961qGW4pvNyBiYGpEgsX3
/seBYuyB+3fTomEAldWn5Z4UZ2L0VhxqhMIEnlYExPn3iCCCHQ+LjjeFMGk7BQWfjylSFn5EWjG3
StpZSBb/QzkDAd60sE2Id2J10ZT8K6V3MH/1KBeS+r4iXT2/WxAr04bfbT2ZU45/GHNYKJTFCtBE
EXdR8aYpQEyTY+jt0hoNMjhvLwKqL4Zl95p1P+bfdSFBoWhPSm96s5tq1Dki/fkqmB0vL6tpZgZf
HnT6drFR0giT1X9gVRuxtx5llEc3Ey9/f9JcB3H1Sts6G9mFhtcRvTvNs5hGIRMlzn7hG3ZeqiXn
PzcTeEvDCcCC3oWFekwUHIdl1Cl8S5n40ZTYDaaXselnyOH4wdThJn155yN6oel51E2W7tEnKgX1
KHQaz5iwHcJqpL71sl/iF95jFEFRmJz5Ijy4amoLh4K2lpKOYeCSyLUs4YdqCe+V4q7pCIIQJM5E
kVjI6wRierW1tksAnM8VMuYvjBv/Kw6UglJS7SD2+uJUrwI4g6JWYjmwnXKJrFsAu6rsH/CdtcE4
tzUkUFxb8bMdxPF5McLola2W96Smg9cUvlnPmDS+fZf6kTOcHecCJf8wH7cuz0DebmYLF/F1p285
JOV39uP1xOnRSaeSmlVIfEQx5Rmt2kB73mdMc9WYtUYXbAlgWFGx3Wj5JwixRoXTnVgHaci+vWh/
Im4KbUNAWRSDki59ZENmm7Dw5lFRpqcOjRGGdeRhvilyN0V8BnHsI4fRCjvAndHzQYwWwHHkI0ER
8gz/kXEw0MEdgvLygUIZYFdSyXLe1zE4s5wtgAZlgZxzx9gTI7Wz8wN+RaaF8R/4rsw7xC9TWRZR
hjVcwE1Yozns46DYG56Jyu1S/e73LA4OaUyJ3uI55e8eO4B7kcWF8Cmb4eAO1a9DiN53F6JFXrqo
Rs/RyFoeMywzPyYsn6LlAd6V0Ayu2elzSmZz3omL2nkusYkkc53SsgnYZB1gSqxyPWakAZjvt38Y
31Tzp3ZEO6tOhhClXoHxLY+PZdFeK57VN3z7mAp/s8/tV+U2zGWzjIyOtXhBM/DvMvfKf4kPSn39
S5Svt167Pcldx66qFlD618F8BU5WUxBmFKDHYg70U5//xMJzTyd2zVy5fxK09gV54P9BnowUN/7O
UUoPH/BJLlVNLIH+29nkVtWMiiadQslNjAIFtY5usNBSlJ7Y+F4B3Sqw++UkbRPBcf1pTBE/NtDi
9P4KfiWZfjSAWXaQEx3F0K8BnFg31i1xjuVhFwWiHexXmtpxqsf017/epO90T1xaTi03UJqVjqUm
ro/KZGTd6RS2zHhJO5zRymUkGwtKaw5wuqui2KYVeTFPnasRa7IWveidFIlGMJrjX/uFY2TvNKQe
fWxldvuN1MjmkO+BpMv5sBTJYkHpwMF3UUet3UxbSLCMt2YehLh7fxODzIJnO0YySxDNuS+BFVAm
fPZ7AZPfdJcRvL7qdq2V4muZHUi6s8OnHqf8bCOLDrBVL5RDogsY0FQt27vpZLipqSaRxsKLcHQB
RyYCl9DonQov6MyTGUsmV3zkBmWzFudp64cu2GS171rIWdgepgj3r7BeetbeEpx8zHyBj8x8G/fM
N5Dld/kQBsTlj3Ph787VO/FXT+i8GJCk7AHy1mleCcVI7i76sp9IJiXudHw0+iWfKEYtdG7rlgu+
3AlInWJYwlMpHTKlzhkwUucpx3tWnWZPDLtNR9+yeTAubdlvrGiIiDiWhIFZZ8aRBdGgWmkeaqD1
BBU15gQjUwww60EX8VwdwVBcyYAC+qekZisSse5ZbRl9gX3izywhwg+54mRsNlRxqHRX14qmWjSR
w/Pi2f309BWr2NwJ2/FPUXdUsMcbO0yGft5D3e1oUBJg5EmZ19XjPJi/j1sb3lufdQE1uy6rsguf
lQ8jvQJa0IlWPeum7fzO/zmICpurAWQsH8x4ftvHHONID8jt9EgtBvDS/oAnuJuzLkFbBFGpsx5+
OqnOfK5Yw2TYId8zv+hYLfhMTlWRnGuRCxrgB55bzNZzEcCZrq1oDpBGcd4mZYfS/uFrNGpcGlAb
SSvsIVfrJ0yWmsrpXQ1HARWHKFNoqoIiljkgNgoQyqUH/gm7+v0lJ6+5l1IrscsiF5mp+syJUVgT
d3P7tP+GUtGP1dOrU/qImGORhA6NxQ05rJ2nONlf6YQapOSKq5RZuVzBAaoUR1Lu0tA0uLtwd0Yr
6MpYrPnCmEaPBrA/rFpgx3uRWoH6hJANMVsTegyndG7WMbHuljRWafDH/NVsHnA6pkB/rNC1dm3n
Y0zyKOqvw8mZXZamUJRmm0kEeR0zFN/2Mhja4lrIGjGg4BfokQP71+aZJPH8KfRcGa1iGQzGqFZT
MamDiq17XwxJR+7NRFK5wiZx7zhTSXroaTi+nu9VlKNVap4omQJcBeejdPG/t4hdS8jlAcUOu2cE
5qUsUD9EwxT1YWtu8p5jEQSa7BtTa429Xi+11yiFBencwIJqhtT4iFwkxSs7w1QpO/J+igYU79M6
khITJF59cVfRI+UNSwU3DvOBXNezPBgLsgVOyiJPtP45BT5DCrQP76VK3FIQS/kbFTKxQw5Oguai
8I/sonSm1t7KsBL9rjg+yjzKN8p01d3yP5bhKlvEjAQh0utpfcOSQoRyr1e363SCsdtO97syt4Du
xhjdi5NWkcFjCyFUqURcExDtDyYnQv8vST6N8PWXN+g061Pk7gDKj0fZpPWJEwbo5FIjQ75SW5ym
ihd7Tw+vJs4n6o5LWonp96T9fBLFZ/sM2dchJ8Mf64urJpCFAM1jab/oGogAI0O+pCN52Wibf6qv
BKrsEYprol+yTlVhjA81SpI91XBh9pNrfKpThecAI0ldKyNVSbws1AAWq5BPcaOpOHFtK+R447za
RFxcJSbkQvcAq/S3dmlV4y38hwkIb8AW2eHok0KKwHGyPnMr8916GyNKprS+A+WHCV+Sg71RjVLG
SAXrhHBCNmWxc3sheAb5bnwvVLGmJ2GXamYSMaL0JWJfrJHePFeyuBW0k/kUAH+lf+D9FcNi2VMg
NZ7LwprsuKFnd8tZgzEkk0eN4BUJmxr078X2imBp3m+vNRVJ0alMKHxKVw4ky44IeM8LKvzKTiZq
TV8kHr69pKxdJ16h5hLSOvGIv8s7BCPAffHtHkQ+kz/SieyRb63WBNKQ6el/A2MwHLHqghmRfaKO
t8JSZV88zHPzRTiIkK4efRN41xL/9ljOinoDcoEZJYv46kp/JcXsrrMiQlUn7486JSXmK0b+7XoQ
WDwvxpj9STuzu7lpDk5XhtNWFjF5KIiTk8HvFfYe5qvI+rIYyzFKNbB40mS0Gw5aDp4/r4EMb2bP
rKxqdjVKn8cfPmA4100mpVAcXjXKJYEci85RLveDTaaw7NRaknQ49+xyiso6TASRLC6Czamr2dkS
gqdojZqU6bG4mfeZM3sq8f9qPF68OsmA0rFTf5Lhvx5tkkJDEkMsRzplcO2BcE+WvyUQPmw3TSR/
KKLOOolTOuyU4/Kh258Sutc9DBu5L3DXi1klkecoc/mrYUZH3tCYwqvRwBcSn7cGsa7BCY9KuyhT
oSnxPqcpjtGhktJuQ7MFWADMel7yoALxJBCGM92/gvj+eN3ukKwvV1t9tgvpKR4if3YS4OM35lm7
Yr07hh6UM44Xiw4LkYlKjFE5eCpbR08Ulmb7IuAAaAey1gNhEmsnzibzokB1HT9yGWDPT9Lezuj1
fo1adl/qAXYbgYNFBK0I2YbxRLR/0RvEZDgHmPhbeGCflVhRBN2pT5tUGfHQtslD3TKb2x7VHcgT
MCryTAnlbxEovBGDOKzwyWvWQcBvjN+MhykO9kTR++PQDFBN3KCgU6xKGLD1kFk+vmh2TkzaSEjq
Lzh3e2S2ChrUCAdyALbzCpHFeKEdw++F1ahuSA1O6ey3W94eO1PZ2nv2is2EO/SRhMy8YostpkEC
79AxH4Qo0VkRKieADGWrySSNrWeNFSoq16hXz5Lqn9xFxfv+xXEPfEFXI1zn5QSO4/c+VUKNVVJ9
672ViQq2sYaHli53yUiAKVDR6EoQYopeJl/Ha5qmeGGwToeTUfqMRRtv3mm5F4/Y1cA+KQ3KIRBy
4U8YTAA6FjAPUAhrexWQqWbTJA3ETmInhaDS1co8GmvTHdG2P7fpV6US6wjmYdgC6BqIJXfqlF/O
SVoKnhoA4vNs9K+UOiiEwDWIhi2Nu+9l12InLjNO6luA7bdy/0hL8h8dhGqAo6+dwhg1ya0OmDUX
bNSzGiH/Des1P/QkbD6/zpXvPcC3ryLnroKowDafEKT60VL7mixeBd3ERjy2GCpv3xQ5xrDqwb2I
QT417LsCCY3FMfp+obuGeMTg/+gr1pc+XaSvjaIn4q1qh4MmWlUlg83/W15oIeXNZW0QqkSVFn+L
CMebR8EmX8bhp+FU5SI7QEbI2Bwa1hoHAXVFhFuyIY+uJXDvHVyLV41Jyo96qLRn8ccuDUTPXcqa
XAh244ShHj/0fhyiZD3HT/tRoeqCi87mTcmI2trxqB+38RJYySJBjTGshLLFSyVzAu5lWQUcbVPk
lIoy/xMRacDGgL9g5kXuqB9MWuXMrYTrRkYJ79iA866T+phkIiqvl7OXNkZJR4T3AECXpUinYh9a
xr1ZlKtMXFanpplcnNV21UeAsBKD4I6VjyeKZwmALQjYiZ2F2jiSvpudnwW7xNYhB7oGI0HeuLb1
aiggxYjK9PCcRGcp+lB1iJwB46FNxCxjuFBjNkoEegpgfQId1Wdj2ChEqTuFTfGv8Oe98csFkOgF
QYMVP0zSbCMQPOjaYuyV6F6X1cLLtpquvATo4S/31tE5oq0mqcZJzL7N4hEKxT8VSVM9mRVCPv7s
+Nqbum1jDisspWjueQyzo9IM9/oA1bCXK6i7VGGSK3hoL+n0HVLzohj7Zum7v/dIlfyg7nf3aObL
H1mObdXcoTdgZdv9mksHTtphYpPxZlUUujBwO/PjzGCPJEyWOPuo9n0vyTBvjqKZAlj7ikfnm5eS
b5DEAjjxhCIWXVu+quxapRa/7J85UH5QK+GWwQwz3ohuWlug63r7sHSUaANzUtRvPQp1cZZGwV5M
/1gzZ1MjBlznyPnfEF/PkReacUQX6Iwj/74gRKtMbZuNfC0RSfnJKCL80Bw8GnzEoH7Vudq/nZM8
0FUhtsjYPDwG1k+Gnx3dmIvH+lmPQPLXv5bQDUQxXohuRwmWgNsEsAokXN0v+Dhf7MedDPTTbK3E
N5dH5A5jun0u0ayRoT5abD9dzZF7000t246+Ms0ax8HTKdG/vcGjfMQy+1y1Tpom3C8on/NICZg9
EaIP17SgnRWTztHKss/ofs3EO07Bxh+EMBbAXRo3eXBTRM4s0B1O8rUke0nlbvo+QKNHQ3hrtw8o
4eyxqlNIvgfvrHpn4QphHlpUtAwYCqeuuSS/2+Ze2s8HCsg/HrvkIWT2obsriA3mOQcnekd+dDFf
NBBa14+M1+CH7Xp9CT+AoOuohbF2+YklMuRVqMvRDsEj9TE+VX6d4n3ETPnSv1oMDxaOByG5e8Bf
hxcxf+pdg6h/ApDPJZZMjh23m/2slYqENUNuqkxYLVQZd46uEYx/v+z7+41tPZ5xbbLff+EA3VnG
SX4rSnB8qZlRAowk0xpO49hhjwFLH07cbB4l6YqtrpiLmVvdR33K9vLYySmyFWSHrZV8UmR468NM
quRYa4UBH3kkf/sGbAtAa1gw4j8g/adqhAFjEhvec73ORkDO2df33yckzfYlZm/pe0agD2fWqARH
l9JbrmIHhkpk8NjN/PoGo/obMxWFMhB0NcEZGBKLEzpj4iqZPAq7rQtN5O3qOQ2iTM/E5fwEHG9B
gNFtso1dlnQPZc1uH5VjBRYuqHxkgnp9ui7s5ucYV73SUvkQOaxUfPr9Xj9gT3oIRvfhEuPeWH7Q
sDdn7/WEfM2jdMUCHxNphnhOAKC42nNYj6xdRlV65JpIKicsVOfwzAdIR2NI1iwTYOTRZX2lQBB6
+HypOmUO4cGAtlmxE4fA1eWNrFXaKl8jQhTrKQRZqEmWawTGWNKCzOt0jvSLK5aTQOHBrSy2X1Gs
D9vyGFgIVwHwVP22npb99t+nU/auBrgCUt8D6DdMcq5/IBItPrF18PHJvvnvOg8fnTu8zWW28Hoh
R7g8k15Df/vUdne8yALP13KNnIDEvC3TWLMjcCj7Y/loL62qzfqi+Wmjt0EybtgOBT54zROTIIdU
uoGL/X2DMI8laI3XyDe0JC+NLngwXKTtCSjuqN3iXCV1/Gf1TzJiGGyRKI0tYrhaIJ2QpWkXtbGR
ZjcqmLAKDf4w360Y0ASu+KE8RxK/1bcXmzWwSZCELr2sLLRE+aWE20zM5P0LmRQRjGqnRaxyHGvu
+5R8LrsnrMhHg9MpB8CCgh8iegVyFaU4aNZz/VnHKXnJpUlTC5awNX6FgMFgGZCfReFj0E6GdsrS
Rt4V1eKYBIa8Bb/bA+EjGFx954qb2kMxb61fy5PQw/wWUZCxIdB1IRaj/ko5RYHNgVCePuLgEgpO
n5KhUM6AQ5wogfrbsj+EWsZOyXktcAcZL63YMINYwskn7Gyqgf7C550dWI6Uf7BtBB7LmadLLaVb
f7mM0gXKir2tOEtoZz4cMcu5nCsdth07yrVRYn8+x8BrKm44yB5H+aX8CDLP+9k98LJQ+DwQTMGT
Fcuh5N7nnQ/T/JmI8LSkeDdm6alPdWwHRybvZtnuRC5z64UFxipnAatVj1Gct8o5iPUb28DFDMO7
suu0PeKmaBpMWqJjINL122eeGY3/1gD/ondVvIGmAC2xjXY9KhcuRCmsWz714sDE85MF7qjIRhPw
EN/1Oyszh2uoIZsXrLFe0k409jp2BGrMkELOsFaCGDXmUtugRqP8Gle/PM77ubH41UG50PnPs1/e
fWS7rC5FKM3bAJcAUbBEkZiwqlzVOlm1314roksqPE/KZikSPtumbcDwtafmvCRMcwRLAsJjf9gO
tGHUV5gJD6ep3UDrfHBR0v9ZYWNnxxaMPZ0KSCdNdw2i7EDQdnfs1JAakT5j8cN1opiWkHyz+AYY
gqgptRseHFbeU2g5aRMO1eXKpJSa8SEhLxSlq54QUmpB5IGiNTNr5QnlklnjYUSIGeG5jYnMos12
RYSaugcND6obaAKyLEcqXjwJ3nACRGr7XYFKLqkdlx9RBWkRxpqVLgdxZYVi5BqBQUjznil1Htjc
xHuHDdxIjTu3RcuN6iqQT/69Pyg3qyL6guWKZ1onbdsIIM3ljY92x0yI087iuxlceRzAwNLH40aH
QnEp3bZD3FvaUX60qnRn1UtNUussnN86ygZlbM3km7SgLIfzjwnyuDM1RutCukGaHp1zYF/ep1P8
rsHfkDT03T219hmjsecczEmmHS5wS4r3VGjsGWjl9iSsZTlmuuF8+YvxoI/44kQtkOsWbShWsdDA
4Uk/9wjGkGkYPY7S6n6HE5UytEBopYuQHpfwFdvPmaz0V/9fe6hhZjaKb+Qzj0wAcflNruc/SjHj
PbMBu/Ri9gosi8kSDmXoblk7saFThjdOG/WzvT5jenOzE/Ta08S0+mRs++sL2KCZjiXX2Q84ij9A
EZUjdyjgs8hxjH++WC3oM+QQSZnIKAQORXPG7GKI8uWXl0UA0yo3USXbU4F6MiFYy0wC/ftnVdcP
TFSHhK2MHasid5Eo7kQuOoD2LFd4AIgwuv5KN5OhjIF/ISEGqmEyM+XNgohhgojMfuV5WEKC/Azq
ZOdiWLI/sRceSwKhdLcPFTcQso+DCXj5D/sX5WTzPy3ra4sH8XzwzjcDZXsBCkumJgF9qTREyY+s
9Qiu/ixNm00jhCRl5gRti1OZM9XS5AwKePvVrP1tFkxv7xe4fdp1eGFCPuyPnokdoM8aqqy2M4yo
tkpDf4JQbOmObr6XOd0RezFdsBZbwvZdDGgGvhFve8DXMJyb4ow03Wjbaagwgfee7Jerk1B2A1cr
e4RE2xahfOlm+s1o794/oobBsnDg24RcjF6gQ6YoOZ6Oq5xI1gnsPT+EdPN6ASbaJiyGw6Bv74wA
5y4yIr8fdVVOuQ+A0uB+zxTdrT8GyZcjAWhVMKbCL0qXXt1YXQNMXdOqbC4H2gpn+fgsLygqrBEa
88fEBbUbHwYx7F2TFV2rm6zod3iXGOuV018J+giRt05NHB0CKLuqJWdwmYG9b7mkxVlieiNlsr5G
mp72hsRpt3QzmOlmfXZrzEribEz/oeZlc/GDmYF1XdC4UFkqDCkTOFEZsGQFK7QlLc5w8uOGUNCB
AN+4ILqUT9/NA0lxWB+OfIfABIGMkderLHnzMiCwvWGd3wqnOdWe483Udu4qxZgUX3GJ5+MmGiFV
/NCWh4Iw8OqgaX+vvRBODPeYzdZG0RWTs4tH+XH6Nu0f+WM0PUM+xaeIUoajjfMagG7n0JoZiNhj
35mtB+ilAcJgjnYQNsqebTHLAcdJBV9BnFsl9u5hfmQNQL100tHXtJcEBbbSSnE8Q+R/saZ51TPn
GwMnaA6FoTgyFewkT5bJUZ2Qg5by3i4gKZDMv1Hx10gs+DI0Pd1apJa3Ui7PpV/pr7VrjMeDy84+
zEhuPwz9K/jZ52HOpZ7i7Y3ZCLkeAe8QTSEv2x2Z5Wx6O1NQavarg+oi9XDMhCjgxPEsiG2UPjKs
QrVy726WCoMy4x98IWF/54luUM9AUxQFRS3GyOQXyChu5JFhgxtnpcDSB/vVmPoN1nXaQTknU0Mw
SB0o42w71zvbqsLTF3u6o5GEN7Jquu9bq/njf2ZrKT1ayqeBzDhMl+CFz3FNbngVRgNzpjcCkl7b
hhLB+jxNeJ9Z7jvIQ4lq+/jbABe9xfc0l7d151sy5upiqfFl4mUjCwrVMzLcaZmE3fhF2O6equ3F
AhtqWxpQjqV58TmAPRuCiOG2sWB9eT1rDAyjFHpmRzfcg8mUzC0uS35AtiFbkMo4pd/G3zr5KVJf
W0uy/U3i7hMZmCfhc5ezh9kx94J81wN/1AD6ojrIo3dixy+tkHv3C54CdbcziyYm+SBerJPOi+dj
RKq4sXHoWglpQ1Jk+xuwzMYo8KEzy3keVDBJ+6LLBDADuGcNp3vrK1hXqmzF7qJAzy6C2YE+1A4S
oB9K6ET+TEXn05sPz4JcVf4BJUo7uisZcZuTtTjuUHjGygCKzIGruHGy0ZYRcFmykpigq6wQeyne
4+8QiJF4k26GpN459B/3aVnh6N+iCQjw+1XvF7yUL9TgnTlTn50WE1ElINWlte46l05ZY2MLeEZ0
UcbCu09oIJ7SmVeD77RFr5SH14q2+8sOIwaROUYew+blNO/MIPfzhQ1zyQy5QY8mCqrYtSxB4X8r
NqAY5SL3H++08KBte1WQ1OYb4P5+X3YiisNVWOTgIZjOwOVfjNFQ2UZLuQVK7deagwWFtKSDWVY1
k11UyvcTfARlGE1p/Lz90uKhdjtq1J5i/v/+KbmtPwY7b91PK2APXpfhojVWr99Yr2dJAiOXyCTv
M8JEXN3AByrPYKjTz/eyF6sMYADy7c2mEIc4ccE/0GPHdqfnsbkY27E5czNCCh47qJCAnZSCbjt+
4Kq0xzBKbq5gg2wcimmTZIeaREGs4buioIpu+jM3s3sSKBAZOEXHXRib5CFoj8N1o1sBKQ3VUgzg
oH830vntqfRRzvRQR+8hG7xV1OISKvOD7N0D3DanXMvwThUVZotO9YHx9tdI+zaKoQM8xP8pd2x6
0EV+QI5HzD9egQxa7Z7YD46knTjt9uBFZc+rRHZouTQIVAMKH9Z0xtoqHQvppJ5R5ujdsCmw76t0
+EfcfD1pfAbtRlJQY5+nbZjPIhePd8Imebe8mgXRj83AfE/DM9E+38KePk2ZHJ0gPH3GCiVuDrXp
/flm9SkXXV1uYUK0gNWsdVRdncr9tvRUSfrtJdhUA23yn5kB7wFjyRAdQco8ZpPaY9BRIpFH1ElH
9SlpiLXMu1HPYq8Y+WB0JwHMOhQCR9baFoBqKtEchfSdIoL3cCbx0iLj25do677beVJIHAAcqAkT
BVEbBg7DqSkYvueMrA0At7jXX0H/tgusXPTlSnW3Wts9E5oj1PlKxFyCo3SXPHCnclbdd1vK6WHD
QtKkAEB+ASfHbiVdT+S4A5UU8laLkpWSk1AeSGTL1bRSAMap+9wSjnbrqVix0rmYMRKvVotgpFBq
dboEzIF34gNKqZiIpUAPuT/hpfmxkQJvTEwMo4bwEvUs6Gs81/LNDZds2MWg/plrTWAooKAFmYSo
RbUHzJg/UEbs9G9s9A7HSv9Mzsrp3WVPv2T+AaVFbTuNLVPo2e7ktXrEXonF+dQTNvqbQaWOfH5K
hvBgb0jJXTR9ZqPjgPB4zeEsAcKcp5qHKUTKTBPBTUzqIp2CLE/2CvJUyiS6Aaj3IF87594z00oF
RxXG8i+EYgH14bVsqCnKixEbgJVy5WQpmnRN6BkGHqBWeQTr3ImpT93nq0AD32cCv1YEhHlXk/c1
wrXkebrsAIQcdxSzSORc8CSooi9Txbpl2+ed4YesnM01Sx8Gi0nKUxFtDwpjjMYPx3CbNUL5pzpS
Bin5/SYSdoTeVSngRk4QqpEgSU0r4yaZtxbrmO88/V9cuEPEcWb51dNON7hSbnFyxEwk89K8doyS
dxeKIEYgmMS8b/G8d5h/Er99opnnrVORG45xHsbl0Ks1KbPJQr4q0zHt7o1i6uciZO2GLi2kvjAw
973dj2CvSrgDUoufBtQzmqx1vvv0lU1dfhR295lr/QPdUewV7lC2NIjjQLbqrjoXjZCaorbSEY7H
CqJe4FQPt27qE5Hl76ZltBtzbmk17xiSw93wytSvtEq8ZP9LDkNJASRNORWJqsvNFklo1gJgXUvc
rttl04YfdKYyXAHRCit3dEQlu9qltZn7s4uPaxlQ+vTECoe6gYHVb9wOygod7HzfOQNsbdFdpXhb
FngK/AvUZVvlTa3TY5u9Elg19Gc+vkRKPkcRM1RsbVBQxK5bqO/Fm3zDA8nppsfl81xIQHDNMe5u
uPN64GClSE7gkkX2S4mJlHKCppg++w4O6Ft/mhx2qAvdtVsSUlrx/xlxiNOwkVt8QZb+WoGMvRHI
8oaMCoc6c0HmChf2E8n/ZlzOxXNBkEg5xKM9BnSRZLhFQNE+vB1nDymKNLWVXZb3PUzktOdB0HhY
MMcdYQE1YiD4OJE19LpKi6JTsxKclo1h1cQk7QaRzxufA/jnlgDeyHZj2R3Q2UwSu3WtFnOsIPj5
dPFGfq5FxJpQKziSkP95dkDRXooXtcCnKp5RXRCuntbDqfF9F0QSUDfibJCIUs1vQCB/we5wJZq1
zdg+n2cHzKukcg0UzM9E5qlywLeAwbLAw5pyWouMbzy49NTotlUZJbq+nX+CZDZ42BelEw3wb9fv
FWJnEOGVWoSbO6L/ACoCrzJTI9QTIHJTtpPLQCvBl/yLSVUMuWP8T1UI/2SO+K5dtkiT8u0W41+I
vgnZTidlOiC3LrEn7CxR6PMoTBQXkSDfdBzEzNAEt/w0V5jf3ReM+f4t6E7/PZGEKQkCKDFoeNEi
oB31rCIFCh1e+iJ0H5FoOyLsz40t1zdON9uvDH/ZSUN7oJ+WJVUwDwPrpwgXIUpPyWsBqOlJjv0N
mXBhF7OOwvOVWGPZKc3V8YCUUHaLzj92nQSwAz4Lb+k0t4jAFXIkMStEkzZkxNwJawXymZyc/0ME
21hMGa3Lfe20VwmEHqu6/gQXwp9vqg9Or/fbtbNRr9AVTazfigF/Jgdh+DzGqy1jkvLLY1gpUg8b
taDvYuYaFpq9fm/9C0h/u2ThUGJd3Gokc2ydy4jyC+OSCiMb0kIp8t7ZtXWDgwtLJtsw2eneUCay
8HbI0KrjaOEmA399eZ9Z7ASnNOZyWZliIyxikdNs0fP3DAXCKNY1873uMW0AP5qlssXNkn3XfSvY
3Cez2ur3V5HC7haZqqH187y9eorO41ordC76xWnLRnTVOkflvHlQvL9tmMRnZvh5Fa5C8/qffSyf
Pj0Ntc3B95yms5a0wubv0aTKWrVfhBVNApLCDPfIjpq7wJt6yarWSYFrNZNIU/u86Fd40sSHle2Z
lcH/Aya1Q7HJa3onPKmAImJSqWgOubCibwz07XJZzStNVjDBTzHMZpjIxbsJN2dJ8/CSE9u4WBZJ
g/svqnH6uBD1pv7FpsH2Gk/9tRvwqxSYYq9kCY+deJyqbO8r94uveFWWDb6dKi+bEGMe+hXy/pB0
mXYo8wbGaZ67T8vXLkF1JBKUCViFLyl9ClwojZX0fs5fyZJh7e0ZBF616IJmN2R21LAj6dH7aEjz
sgDqKTM46tKf6G6RCXxI9l/5MLnxLUryuWbHSpljmI9tTnSuGq6qSWznZGjtOP9WQCpSrZgb3A+0
/lnLKwSd3ncBifP0AsdntzalVi9/z6H/5kZxbDwu5JSM5DPR1cRFXLYTtp+0wsSGRbSZDVRHZKCo
HVaKcLiXbg6JdIcFIGZMBb06xu5jpbpSln3u5AXNdNJ1mlmHvRGZ7NE42BChpDw/It3jM+C9MsqF
2HFqOFUWz0/U2ekrvW+YdnCo/VBhURy6RapCpnvFxdN7C5qamKMQI+IlA7sBkRCnGjROFECW8p8c
QqPgjAl1++DK44Z/UPyyDJ2Ge1zDb4jA9X5hm/df3Lbrak58awxJ5wWsMgFyPohEv8hM+q1AHHV7
l7VcvxeP8ZiWVEbBLhKORrIygBF+sn0OTUDyMRoLagL21ew5V3CQToEMUL/47lBkwK0iyZSRjvPB
4BRQ9BAP18N8cGRExAn1WAikzZSZEGP4npxEsIllwK+/6/9Rbp4fm5aaBg6AUtopW1yOCriJeg00
hWcG0j8QNG+T05FJWj5ZVuryUqghEhYFBd6WCcOwALJUHh1yQCTNB3I/cB4EubUiecultUHKF88X
sIWOD20nQqA8dioaIl4lWmwbbnfFfwrWgzWijkTmGJKSrbK1uYj1bP//e7fOXDsNf5+lVFTf4ylD
G5U35OVkEXIZloUXOjBY40yyrCg55JL9ylyhsFATO/txdDm7Wvs13U+fUwHIe3Nn7jUs7CVQU2G8
h7aADOIDe47U/6ULue8QPQ2ZwhEODcddT8lUH3ZEr0Oeb9/iLF6CBYNd1XUT+fy7FXH6KhnRr7qj
eX73NhLW+z/ZCpdhOGQvC4kAgK785DI382ciPfRnkM9q/UyZBF6mWEuxcHGYQySuurQqJdlXblRL
8ALO8KHaCBT+RPQa/5PnuJ/3nXJuhVZcd8Jb0kxNaeBoB7/O+TSNEmmEsGlHpiKi0SgY/Ni/K0z5
JEDQ9PzvunbtTCDFp8eYB+HXl5Y+ujOw2H2faA3HE45TXCVr+OL+bIBQhN5IkM7tyI771HgPRagV
Eq8L+4v72B2tAVYjOFOHbBMX2dvvkoRV5Rh3mEQVIxBhhbMdzktK4H3JEsvf8oIMcIh4bNwOOvaG
a5AzwNEkmjj/yk23opg3QbcPWdJRZYiGuHPLuGyxFV1ox6V+CwpVFWhJ6hc/H7+nQF+Zf/WVa6bh
cbhgIiGiXVbWCDqAOksW7y/bMtAO/cyrSUYXKxtSzBRCpSLvWXLnQ8/96J8Wyjv+ZR8AoaqwaYgN
fl3dPm14jkNnd8dnfeh7eqq+BrJIRijrk3T06cQJ/cnuF0Ohi63eXa/ajyBZXXZ15l0jF9e1oO2M
Ws5jhsUjVxoXX2aeF2dhb/4rCBfZbGGIWykfH5O4JSjMvnk2S+OEGVrEki2o83WcyDhTRTFsegJb
nLuTIAtp0vw7RZobez5oIgZFHcRNsPerexWz3qeiRmWQY0qopdbt9Ay6neEM0DWvTQaD8XuOodgB
RCr6ayWhBMOcksYXfb/IX/ioirGrtcssJrjvYhuRYbnuLvb05M3KCZeGN3Ro8SLCbUhx78vA0lTt
Po9ZCSy00Y2xkIphSgAA7SR7LY1wygo4/p+nmkHo/g9acr0XRzpfwp/Cjvpn7kDRZrg3MQKVc23u
gidh2jD7UObRUdKt6uGSzNu986ucEfaNNwwHzG33g1iBEB6ytoU/GZjT0sPB5TX0XdcSz3peYEb+
js3cfMBx/4YZZA3ztNDwRqNq3TLzxlu4J4VE04bPQdI8ER9KwOVNV5g7/zN5ofs8AqhLelN+avKb
XXW4hSwuNQ1vnd8REIIzdEbu13FHfe8Jf8QR62HUvDsgp/3pE523d09W1ijmyqj0AAVYFFVv1qpv
qDsduQY3Nux2sGR7lOAloIwifyNf8BbE07Djbtzpvl9pmVX/mFcjj1to++hMLme0j2sPvUM8VW3k
ZuDQi1Wqe53VfO4VNGPelXrP7zjrOdzr38dKEhLpaluTgmpbhJ3WaC00GJhFXq9UXHBEz5JhRUTC
hg09JXfKOrYEyvBGr7rdaq5CQfa7GTzqvOlTOB+KlGBxvhg0qq6YIGILgKOAg8t78Ks1uyBZm3nC
ox7KyFqlAdn7J/z8N+TspqusJuL9H1mAbeoz9RPEX/G3QqJYmzH/B/hvpCb8NDn/74UAIJhUtlTU
IX9XTCDU5o0dJ1MqGwhOgkm0xQwBatnzlPlixpvgOoTG30CvalHGLobPRuQ7+7EURSPkOEYLyL6M
Rp1PW583J2qXT93hziV4q24d8LPGpA/BHEUnRaEUbwEyukcPNrUVzDYskffWXXQGvSn9KAFvEm5D
H4NNX63jN6h+VmxKgqF8LnT/fYHNCHOAdTsKi//eEykrKLEgDFzOQRFaJ2ibQgceOwMQE3BmRHiZ
7d24WZ5ATxOYLjPov2MA86RfMxuLctmmVAcGsGqd9aKqjbY66R5O+QHiEKrxF6YOSqdd6J/YACF/
OuwBUSnnlKSRMW5s/18/V5Gcjder2M9x+tht2kBwqmJnRqT4rdrtptUw6J/8yuMR5sHR6isnZgLX
hTYk0zFNO+At1CDH7UWDK0uFiCs/MMM5t9rN/5Ci3gjAvjqy6+SR9n+LQxTKn1kJkN8Qoqvj1JRG
QUqP+C9ozBK9j9eIqLQsKuiinMOAApYtXkK9r06it3TPG9lH69hlvns7DNxS8KIMSnALhALzrvLy
tz173xby1Z0rN4g/koy+t8VnlDDPycJECDoqu0GuLH1/Y1AmlpGI5vHQ6PXvm4aXqB75VaHdRmNe
DZ0p1VV87jqZ0w/klSG9Sc8Z0ZYNHu0d5wSGq8JuFU4gMlQ/jcGy9Ft5db/7yyK4tYQVhB3rMVIV
gHansN+owpwgTsc6YN0ujKuq7O1H5Urzas1E5qvUQoqMJNuqUxFd1LnF9wajRBwrM/BwtYWhCnFC
4nYC01nDlpvUWQsxbIxFZEfILCKlYOU5zAjduXaVHRnrs0vQnEFI03yaqv2CHUiOwPliVrYxsUeO
jhKpyBIeMTHBx6tgmq/I1aXhfCydusR5RNqcVYL2EQFzmaJFfhWudRYS+ZNNEBRraxGDDcg2O9uY
54r9MS87tyQXb236pXfgIR+E7Yj/EBU1d3LHZoH6hfgoVXF3cLfuwfzm60zj66cAJGV7hPxnpIWp
hnGmRFRCK5P8dSpB/4fMQF/3yqBgN0/oraqNLEhtQlbMJ5wWDI0cqYmS32wnv5DJ8MGzZVXFx6MR
FMw0DFN2Xsfm3TXIRgxZzt502T2ngR/EPEYbuBMSRrDanv1/D/vVLNDtfT864/u5amvVhYToaHmu
yhdjgY5Z+arH3azwnTim1mWyDaZUiRX6/zz/C6XrFcHJ0qotAHaCI7EEzklDL3wiKqtGj0ucjpM1
YQuTsCe/AIWerqqKU7Y5j7RYVLmsw7mnywoR2rHqmcOJm0dVXxG9QOjf2Qknk1c2bj0YY729yil8
ZPbEoqc2q8DgBlhxfDUYxcp0fXk77nw+/VV5VFoU/4TsqsbpCaXNmCeMX0vrl18/VU3fIbuIG7aB
G/n/rZbfBGM1IfGj+S2UmayRe/hWpDioWqBQJQHT2pwHd0ZHExxpAeHLny7/yvYqSx6cAoTRbAmo
LtP1dT9iTSHBRJRrFd9ksNUBLEM6eKsfoQKqG+MWj/3ziJLXfSRQBhCjdPQmPUz6bt3v1oWM1Ugr
vjzYbe+jIarSfOOOyT2MhyXF2rkJ+rZGltqjhpXCwvwUSrTbbTuSKwSuM04SSYoqyWuzT804pbNQ
3bZ6CJrzcg6ryxJ+IbUuLqQ0lTtnUs3g1kGDvfxBXCMHSppX/0YatbNireEN2uNUMOOsSAv6+jXs
SyjttBxbO0ajx6Hi0RkRARY2UYI/Zgf0FfW5PmPygPzxGCmrdRs7/lmj9yFXvPhm8R+4C4qm0oXg
khf7wBrT6fQL0UZ7DyRhSmz9YbDjodNqmQD5HiLtaJUZIYlyD2eTp9Etmal2Xhm7hLKfdiXqQWCz
B6UIYA/sGudvVtz44XEJbAYvVG86Hq0sHhhmV/kayPO6uk29DnJmVCntrcgS2s6/Oh7vcP6PqW2H
HwzWVZjy1S+H+rj9M9Rrs0ZyRQRjsCIuG1kuWSs41CmfbLrkG5diYlK9139k2tYW/pE9nTVb0pEm
bzsaFXZM0MAGsgFQgRCr1maV5wCI8nzISKw+Pf8t/jL+xaWBS3TjiehPpeObUnO7WJ8o+4i9uZMU
oa/IVbq/9PElfsY8RNuFssDr79ikfJ/8YKRTjmyaSvOPmKwPynyweT6Yuj2kt0WyfLTUWKW4+qTh
AjKyRYeE3gsfmo4dXD6/BHQ1Cc5Vgflpu3/KVyDD+Iebc0YQ4uwgV4AslgP/KUZ2Xr5RInEf4kUW
E1EWvpDpC76Yoabhq6f2UoTcss4NIgDw1JGWrTk+meIh8YsGq4BsY7L96aCpPWgMRwiCJv0CCBcP
jwgFQppZGh9Jgdu0Sl5/iGtd4aFSJxNS/fi5sdjbAxODw1eXWFdXu2ZglqtX1SV5gnFL4gGSv7Y4
lG4VSY6dcRbej+3HpkgDQTIlD+79x90y8cL+TBnKKz4zjIMe5izm1ogKo5JkxUlRjI9V1v4SZQ/+
vpUqNetVpnsXz5ni68zwxukCVPgqRb7MkC0JUD0sf2XrQbSFXbkwLMDtIIJA4Dm3pEDS1oigUmCU
plwTKM4epyeVMx9Q3OcX9SXgv34TJQLSK1xLTMPLc8wQu7YwKQdoyd7VsMk4pBcHJXF2Ty/JPi5f
+qwLokC0JpqeD7FD20+hOMLHdI9d5AoDYyMThfzEvH88p6yZyaKAwFOXiuAkdHAywFCj+Rlz4lQT
s6QguI7G7u80fOUJWWKD4Bs5Y4jC15M0PPagJBd2WPA7tZtZQnW04whFADxvJ7w44mIsH57xtqZP
1G6WuGKi92P6CYz+WbP5ENYxzMkrA9fWkEERClg05zZgJuJPZmhCKp6nkgCgMm/TRb0KGSosspvQ
GyRmfGnOlDza+r3aoWbz+sCSCQydQPBdXQPlTLBtHBjeVjv9jLpZbRhGH/SRAW1eLDhp8SxujEbQ
k4nn+Yovw0AbvCI4vqXz/PY3IhWmPy6TWukE31CiqvrPbzLlEc34WhvwAy2yyJYAH1Nze2H0s410
LBDQS2ufAMODMljygTM/UmEbx8IAPPEewJF1O13RxJI0RymAbwr6GEU+Nzlo8YXQ++zTvO1bkpHJ
Ur8aLky7DkBtmsrqy1+qMclmdX4/Z9+iPtJis24SXP9J2b361IJwITM0TVCfa5Eg6jCa6bK78rC8
S8U7M40DgPO/YUqIRv5rbCNtJ7xDS2LprDoWsM6bQy7ZKU9O2JyPiDHvsLjGSK3mg9XlUvfkn7G0
Ywbnkd601OcF/aAoIHdh/hRdSdLI4PKAblbYcWC/AnC0CAsKsYYX0o2wV9+pkuqZtHZaLQdOzMNR
+ciTCysCVV0f8gpEO0jBXcOTa6TFd8AEQt3Vjj9WJTNRwbSQmb4AJYV79ic3EKi4yuyXv2U2XGJk
PtjhdaHUhzmmrbDZOrFoa6yCRrVnGP3M/w5HkpYVN2S9rvkDRv3Nenw1FgXBHVfbRcZcEvtrKq6t
vUuSpSiSzzq7+InzYiIHVq62Hj4Okb3kYRAbTvlYRnhgOnK8KvIurH637WqGgF28rrr7055aI2fL
Qkn1PPgRSe1eQIOXV4J/kme0dSmGNKzT/BufzZyv+/gzOuwkFpw2vRqGTVVUIksr2rRHhzq7JwwS
/HQ2GFxDmNrDf3DXWJZqckCNO1kb5HChTcdzHQCkKUkBsLbNGnUipeGR/8sFXImJLQGdy6cQzMb7
l8Ezxwhxb1nR4l+WkBR7FdWg+FbH3ahdy3DyfUiWqmFF0EWlSJ2EnqbU4YJ8dh9ACj9bjCgL+oGJ
zd31eeJD8+i2GeLD5FFfv6uwHvmGt1VrxXNWIspWweCQuEOFxLDAk5/6TkgAotYYK3CvwKCDRwKA
3DUVtCzucbYqunK4VEui50TFyF0oUrkTndU0TycjuDTMf9//f27fkUSo0HQryjfJ2SGHEjrAe/ph
+IP43ht5mkQ3XYR7bkO934cYerPADmKE65+/Tpx5IYy/qbc0zOUKLqB/3QvmGnFAkJQn2fP863pz
S+mgbttkSBQaI2rrtv/yDlWKuLDmTHAxt3w3HB4b35lMhY7W4U0WusnNC4+RmMT4cHfelvBN5Nxy
WaXX5tldHxYeLAchHEvBYyiYpZ8VoJnItNZ/JFBec9rUGg1xDm64qTT1dMrfpk9qoeQx8JLcFxJt
huQDtegIi0PInWHL/mUikmqjcoOZRiVjvrWYmPXFvrxJlJlW6G3mdJWj+CnlFK+K5nTun0RAqq9I
fjWQoNnzK8JU4OkmvJ6alsqCQJeJpWLXwt5p3cw2WJOnYyeEW+lYp4NpJ15fEGuDf5E8k/7hC4eI
kVZqiVngK8g3oDdF5gfduaYV4m/QhVbdE/3BgUmQpCx5wO0HS4te/IKwp3HsxdyWM33JLhkktJiS
Aqsqvvxrazc7CGFgLCb0PbUESZHq5Okxm9MChfAjewqDgoZbDjQEiPZK5mnJq9hnt3D46T7Pd4rh
O+GYMJpSP1uC/EPsa/3fvzXeGcTQUHGccK8JmbCdt5XV3vfcoHhTrwglPLY2bcKFlHRPIPYWLuEt
uogq7gbg+pKIoedkQLG9Rlznfd9DAzYGaVNbyNsmq0B1FexH/DiTz+Tp57fLy00rxDWlqVSQBN3U
0wyKW4RSk6sSUTEFV76hX7pTwqzPKR9MDgQkJFOGBQygc6seo7JRv0ord9QFsijMaaCFqoX3pYPV
+Fd1WJtmcqYBTBjtYCap0R9YfjiNI6Q39193qe6aCxeLHvSmgKc2UJvmJdI+sOdeDM+MTGCxKdGa
cGCJAf8LUsJ1OFWb7+Bhf6oy/L0gLHgmWyjdpjGngXIISOBytM08NcyMFRaxp45SFZ0PQgRa8sGz
PwpIeE8UDnsR41lUs1m1dZtaaesMGxZ8+O9lCd4Q4TPKKRWRa1DDbQmMQgKMNahuEjMYI/JHeE+P
mXVqr+Q5eWxl3KXe0LR/jptO/mFFPQpEGvxFYp36b3HJ2s0hLZMDEiSCLgoRVqTx5oVq60prLO5k
22+BNJFxWlYCgB8U8SlFPvHsPjejsV6xk0Kgyy+oZXFrqk2sJX/VOP4+kn4bM7Ba9+KdHzbmy6za
c40O3UJReOWxWQNEtlq/1N0obkCxp0tDHWQhweBgfBx/YkVxLfs7BWj63H72OQVyJsHkx+W27qqj
Gbj+tDbaFrVrygnztRouQMxTiMMSXMXLDr7s9vYNu3i3lLzqKBszl19Cz/haFICcmuS1am4hQs0C
/9SMyH+yOPwXFrd0nV6bazEcB0ZNeVnOmHgVMNFQkOvuW5r7Gw45adX7WFS0wF2dA66t8O+ZWpKC
Ii0yOabe9u/JY1H6FEYn5xA0dazguwQwF7o8fzmqjn9x8EkYxSNX/NkDyUxn+TRSNpdDK3P/OnKe
yBWWXEKk3vKUrwfPGhc4EbXytX9wXVjkbzN+cTWJUzLbwaFawV9eeI1Vhggt3F4sRqa8y/MnzJZl
Y457+Npux3nFT86OVWmRK8xWdXB4YaQcgNNFf0yFSLBPwggHsatUEfbXy/1Km8A6M5u/f+FUUKyo
jujURvtlnhjYfxEbn6k8NLHGpooaS/7zhQ08bubQd6wokBx94NwKpRKo3Z2VMWepzJAkiJ4smD4m
56U0arOaBhLnHZ6pWj1F77kelZWfHFvA8vU+Ir8YBE7fv3AvfbDY4GBppB0Ps7J9+d3Nyhh9JQML
/5SNTIHxlN/UeRY30a4sLYt8+cGr5dBCtN6Mv4G9Vuym481Weayvy2IIK1Bali7k94Q0EjYlS04D
15TvkhAnOOpd8XONzLoA6hIwDY6UPkw13iMKd4Xy0w8kR7HRag3rn6TRwa3RiNxm9zbJV5ACu56L
rD/Zq7z7xsssgCsofRt54xJQk8i1HQQCtXvNC8YAoPkbTxbScZHL285jjlCg0KqBGJLf5zqPAIaH
ZohSua7+Ybt3rIJrOhtPktL3TnxL4p3PMtGJPtrkfZTs3b9IwURgtKRYc5qFqdopKT9rP/d9+RaF
kADAcJvKriF7orKfzyMmqcPeEKIaPMR+RkV80AnKPsM6yMv320r8NOwgM6kL3Usv4KX8axDMf8ZK
oMukC4pNq53lwIhhaLawvWlhc1aSUJwXpzlgc04k/gCo21EyV52r3w5aNuQoWhhoLng9NZ6LiKQx
NmilJ3w3eDiQL2ouSPnuz1Tkz+g2pg+vGxU1uvC9Ih4HlvJKZUTF4vlHBKV0dKVWwmDSSuvELg78
UpIbx7GJOTE171bUt06i6omiJwcEzAsyyyrt6V+z4f18Sx6xoZRnTvDBl2GSDZr7HTNb+R5YA87T
5CJ6IUZcf5v/hHhzAYij5Lxo5IDKEGn9gZDTj9VrU1nusdCEzT6dS12bXqKVjN5AK7gl6/KilFLI
JY/ECU6ia3jWilosftlLaBJRYw6Piu/YMJEHwSmSx1chJEDJ5a6hRb5G9emu6Sb/mcHeNg1D4p6E
m+RZqvTbNFRycYTLDeGlK0PPFV+zgFEKl09bADgg0iSidwNVHeUAe+6gyEeWJlCFd0LxUdX7KTrM
nnP1ZXEgCk9t4T7DyrN1Fh3dV7oFEmBG+ZV/2oTwwG/crEZ21vCs+39Wtexd9hZhL3oNG8UlBTgd
HHV2UWjA8+IpNFYD+D8M7CK9+7IvOvhQXtXzo7wSZx7ROhVggd6SiBn1ruMnrMtCUU6CWScm8br4
EjCWFlF8m0jUBbQMuVZ9M9TVUSTnNamaPhjaGAxhyWOA3WQcgTKZK91Lp0ZLFF7FkbvDgRYGd3DS
L2hyWOl0woWUATRhepukyAb4XvZHJ0En2t0Bi/NCpoULwe6ci7WMjoSZtfWUPxaHkzH8S9iribF6
3ItzL4cWqbI9O1H91085yt+ducqyQIg9up/C5H3VPGKUgr/k7vRXy5WRRtQS6VOiYYc1f1tbLQwn
GyucbV8fIwImKk/o+RYT1HrMNZc12arNO8PLD2/NjmGbiflmlwjp1Z0XsHc4T1EM2bfzpxG3mHzp
3q/0uzeR+Cm36/gEuyygVwtutG5x32PgVkLXhYMIjTs6KcBmkdCzJJUcRIOCGsdCQ8R7332Uz189
MkHPQ/ii+RatS6hT3H9wRZStABetFa+eo1UwwzD0pMoN6fwkpiuOF9cSnaOxK7Bq0rS4fUstDPlQ
wC0J89h30EGa7NNIJ4HlItSRRyH99To++M1KgUBGu9Vm4h0Qibrho+BISgU62GdXhm2otZ+29ps2
F9CBH42B9jSaWxWgkecB+xLZY31mec78FNubTcE091jwwOue+u6mOu4dYFV2MhhcfDp9eH6VLXAX
/065JCGb5z8vytKLqMZXvl+AzcPxFAJZaDHVbb4K2PSIdTlj8qpP/96OTh+kRqNaAy0g7egmd3A8
8LeHx6Q9xy9AwK6BLuVAzKL/7Vz3J07dsFZftHo3/zwDyatb2YHGLJMtkj9UYrTV3zy0MXKFOxJz
Lh99+9/rJiZuHM+PMR3k8kbnXwuwChn+PGL9En5BjGvrtJL5jb9jRfhUPhp3fujAI/pJG3WC0mLA
uvtPeIdXRfa+hea988tllp3uVKhrMlWGVETQ69qHEtU088+Kb0lNWjpjF5pJ5IG37AaKeoTWQLqT
CL/ev+DW0uBc+Xr5b3/AxSsiw8WrdGDmxwrtSFb8b8fgyh7I6PrP6kGT0bU4q3uNTC6dOYTncRVw
TxXatxPQSRzd/NwzSaREhmICw6kjHegKu7R2UvN5S5VKKBCCz9PJOt4hzWGyXgHPBkTOJyHPz4Am
5U3WtYK+nfAEChedaQ5OtO4FUNEQgUmg12C8ILzH4yposG+rdDW/QTNVyID1rkWO685k3T+nkpul
J0vpdMYMGRVsCbc78+ubR+mP5tBdv57flu3HVUi+on1JxGO5YdFaG7j+iYtbNUgPV8BrpWHK/9a1
4iRpZVE2v9JI5Lf95tXZqMWnjaTLBfEovNfxgBP4CoZjQIaf6n8nhzU03WfbTcBf+oBZ3ScxW9Zs
3OOzyyzE6JnmadwE0OR+TORqQhBemsMDq2yX9TL/zDf4pUqe0g72de/T4fvdNgXchcjNETsCNVI4
5V03wlMMaG0F097b6k5k2dAvET+YWxOoVUb7QByPGmXfV36WWe9ZAUd5qPw3SyM/WWUUwboLFl8b
1aBp3KROXvEQb8VHT/Lz3hwYC3rRkLzQIc+GPPK8e9BAFSV7IctK56qHHTqrfU1M5Q3//CbhKaAL
VlrmAuLX0/b8g1BwSCj+M9v5vPmEpu+i+JJKOnhCRsfSp4Un3sGfRLH1laIh6bQ+LQBlrjQPjx8h
DKLBEGjo2Sj+Spwh8bUl1sCroDKz1ESN7yxY6oUK7oZ+jtB2rCsP4251buJIrZkru3/+ukT89siP
Ux7YUtZp8jibiZ68zr4Mn/k/pXfZa69Wh3JZCbAnaQEiu8jOBWnshsXlyXmDFpriKvVcFQi3KStS
mdfxw+o8rU1aP2qefMLRHHMLzwLtMk4q42nn5Pa3BDW6FtMNyXVzll+ad+7wRIOrq0jcAUgYCV7g
1B77djFXhJpb3PySA/sFD5OSJ9qeKA6ieb2Q2JOzMa01+6oEF0Z1nV4JzrVukq+bxYRV4e7f4J9Z
3m1w/jRjR8kV9GamPu8sXwuS25i3sZYiZ530RvKcUdEdY+LJxXBpbPHoEdbVAIxCADQtI357UINV
AqyAMqR/mZd4N0PCxRL1he0FMJgT+wOUqLuiCG5nP4/FpCkKyHR79Bl8TK8Fm1ffBQ9/im6jXoQD
YfPexBE+14dE3Z2QhhQBbxAkrOYEE+lzLY65DxSvRx62yvFwIVc8MIPbyco+z/0TEVtxqtvGieZz
XIWzXCfZCRBGnFfFaZSr1R0PrcZH9m+6Suv6HvM6DaU8Wyc15BB1V2Tozn8BlPnSuyiK4qk7uTmq
hUEoq+9UdwvwmdiVpNLjCJEJbpTUU51BD3GqYSZAhe4dnbb0zt7t4E8AwvHU1EtRqp3BYPjXvluN
FVqMwfksNdFhA+kJ5UHXUkCWKfovbdtCskfr/ocsD2WLl53WDkuuLWpI01ovMbt0Rm0AE1R1NSpI
1D9bLnWcC7KXjWSxDbHYATyaeI+zPJd3628TKxj8M4N10o1Q9YNvY632w/x26bj6sRjNw9h8vqym
/K+meAagsxPPMoHl3UY830r9bCayor4JRZzvyMnvQ+D4aBzwPi7u3ejbbERNlcroLYV5oHBb0Hee
+C/Z2JBWxpbVsZLkVk1xnQr/yoBuDIRveu7Tx28WZ/hpnpUwD8k2VVJMdv7PkuUtlBkpxSGO/G7u
vcBoDxtbDstVyLViXR9UFRJH/mQewYbKtHrF+3ozjqiEIqOU4PQqbQIpZU+exqSPWVrFMulrVaEF
DcXyzbWapKWZ84IJYve1/5PXUG6CtZgys401ELPRbVPm30x7ePKmJ5BiyEFPQhuQn8NiDRZI1nmQ
iAuDp3avNoJ/NLkUqnOdYQZHAQErP8S/GAICa4H1jVHJRvn6YPK49xz+lzj9nTKOgEABJSnb/tp3
VkyQErsDIkxX10tcH9pE1eT28YKAAWj5srAjtM+MDL3AOQ1bqt/4DmVV5P2M1omLfcyp6C5zTBAO
UWFN+JhI2ae3Z4UzQv4+mzdSBes1tYVDCVlSrZdmqW4Sgw9/U/nUbU07RaIemfRSRvF2MgUIeuL1
mXVu3RohT/P0FxJPiAteuFDVL6I6tg/oMEuKm/k15TPBt/+c4AjSJy5GUiZKkz80ZjOeXg9zAvUu
+hIvdiLfAgWpFRBqodvjaiyLVVbeaj3a6o2bTUiblaj65Dd42fU7JU9pFbsgVzO8gMECe6M/FmfU
aPeif3FDkKmbm+zN8O6raWl11Hi/DUoXJuMl/y17TAIruaTwZ6k2P2/GzKS+IRygcfeFCdc4JHge
uTJLfeOpFPPucyLUoJntlvl263bBfwVd539U7gIjIWFOCg4W49hEgfam5nqRDZuSUii3iQVzkS12
imCv7CAO0gEmXUyYGelLBS1ItWTTKTMMTBsGMB+h1qP/cTG8gLTbqBY4QFv90d6by7Q0s4ppK98p
sCmUl3Brq8A7idy8PUWycqC8xrmhXEDrFEThyA3dOZ7FlgbA3KYcktxhLf36/hK+v7d486hsx0Iv
Wuca5zjRPrULMTCPn3Ri6u7HHndIrX5lE3pMfoIYwAeZrlIiJ9a4LCPWluGban8sXBXpKtCZtKTc
xKeOf5XYprw+44iEuxClVTXoXCl5TeW0S4Y43i6L2klet/HkrlAsq6EVZmPHL2UbhCpE8ZN6AbY+
ZUpRb5v630K+m9RGuAog0foyZzb13+9TWkCa6vLGksbGlvy34otdrzxxHWm0ceemaqyyvTDm6tD+
x1+4ewGCDfDtI2cqaGKXThDj7R4Orhz8aQz6Vewzp5fkYsIczrfC/q0ACFmRtH543gNLJC9w9AYN
Re1YUIJ9LYzYSCCinyjfQmT6FinAhHo1rOFvwBmeSTrHPqK6HrYMiegaEPu024sbhYIHl7O7CsiG
PpMSNd7cqi/+RSaIS3+6e49NMnWdfRH9X4zpE6kyhLQ4TDk50wOhrWYsV5IQua+vYVQ0h98qYM9h
oiCPJ57bgLpDQHWHdckraPMmmsA4FOEYfod0IZTOu6VpIr2LGerbDBuBJZmxdGx32CF1xKjkkBEd
zDc+tfDf2ttXJpkATKDdrQo5ya0bzf3A06MiuXkSQjOjjxybdKZXawmkMH530t6CYoo7tIn6dWfu
wMt/TBUFbgZ9Ry6BXMLN1Oino8CfMcoMcUcvOnWYuxaJtGN1dGWUcirGXYeFQuFSpmcAr9ENmZ3+
0ak3Pp37Khq6B34fVDA+aHnBtoIUgBe1D97k/op+cuOVB8kOm/1BKKJYiDVREbWO/lmaBvma60tV
vDcTltzhQjQ0v+mbQofjOzXYHCtGtVhTnkQ05ZZMf92iVbQbMiTslzfR+6YLWGPn7uEBxQi3l9ID
bTy6cwUWWxXu0+AYqt+qC1W8TnLBgKHSNIjxmv5fxmlhbnC2lvrQpsEPLxIulkVg5HK9lqK8BJT4
uD2iAEEMe54THO+J/e5CVzDuIF2ZwpU3YHt6E+2Uus+eb0f5x+TItjWj7OnJgkC1RPKECr20tQaa
86HrViB2SGPhLlAGkXFwxSakhF4IzXSl+5ECgezLfjBpN8ZPIz4OGyVPReTdZOuzHkudswaznyoV
R/Ykl24qY3qkOm/t/WH15O37US7i9ogxNC5NRGRAy2+c/NNxRCOyFfuKuI8zSYnmRVi/bm2SzLQo
7Vf0PsTDggnYT6lY17zTD4+WBV3EjVUYwDbbfPIAtDxLLYhEzfZOnBQTExQcMRZryieIrgXIjPay
XXhZKFQrNoMfeUcQyzlsvzxtbv45KJHWcZNQQkJCukyOmVBRrGO+/aXROd6coP3BmS9PMoHjSMI4
LLGrMW0YJclWXJDYXldLtXlbIcSzMuFxsmoC72GTa2MSDNaxg6KQX5p3qSSkJnI8Bl7yHO6kJac1
4ReomgmZRLea2EpPHMvUNnksqsrYYk7nwZXxZnzs5sPGnd2Sb7emds4w2PkQmXgtZ1dl1Yux82zB
TJk5DVgBMz+cBHo2Ry0hUv+GYzMl3oHGeUx+yphTLvzScz3tsUIiIwHl29+JA1fAbWVc0nRLz9CL
c4XXlrgTWKSfNpK3JGJS1GOCd1Q31f+Vme9WJoUbxfPv1+eE7FxwBRqJIicY4ThI8MU1MLHHkV66
ZrH1BgDZOy30cLIugYcbjScCRAM0RMa9OxFuq1fx2U40pyXA5EiQ/YY/UJHBk/dQWrzrPvTDDMm5
/+Y+V9auLnoeuyg3UN/r286emfHVOSJoMobu+Cvo59lCAJC2Tf6gMFBItaSYJHCgM588ZA2Job5q
s2DiI7XOeWVnRHpWloRx9kgcoRiMAdhDD34EugHkxXKIShfTW4dwpBWCQZ48eb6wrkRBOoLlKYr4
9DoFBG93v7IalENo8GDkhrTBr5kfdv8vTjW7w/5aTopaT/C2BW0TmivlSCPduP1Zf0dldiPnk5vM
n8wLx1QcIIOGPJwt3WZKkuSrOpR0j4tdk7b+Ai+FgV5CnOAl0+QVTUUkoTH/EUVHB78uU9HQ3t2+
Fn0WbXKfQJCkLMXLolXlAFZJrWWh7E5kpBGMLFikqTd5WkoK/7bAt4lDGnPXKF+7jELaRNtBKTFy
b8387aHU04dHy6OStJz3clwQ9utzmZd8gGgtYvI+7piM23NYIZPStLXVSpVVKF/+nTWmknm77G/6
yx6hC6nqkSG4TO+a1H3vlRZF8sv0hl27IcZORzC5EeuMAaLSdLNhIN5MxxxXGeYHQgk72UZq6sQF
GDsHtnB73fLjhe7AFyhrBWFdHXsnQFBD0eAXxYIAbB6cbA5IAG2n4IUiaUh41A1k0UvEFZ/3F9Pk
CBJF72z64BS4yzCEAhRUa8mSA77ysiLXETWd0A9i6xUTGbuxqSmwfTmy9gbBays4QzEvshTvqISc
UlgFEKHxcm/evMOkn2VFhasSXhS31zDvuPbADw8Pu/YZOBG5LZ4fpwx4n3HIagl9GLADTebpzXPF
d5iO7UCkmX/xCgUG//o4TFygu+QSBo52iDl7c9uMDg8ciyjmuBCAvQoAB0XatPLqAsUj5G6wWu7U
31qT8PuwR1sEUuuJ8ZxemeIEwMKOAGx1Zq63sGfxk+jwjar4zTW1FUtytPHsOzJlTgYXehx49CGa
ULQ+SPJ7AGh6dF8BDrz6FUK9TKecY0m8vTHYUhxwHrbQy5mHlG8PfcX/FINVjj0tXE9o8jtylviq
dozHwaulzMLC5Hd8TJHqVFmpT0dhRx3gPKL0hAvTkg00tCxPbSZzjh25kmmT+dn2N4lgUxL8Reqq
BrOTvF/3ilKHnngYaWldJv460RkpI7/ekl/SDIdWRRIUeh0WFshViZ2YO4/e0UUX/BHVqHKsLPin
Gkki4XaACnjUFmQq5cS+wp7nU8Z1JXuHCZl+OAnBkGzgICc6fenAiHj8/3SIfq72Vgg2vzWjrKjN
+lu4/axk3jIpVG/0SD7vnDqZ0T3laUX3bPskDU4UgZqsFN5kXf5g7pAJk5CV5MfDg0sNHw/qLkG1
ayyeHNQLLa4OwIHq296Spimree+LyBmdUJ/V0AiBVj90KoLYNmP9Mfj1lIZQBVk/xWTPT+1uBZDI
dCU+bmT29LZkwFYgiu8skVkbTHuC6nuVmY5/jHe1LdU9t9ayT+pWVd0dsUd3+Ao0Tlh+n44MHFxh
KRJVTyaPn1ld55C4RVsBT4oz5zMudssruzTaQCeIjDd8zFbqT4OWcA6o+EeQ9ftYPylNQZ5e7L+e
3es7gkbNvH8/z1sfnZ5G6avZVkjaKPox1EvP2b1m+VdTSYZins/zxKGNOENQ8NH3CjM4Fzc9UwYf
22ehNTO2GzNkmzxM6kGjRs9Xiv6oNR5Z1ZdknnUz88oyOZqKh1uyqEkp1Yp672LtJMlSYvziohol
cGdsr9z1qDnlrTSoiCFMIkwQZcs7StiZlFp8dOG1oAOG0jJmB8ryL7dlUNdfhNFzVXFt7Z7kLKOO
Q+QoaIde849qt+NtoddMKqO4QT1Cwnjl3NjlHhDUoSS11jMimfBdy5OErZpVXYM/IRn3blk4329J
GXuWgJNZumL6edNN1zfB1bi9YgSh2Z2HpDMzwxwteN8eH8WCGmpqwRG87UkZXOuy2o+n81avWbuz
Jp8PABZZcwfkqjVxXFspRW4BDAuZswEx184VI2vjXbV9XJaRGirY9JNoV15/xXDGNDWhqGvXU7Iv
Ga+C7b7zeyW3L6+z4YK1nJ3ZBndg5o8dRjk2MwRuYZpPzXsw/XcAxKeKI7JPJwQbIvqpbgfCNonR
TdUGumzD3DoM/d6S1kKjzqqjZNdBO/iz+wFUEkNa4a/EnI/5ImKgJMtsLP/0NpkYj/nsP0NNdGwi
SKpy2pJSEry88eqvd/m4S1vTRtaKDsYj6WtSUVzqK+eeK1dF3LPcbNlNJYe8gE4jRNE22nbdTTsR
7/wsTNMBE9elRK7RbrV4xzWiTffRMbEmo9y5WzpYX/jvXwNUhp9ZkrDsskt0bqeXnS8C+ZfC7grC
8TJJJ+XZ8gViPEbqwRmdWRReGHUuyfyN7jsQ+fIJo5LbjjjyyLJfyNyJ1gQsi5cFbr++Epdr3wAD
ycqcvlxiR3mukfNFQb2TRG5OWBjQmOTcmAAQAQhufS6ci1aL+b6HXFjQ4jv5lVU3jHhIs2AttLPi
b5g/bvSJuDCBZeGxSg4oZ0ObeUlIzPrGKtdrmn4GSaPMFUl5XHKjurfryS1q0hGCa1I3nBsksgMV
rBTdsTcIwf5ZvmfoHvcAiuVetomeHE0CoR0CVIu5upoM50B3GHoIrxE1t/64M8LbJPwpAtNwMzS/
W1QhisklHif6t2x/dLL/6DWGlyLuB5Iofq15SDlFEhLWUqg1wdEiLkywy7L2mKfo7SkbdpVOe8CN
6kYgmh7rqPtLuvaJ4nygZbmIGlvWujmZxvH0UYazqdW0jOvTR/MQMiIyzqBCHH3tyuRPYM/TNGML
X8NFeasvnZANV6UEnpNBUJgkPsO6DSA3xyQ6wjAxp+vsOqTQnWxZArlciNk4B518Avh8le+60SKh
QObHGtw+HKNJnv7A0Wt0NBg+wzSaNzqDpijP3XergzJUiG43QAxjfcFqr+wjpm126R6ksTG4U/Ke
wdgOe40lSSsm5s1MwdFxTTDgcOW3LSngW1WO1xDyQ6RH2OuiWyLKVRmaH+DN1dDOwFVeHfP5Qa6/
o48ziDZu1dO+QztUbRGwW68uJIOoklacQhMtenOr+PUoSVgS9lIPOQtY9qj1zeDDblFOKY8kjyV6
aURWByd/Ddll+QOqnwcbg51JwLfacZq2JWHpT3Vgmwtmik30i2iiSmaPJnoExeFAx08t4ifjS4CL
5WQUhV7dCS9nTFI8rBOfry6dkqbycOrYqKYo6+EB87c25Y53ffM62Nv6t9ZJy77E4uMyxPASx529
xgx6VPpygQSep5sDrU+IZOkHPNrSoHbraz9yHfDKhM4L0wGasU1UAZSGn+o7iIhLqkApgw/qVqmL
1eCACzjEt7c7CKZgZN8NnlduxJkUhpQIVzDa0tOlZpqBAvbweuKITY/m0PBBHd9kWw/JRHXMEr2a
+LFGZgkVfpdkhlC88SinxKPMMF+Wr7EDL2o2IlRCcbJwR7ZKkPcMFejOLlFT1dan8NMyH8NnoXPO
Pqqg9l2xl/r4PFI0QzQCnXLWhKU1pa+2ZM5Z5vkT/EkYCO1GOrDhClqNJWpcWLf/HBy3GM3T7zKk
qoImHXp0or3v7zjepu3zWehf9dF8CgHPwyQ2dUU9OXKLmdKQh7vNVJ+m6a/SrnRJV3oCVviqabRv
Y+7L05dGBiCbvynnQIqrDnFAT6UNDm32G50TETZDXOJFRHO1lwcSla+hGGWfgn7j/fw6JmjAaeJ1
d8l4z20m9GiPr3UFvmkxtGSFTtHbXLvtQdd7wqKi1mD40iYi51A0hcsqal2h5jbsFbE80dtg17lI
hjw/FvT8+klcFb09PiKo3T/g/RETCjG1/U0DF4AhIglVfZ43fKiBGz6odP/JyJJ3o5+z0H1oUA08
44pm/2oxP62hGIo/TmKVftkj9vCzCuo4I5mTF88CyyGDF6pbvRZkypCGyYFN+VPwKalVhYkqfHaB
70Jtiazk6JlLu4h1vF9bk3R3tp2pRqdhRga2tcQBZKHsEvkGg3rcFKHCUEC/cTlAKZAgYyKAMGhm
3QYUiMWy+7V+UI3RfkSfxnsPHcck19gm2WmhtbBKPWJ1uqGmkU7U5dnDzMxbbvfdSl3WjX71JsAp
r3L8eu9wXEKTl8T7OP/luGgGbP4exhSFr6a3yV9kMDnQ7Hl8+eKrjpueiijcrIzXnMlBQU1DaK6A
TlWtMpbciVOATxYz5TS4ig5n9vm1dr07rw36ZGoD5fTMyYV16d1Kia51dwUpRaXhKcROm2q5qDS1
ITnwWvbPKAkFHePLv/ZmaogMHynD2xGWH+mmDsAwux0gXfm6OnR/KK2n0dvgJHyP6A0pKnPyi5oX
9cmf+ChBlaX17NJlH/c+aYo/bo3BO82Ip0jUGzFzZn0/vcONdZL6mDiqxqga6GROu9pxa4m/7+RA
SjV+zPdr0qfmKDDZRVrDHAHe2OY+NJFTCKZPVgS16CkpOBYdbWsP6SjOBXrIV/iMovHnC2B38kwi
+RgWuXMm/7uavVC9Xxsq/eGjRKuQ/AKMSJzzkR3rW2Npkxh/xJSDG1ceCjNdoG7tHg7HOEzpIJtz
2w7lsHZU+I79o2EEHmDM6DLNBjygdgtx8w5Z93bDfL90G1LZX5cy/Cv50khHTGu+GfG83CaptrE1
gfGV5U2OjD09c0SHKRQ4tjGVXhDF3RFN5uCvEdBGl8fyoCWXIxFEEhFRiYcECPjEesO9qRRFVGb1
GIbYzn1SpMPxtLaSopMfvGCjzYiRbRo+Nq9Ailo/yqrVsDDpviBAinuUVVrf5v6tZmqYdUmmnS9r
WK779nL50bj/Q69/cRiQ8/trMsjM36apSvE+zZgDPBatGbyZuzXlex0Gj2Zgh4JIjZLP+ByBANye
kv4CTf+m76nJlNW4X99mPiLI8+xapVtX9otvRKNBj7gNaoN1RXTFAY+8Dp9hcyXdwoRDpDHQgdEo
LZDbFTrLCUq73S/I6PjydY4kSi1Dw+7F75NwjA2JQXhjZI4lQLIKyUIx/krpkC+egzB6OKUzJ8h6
mnNL+oGsnoJugQ0jYbFtgsG6a+016iVfGX1ULJRH+rvE+FlKtTNVWXsJ0sV4Frh+zhkbwc/Cf/5T
1xxMKNZkrE9WcHX1SEQKgeDo34xLvOGg29gS8wOu7M3CSYlCvimrhUF9Fest41MuYTFhYvj4om1d
jo/n3bh859IhtXDDd9W4onk18PuXChBvrY7KreLxl8N0c7iMR1pESu36xgYpZCTARlTawqMbNodr
Bc2YJSfKYierUp2Et0OmISwAUyAQQShaYRPTWtAzGH80rgzQAnDrRiOMIsX+tjHQ2NbgwZdQknNN
dccsUpQ0b9MwILqnITq7d03wTXdglKw39bfziK1DNSPkJCQDzXJUJ0ooKkjV6coYpj19OZJX1hVT
r1UrMJ1Zl4P7eu99XADNN9cBzGpE2egXGn79cmsPjL6XItdqBQXIDY69kpyuPOEEydb93YVOJc6D
P75CvVyQPePpPnmEcronr75OBqMcKSmbpfCPPRm13Gy3ytZ06YwADnmHZiysT80AXfzA2J/58oun
c9p0JIfYyt5xKnk7uyRDlq3tHY05pu6b76lN+0MdX1yE3IVHmp752AoLN2loFvJpuhTYFCsT4ZS9
LGproX5zuBeFJKD+rlzBH/DCTHB3tMDUO5acZTXEn9x2S68wQctENPmg8YtOKflMhesF1PjBNwLo
7smg6acLT7oxsnQfW3p6xRSADuSe5p0uLKOz2u3rW4X34/Vx0tN3cl4rk1ILms+uju0IDD1Mn3cw
zIXsTQUSMyd4relonXxXsaYo25btXCg+uwHfa2wgOuywTWpQ/oJVDQax/QVrrgs1WOyHjq3LcC+8
4GcpmMmuNgtsma4xJHfs03+FUlTP5tt9MxNHdNBykAKBUGdCOWECPOn7BSx7/wjj/fPk1uj/LdrV
0WjqtfFdnCPIOD+leX5x6W5bZ/Kzxcn7vjJM017gVVuGaY+y0riZJvsuxt1ikgXnDb6PLiPBqjnD
RUo7H6opmOV7FG74zRgUMYHqTrwEC9i2KhD4p8FSuHoGmfJRxV/hVFG+B3RPyQE8vLUOnVJ4ns/h
za9H9g3z62BUNjTmNnn14ZmgTuDmkDGNt7BzOkgPVV2XU7mXX7Pra8hU7tiH5ACobXP01pv8pjb/
XTX/gw/di0N+KI54BVvHK7liTO0ZnO+mEUEIolfy1b0fVZPi6oH8j/x5Vgze0DdYBsLj39dWQOGR
G0CP43WhI5xIhOX6soNSjIM+pP4x0nF9VZWcw+RbnXR9PZXsMWgF9v1N/cEevBF7MAtlT+2JvMRb
U9aGeqw+VUiVE20sKM3eoohlQGJ0Qb05Ocg8S5WSubW3XIOkRjozixTXPwF+UJ3vGNPJEJJ5+/HB
Cvh9AVNoTfppbWZRYaGgXBn5LGw08bmnoofkcXZqc7QuCF3gakL/PAcqaxjN7YpIjO6FM4Uwz7eA
XKa1DQn620QDw0r0w6ozGcSEjJskqQAN3G92T4J4TH7sIfAFJL2Io9xG2wsuWDpXIaYvSOQNWV2h
SRdoD8PMMsiiMlXdGBP33022aVqzaEQeZB7dHqAw2Kfi2EXpwcQesja+HVPbWaxXD3PxKjc6xry0
iJYM6awfMbhaOkyr01/XJMuILqRx3kANQbxhIckg7w82h8OCaPrv6lZ0ITY86gFEnubYvuGABbXp
zegl/vw5H+n/CHfjP5eP+cZvkRaL+9pwZgcdE4MSdNp7yWvpc04zK+v3N8m7gsSjjOZrSAxY761O
lQmE2i6E0fIESjcjq1jC1CdXZZ4jf0Id1jK02I562BG7WS+Yk2y4SP/DIe9Xm2Ba5sSNTaMGDkZy
6QXHBJPruYJX7oUr+mI8eooU/rfeXuT+jIifo9tCxYk0GUaHLwbVsBezHD1Lzg+JH69Twp1mhRxi
nNonDe62yw4lMTz5YhX5cWuW/SU2XwY1CSJmTCDeX0tP0pLRDncae3IlAU8GvcH8K3kkEHukCn54
JeZ5GbCHn4A7zc1CvtL7VpglgvwQJ6ROriOl/TCmWbiTWtkLsOz5t3Ies8bNMswiC5vuiMl9qfV2
UswX0A8HviqhYWBGA0juVLysC4735uTaIL2NdVlKQpMNeQ9rJ1IoU4gT47O58GtoZR27WlCX+NqF
wkGkr60RNqNoGMPChRF1XWla74oYQ+uYN82/ttUDe2tFoWUawTSlBaCfHq4FVw9upIajKCTbdBod
DUOlde6wPQy8SQiHXqBd8d08DbNCKbaayo2RErv8XEc+aF8l3ktQpPrqzZVOaijmStSmfD72k41C
dvroybtuA1iFnoleAhxG4Oigja1F2vjIeJ1vqCnQo+ht5wCl8AWxQ0zTZMcPoUTpElEUU7TyNOUl
0YK64oAro7S6vM6RdXWFP7FFCGIU7pVjNoUlwdhP8Fwt/SHMBg6I7L5Mko+HGfBXg+moQJswYMCK
n15snMX+GStGMPJfn1ld581NNFwcTSYfWF4tGYmdGjxy4tNjr0mTDQDyA8IPgzi9dhZHt8CmEvj5
39iJ81kd1oyhvoDr+UPQk7vVF00fj77X9tfFMkvs8lr92GQzxRDrcJeD4dyjgBANUU6r28l8TfmX
MJ05OtxCslzbP7e1jUXrLdynkCZt/jn1NlxVdnN1NdT3Yorz6I87TmMjFEjRFqU18oms+Yg3SAGV
VxuNuiogFsHPZLLuXcgXtbiYG0GTdk7L0gvdWYj3SK8NJvOzmHBWJ7OZVGqKWu9y7iBe0Cq9MKds
AI6S0hQpl4MkPo6mGy+If/nPIGzKMZ9eRLO1XtTs949Sz8JSBNH2DAcU+VLE/rsPl0R5PLfMDHeO
UUtgI+fz6cN45QSIwy0ZcB+AyNOQ7XdXy6G9wB9G9hCuxdZr6KV/FqtCLIS+mCbIyTfjOOEk62WU
eHgQ7VHvAleIBnxlPD7keiHKtmZj0PbxW2Dgnu+yU3SMeGEDK3TB1OTid/y2Gx5LZmSDNze9Y1Va
htnqoistXJ61E+nkDm4yKcaH/NGkSU5mTWuyxgI0rxbc5mpelTOF4cy3R53Iy0z+gDtsFf6LsuOw
mKxKD7HR76v1LBNKE+9ccOd4ysdXOkukvpZCBeaXOCuR243xoNC/mOc+hnpCUa+Xq8LuCJPu1gOC
mXEX1aiRRnBn2AgNFfTaSr9fcOO0wrWfqUvEn6l1fnCi/gJj1anSSIjAl9koHvC8rABTLkiD+2CJ
C24Cs2TTbLiM0z7oj57lkSGyO9PtMPcz8ziPYRz7sJ7rLmwmzBOEAHG98qyzKd5oTnujHB4liVU0
Njq9SDxQJDxTMd/ju+t2CnPTBK73v0kn3L0jcM5RktjKGUDM6dUFYA4r5pAfrlWNcNOLwcrUycIR
pNY7rWyqOak3RpZk6KbeK39B8iFKSJpo35ropr4CrRsxl+1Lk0nhU42t+JvCuLeqDzy4lTimrVwW
DOehqwqlr6QcrF8hjEVxiI2Fa8rOkwobfYYwiGXNVgXQX2oqfmmRcx5BIVdtAGrvrdO2lD90wlz2
vYN9ruXrj96XIv0JaQHCA2NU0Tc1eMAPK/4O33hX3r66U6J3MtGEBGGvTas9zfY4xygyJLpm9LD8
u3nouidTGxsVjvzmNeWWGwjWxEXnxFJt0dpqR+yR3rE0mrvRk6yRDSb3Vjrfrio16QHgXtx6Dfs1
mRj0XG6L9RTBFphsliy1GPvXoNEEDAF95eXj1DLMweO5REq8J7nfOzNVVkMlzQkM2zvCu68CQRvA
uUI2cVQdWsiBG4s5G5eEgzvJX1Vc+6w1YF6qPzbikDyDZbEtSphoXbUJdD8GBx3ACb4GYpeFUyVa
imPg58kmLCXAIFcIZiGms9BpSSnTVhGzWpQcKX425L14xfns+6/V8t0/a5EyxgQtc0VKL7SnMo7O
mmv1dY7MAlmV1qsnDYb2W7WfzPldL5ycgmGt01fKSyX1mSLSTEFE/nX5AmTy8dCbFcY8f58ehloF
KHNaL+734vkN0RD7Y+n78OBWRYYTQsJmdwxezofx6HMOpSkSV40KEnbAwBCjCMGFnwm/aSaNrr+D
kvglUZpOp6LXc7hOazCsTr+/BtxgfkUi/k0bWPQBlfVuzJzcEoficISZ0LhA6NaaOV6sNFuU4Y9y
2/j3HQj/dB1aAulGkG8lK9slGzCQ6TU49uDLJ+yb819ahUW/CrJf9qagM4Jk/+mU1FD20+qbDj0L
mLhmIyZF70rbYoF/GzZHni1gwMXkcWOWvxr4uTmq0QUAFKkImxTDNNDXrUlSrFQ3F6qzsW/TbIry
FTpkORJwwpl8xJIJEtHu4rwnombETaV1s5KFcpz/H4gRQwk7LsimiMQz0pkLQfxbO7mO0n+Cnqzx
9zbpRSXvPtq18X+tmPzrJPBQZCxc3qir4Hym+r25vk6sMMro69oZpQxTxRIBHOoCJv6X12IYxtDH
yfCOIiKtBb8EfSFhyQv3Nh8QlEv8PDmtO8tHFoqDQEExQIUuVshTIBljxM+d4SR7XUmUtW4EjHws
fv1wdtEoJViCpJaodfg9KM2wisfG7xbQGTy2ulMRx2wogA1dHHRB8jOluiijNYVs0AtN/PxNbmps
saFlladMiQX3L5HY/yByp6xY8tKPFErr/hPGfUS0e+U6EEmreWoJcBNGu5PbphAxpNazG7h8n74b
iABnMuIHkCyYcOqtGlDSvcJvckVAMI0SG7MsvFJRRaMYBEyh9eAuPUFbmF6PgtxgwIB83H85XEbo
JIIRs43R3yKyhBbRzVOL4jyruysdcMJAPXbLHNudk/x72+HmlzYaGinl3Llf7k5HzqqoxjeCntZA
xCMRMEmPIZN7z+W59AvnY6seAaIxw7pInxzqEGG2YXWhtDnCw7ZkpPR9a/Ad2dzQ9GzaJbe8C43Q
m+V2CFM49FG/vhJZHW6m4ObDzNoguPA3Rraoq8eR32+fIW92S2UgORM6SPWZ1pbjBCwrQ0Qkw+2N
qq8r8wsE+KTTbZVlbvvLyRXkmD0F+lIiUUIwF+/PDCMNcOJiAo1Ot5uVu0fyZIvPz4lmxAZ0XgY9
LCbG7ZO9KpFOUV4RP0fy3feF/0qPzF+NG9n0zLX3T6RuEZsCaF1vXweye0oIvbYvzf/w3bZ5xlP8
JvUg2f1f8FKuYbauxo9kKQ8ftpsQJRA9ze4A7nK4lRnf88QAPLt0RxrVbPkLSh/b7TXhf6HB8+bD
CLsKEW9uL45ZSl7U7fEUl6cYDNZI2WSru5AiTlVsvquBmbo8mlrNBMfhJMfLCUaS4sbhYTtGvdli
fp03oXdmIJU8fwIZr4v8o1lWyxzKPrXK7DdBGsadyu9Xo2SQGJ8/dy5WZgP6UBUoUNJwFwYgEXTa
vEpykoDDUgQtp7wjlus6x7Pe/ZBEPBlejS0COIWSn25LRG/H125B5ZL0fWJeKhaNRWkELkh4mXBM
LjoURgAulOkmrbwG/doNVdQAlnkFfjvt1tz7pGH3dfJjh5gat6FtMFoIVVuhQwt6yB24/tj3kK8f
ehdUULLGT4TRTxZa+TxaAgMXeio7Izr4rRsWE0BzmLqDBBN7ZwOjRg//rUae47znVm06mskaNliY
X/Xj15AxUKC+vBiTWVEysy0JrsWSDaWbMMACgRbraGUJmriz4CZ5lnbIr0zC3x6SRgLofz1BniBU
Dv5z9NZaaBEiY2nbJUjEOFxTTxWtXaHlCWl3aT98AOghldCFhT6RBLt2Q9TLliDKWoJMAafeEr7A
oTQD6MzyTuclxBJ5b/2jySbKrDhRPyKIJtNpt7dhLRkEXw9WWz1kYWgwUz2rI1tZuIHvApSNSF02
bOp3xgugkAr9hYOCLxx/PL5We0aCCVBQ15/aHxSK2hZYA/uh35YRKbhzAu72EaHKORipTR63cKdu
6RffObBYqXkWXveMeRDZx6ojLxXJ9AxgiD7u7TEnyDmjHRhMIJtjuVT32skWCLIHRUjNJCWTzOhV
QTZ41fDwOv8mcJaI9DskGvFJsRygOxZTxAUpx1KTZVrdWyX2EYxM9MRndKLBXIA43m4EtmQCcVEc
+l9s18PzrK6lEk1Hub/F/viza2yJC5hC0qFeaKurNxNn2pYTYbW/WxHvGFK6Y5SKkV5ry9Yn0zty
PrjZzTfvnYXGa63Nmldke1bAsY7Hm17SLk/VLJHr5Oi3xE4jlBoLbyZ4BmA+MjmQeTw9tLNmHFyU
z8aChjO/g1HneMDqWr5pV3JQ53F57B5LdmY/UvSwwqfJhUNlumxI1X1Y+juE+wMhOyTmHOW4lDG7
mT8lGaCpN0JVk3DVQgF36mhrcWEw1voFSaskODeCPsvxc3OFsgHno03s4mBBq+hUPYzqh3+d/zgg
esHSlatJdAqOPpQnn6cicaPVurg79HeaYhMRThvfJ08gZggrbKvba/wXLUheYDkbmfWetMFEJ7Wy
fnyiD8j1FVCLDHYSmtwgo2mdZbjrszESSjQ4fM2GBd7TrNFehPwuyPRMJtjzXjhUkm/wMPEt0iml
Y2IuRxM+a/ezakRz2/sG2F3DntE8wk+lNH21zyue84zq4biJlRvihg5PSZF0HZaZt/PMVhUmyECF
+4c1ly7uwwpro9A3u2Z19Cxr/OPBTTpf7rjE4uN4/X/pyDChOoxJFSc02ilv/ZoUATy0c7yi6laP
l/JjAUTa3xEpcZzkabDBpkNlgTrhlmD6OB+3PTLG+6aZ+5wr0UZuQIZlLdX4I0p7aQFOYAWtw4V3
Q64Ja4FBpJDJyFZSGJaq3x6Lgjaw2qTduqlxHjn69l3CpeJ9eu/d3dyWwt6rjAk+14nuO8DhhWOw
lADSOLUOFLn1vG745NbcZjUCATnprDt8g/ymVCtEjO92wu6Uvb3LqS9h85OzhijuC5dDD0Bz4X2I
KSx0U/ce6OvYoOLg2Z9KO24erZZicXV59lzOFITL19OcJG2ERxMiI4xIFAK5vm15IUvVhzY1CQxd
sH5MFpV1H9QxUyeQGH0t5EXUizRiXrgdsrAVuXuAhAxAAZt+ei2Sk2VDC0HQawcy9thIhPLLuSyA
oCweTgwC3pr/Ia35scFPktCW+mzYwjJNFaURq5+mg6FEbnJr/I/pz/jw5IeON2lCT535EVRQo4nE
FCrK7sJm2obrO/t6uKMLBnWJRxnmL/+2aCTFnLpjy9KXL5V7f4A2x77EFJn20DYcH36hm8glY3Io
bVsTjEiM+oOONNxgFZWt5x7UTqqH5x0vHAdIhf0r/mcgmRPipKGxxMdlvDZPnVGR9Cms9/ib31Sr
0Fh0hl+kI/DMSxW7BafWWZenLdo9WvBMpyrQRhDXwUg8LQuqawXYU3Z3ExovE5GrGik2hE2xSQtd
qb9heFJ/MFHMBDRYe67pPj5Qe+kbesH3mTrVaHEh8BBEFUl11NCoREuQ1bSjydoRUfrwYXJLMj+n
2ATzRyCT/PIBDqSfiG1EHe3YdEj5aHLFGkbzElPr/QeZi1CE6elGCYBUhOrfPOZ+sSYFEjHrxtNr
LYhiKNCfQGpopcuzWwzRI1+65M2jrPUwDC3B87UwrcD495xNHGxej9WEa5LtG6Mr3SO8TJPH0AQY
N7Ap8uqmo4sG2Wd9YPQ5J0jYs+uBe9dYP36NBVC/Xb7ErwBcwyJM74Q164QszeEhCk7s8M/LoI1a
s0fEJF+YtTQUVQRhiT4HUPdT1NFEnsS4of3Sko/Hwq5pczSBGy8Bf7HL9ZtGrjRvVGCBxMnkSDI2
VILd2ApQuX7xLBKC64bMXY0Kn6WwWWASQrI1fE4A2PQeZX3zI6UrYxLkqJw4gnF6xmnZmNYPq2xB
5sfmteehSrMHQi8uzVIrPmSGQlPfam9EBUcyGmYKJBkHpprb0mqao/Bm1kKKtBtjMGsYCWF62T3M
3D8w89YYEDNdvgj7+oxQmZP26NrFhC1UwIXhnXuZpRDGOhUyV777YN2FUl72nMIxJsIAq4HWVLnr
+fndkRSLmBVle9RcAhD4PuO8IGWdn3tlji3s/HvUtj68MuwW02wsFnPA9cIdvxHoK3+4Y5Uf+W/b
wUXCBwcuPymJXHAudCsGePRqhivI7pyfDRm2YfTeSh/1rews947InHW3FWfiSD7zOcPIcN2x7CgD
KcF9h+On99EpajCfn8mp+pMx2q2NFusC1AxfMudkAVihm4sg299YdahGIhepohvFcuiuEL18OVRF
5D/7KluXGOxjrHeTtsd3KzELGwxzzSwN4JllKNbGfxFsnF//ijm9E9Eu1N0FUtiK/oj1QhIfjxrd
ZBAVoQtIFWNAqsWbcoZX+Xbudu6OjHOTvsZNkDZVxSIJKta7DRPftBRT0sg+zdKeeMwqyt2fluEA
2Ts8X1ppBMgPvuJxL1WrPHK4OA66K0hLp3ebygi+PRbK77BgS4eZ8/eWmgXglRpK2YnG4ewQKbwk
CfDk4o1XNZwhJJvCNqKDx8ZfHX6/57hOepXDqBIjCblq3AEksuLILR+Kd45/caYLUWo4j9jD3hzb
2AryKUxRZgWQXi/IoQ4IR9OIrECAjaYhUPCZFAeJxjNRBPyMzR/JgecrTj8iItOT+WmcB6NP3O3R
m8BCM7vEl/8c7UD89rPLMG57CQp+zi9jsMr4ROrXqcSGs2hgZBzk2mhTkqsACGS4mSTWOLMgrTa+
KTEsQaQAm+0T+Tn1I29pKj9JKSU/WiTcomXdlgM4cCBFuKclSmYzIQsuo6SUHO9zwC9DGLHWQKRr
7qZnDpj9n+bR2TZ9ZwKS9Fal7RYUT6tsRjlqTypGFcIZqezCbiuiTM+Pz0vXh+Gu9m8GcnDvioKu
rMa3WYKFZByaY7JtoKC12r7eFztzDAa0eHlBK7IEHIPkup8yhHO+BVtJPB6gHhuPDtjUVhox3+a/
HA7gsYPf2h4AP3CW/RWe5m/nQIWRjOcANnNVVwBkAsb+407ajXtVV1LNs+6Zq/JteNw3P1oT6EHs
11Nk7Zf2ZsRfmOkNVCixyVUzAU4Nh9lRrLyTf8olmO7ulYWTuzxbNuR5luVM1+BrP52Ynexs/c4g
t+RnNV7Rv2iMfupR/srp0vS6JJfg5OX/Vm714eHGpUbHtmyLQTJBUUON503XokkDagPiMEltZlYE
kjW1SbrwEE83hgNCi3e9WX93U4wqe6Qtt+24KU+fIPswYqDrbD+Bf+rhqqhZDTAEw9GIbVHP/jk3
ZMZGjQ/Apa1+iGmBC6tyWTT7tTkXeE8fZTi/CIkni1zvVyh2Ngb9eC4Q3+hgCPUkuoi9IONAApJq
ZsIKyL0MhJ8MaZnFpX3dCjDjrjCpe+Rlwcuhg0gu8o8PnTn0UWyaNHJE+y1Sx15yQYn9LACpb6oN
k2ZnpfGAx4Fxv+hX5LZHhv90Dhuoqr8MdZ0AHPgc3BMykoPElmICNmn4HP0xpl/71noPtO1wnjoa
PJNlPaA6Z+p1R2/vGRsRffZs9HaIqamqyjHryGRvcxYpRyQfSt2eWvnmwre5N/gK6IOvz4mm/xGd
Kzh2Gzuh6f2lxXAYLQ+tbQT18QDxpbiZqNxp2q2LKOo2NosyWr47FhIzyEQr1fHBpvthC/Y7YJtx
hEC6FwfXOnpS0PrGQnvqrWcr2RYlEIgtzw4hxWpF+YbwPADuSUy1Yup92J3XXIcaqf0l7TwxXGIe
9lxLb+ycFw/64CN+fIa75SQpWs0ztYHc0xUgb/WeytYW0Qne8I7wCTZeuYZxKTNtXwdfb4clJNRF
Oq2JYGiMnXWVvY5UigpATY+1V0nA4XcrbfJEDBTL92iquMpbykzoUEs5Vu+wDQTtWNUyKwpSrROX
y6J2/RplL36EYvzX2zmQq4x4pGa03bJ42NEiaPKrL4Ebub2x/jBuGnolIR7p843xSA7N+tIcnnNa
30bKGaTuK1L4KpmcUW3dQuR0UVJNLBxZjuUGT0quWiWtdmtyhE3/2/ryU3s1YXT3Ig9eQds9Vnug
QjzlRxgHwDtOYDeS+U8v+GC7uU9wr4kWmCXrf3hGxodeqtFabMRGXgAFCan6zNKqZ7mKPBiZCogH
knxgoZ6QmBwj9Ufbz8yNziPknrULnbXUtVt5vc1Y6ONlpqR6ymwckY01f4xntQL0c+NEyxQQ0/Tx
ehsY9B1p2//Uyg26/aE7cYR3+hADjZo9Cym64kVIjHUpUwSgRScjMBmOXYjXn/rt+Ik+r3o/Uzar
axWe4MVVCKhPRyTvYg05g9Xa5Li/Pab5C2iPlt0JSl1Jejx3PmnqUKw2UOVfD0fjpiWDd7uOPmqb
wYFPX/bKhRtvIkAV7Ecyiy0QUKMJRzTMcgTemmy3egwSmATJporEyxy3DFe30RG7a5SFGSVrM+XD
n6lcAhcV8jHSzVDN8MTWPeCJnIGCPdf7n6oSkFTWDQ+QMjvuSCI+siWx+YKUY9ceAYlsbpwRaMWp
xRFohptQ+oAjKcoT5yp1RPaWJLmeF8FHizPlqPnHA9G+eIH4eJ6xZlJzISYbYH14yD0idS0RNX7Z
Le0Is4kvVMU+TlxLw8Tm/Jm+ieVlOizdEA3WaNPZKu2MCkRX5UvwFJ3xgEeeaHqWULznk/5jR+Mv
KFJk6bRO2MMEgpKtGdwt7v/mdRVKbP/QyC0oZN+ApfC5V8qy9QZSLc1JGE+4KNH14rCncD7VLLxd
7/23Zw9wV+ANOLmejfYBcekwxQOW4dUkIBmRXuu4+oHM3P4WnBilovCA63sGMUL+vk51GHefiT7B
5d+nFsWkBc3EHkkS5MK5bBMXoPeTy6jW+Vdv28/MoV35oR/62SM4ArKO8LxkEl8MZUHF6nFf05U8
JqUccjlxsOh/NzMwftTMjgUM/cYt2VCElX6yJnWmvsXbGs37+fKIJna7uZE5pZ43FPwqO4lkgkZg
KeTUNM0nFPT5VEJ86Y2iJpt84wM+3FJdJi3Co7ZTinkb65fH8Ja5HTZ+A77rjjOlye6KdjbxlfDl
UQzAVCCbqVTo/Ved12pPBQAgKxVRwFOkPyiQ2wjzyN5YGfdLZUeajunP6FOGrvGNEehTNYIhLMu9
Kd4gbeEAsaNsmwTCwGa1JDA/77y51hUTE6SNLxlz1iFVkDeRZRz5JmFGsHlKWE7sPQozl9HnL3wb
2FASa4ZPmmcQqklgKNNa9l6kv9hDS7bVqpAeqcZpWOqG/2rjCUkVpNaObTFZJr1YLVVpRpE+uciF
ZWOnBq26SnSm6h0tE5nPYmYI7ci0UL5YpTYiQw/lhIgOI6P2AgNOnIPJhLsoJo3SxnI3vGcNyig4
nmk8SQvp4pFb1SDzKx1PNOclUYA+Fk5v+/IEkfsRuQubU15MWAoun0ZytV3qqwscUZyOGOsJxkSc
v7YZc4ovFezWL08fHicdJpu+K2FlDH9LPCll8QuHsQQR3KFWxxdVHWMAOeIGi/ark+vxFN81yTRE
eZ94yJTxCw/P4IjfqvtCJQAtMKU4KKIATKkaR7/Wet+0i5ZFVJ8hmRfoChiFJClGxZ13ILgStgaN
bWZsJ/3obsvwuOnhE4yVlFn22yDvFfDS2ho/YYcghC6gg92otd61FSiyhzNcmH6xXkeZcDbn6EcI
1DX5dNAX7I/T0p+n3fnZmvzRBt/aad4BTiqEI9AW/Vrk/rNzY2YffupPjyywggbYzbqlKoWnHqJO
OiQdf2f0RjWXsIJD6QVfFapE2vsASFn4lmZiAlZ6wM3t1w8dtBqb8f1qySB8s3We66UtgN8jQB7l
iQlDtunZlqpzZEfhppNr33QVxIrpNqBA/N5JeZuq9vGgSA/YxjERVUCINGNkXececHOU9O3i2ys+
/nvQ7WEglbOUkgYnDBrVDUYLxgpdEfnzPheyO7RxeY4FWhYDjbe4arsEDvHyrrCQexxjR3ouMNBH
ReEdKMkyC9amM10nVvWYeJrRR5invNdT4/I4vBqPIXen6XM/hzhFE0GKBGGes973TkEgQAjNqxrV
aC76JA7wnENlu+gHdrbSwcfRZizk6fEJSUk+w9j4M+zA1Sq6CPbnXCmrDmDrAGtioe+qVTl4j1Lz
JiJH8ImCUDf1M+PnPCyZynbKJ4y/vwFJ/kIKGCHbCPn2CQs1gKGyCcpaLJt4miCZT6E5Ihq4YAQK
3M0GLjdI9NqMwJhtLv75TWK/K7/CTGDBORT4WFCp9yFXc1LXDL+emFfwSsExO++W3bE68UNBI/HN
V3iPUnGglWkWOXfHuPdJK6gE3gkz3NqGcFpp3ulW5tQ2P3GTZzZgy0hx+vlepml+gEMbSjtvFAS+
c411u6JW9fI9cjH4+rERjsDLvBsuwC3NgRfGtx9nB0lYztwy54TcRxiKhWci2kbnRKTdtcivqi0b
heEDTZL0kPJTUJytO00h2npb6jZ/SvHRebBnL94WahVo0c+XE44+3Ole5McTNp34/2/ytTPlHKf1
humnew/M/KgrDcvbW9sPdYf5B8m5Vc9YObz/0/xWcVEp5WMFTxeLL1Y8tEtSyCfZL9jXXhzAuqL8
VQpRxqBWF3sED0D0UMAwglnjeL5Pw+kDPQnZz1QRsS9YaUwvpiU0kPlkKwbJjhtUZ4WugIoHJVkQ
EvD9unwQRqQ0EvPCQVmDA4s9/aSM6Hk0Fb+vWio/AtfRxYsGd90PWWlqOGX16+BK2+9bGIDUu1w4
bnXdsi28vNPgv7sH5em12PpJ+9OqDBzuFk1Ey/HQqYSvu8uCdAVxoTsTtLucgaUAopjx+9e12IHO
areFhg4Vp8nxatAXE9m+/pnfphF2HkGspKcHQEwMwkFickhKQByWJmVudaLjYGbMw3ePLvkjs2y0
9JvOQqQ1Zxm74PfeLId0gBbEDkZpzcke9EKcjO5n/lCbuQhUbJQn9UZKQryesXoyF6C0Nid1MANy
X0c6jPYxp4I+IBTynvO2fw1MXsNuFtohPJtvr1iH+m83lHiRY3MUmgNxoSZDEHckQKywAJH9hX/N
YYxLhqAUMiL38t3py5AcQF+ty9hafh5Ft2Tm/E2gnBjaMh49BQm6VQh/jjv86UrND+2jqByASudw
TY8z0banxeLFrEUfXlApJReuqMTj0nNQLkoYn7NFUHLLAU/+ek/ZTWdkMFo/6G3HAjq3PL+9aM04
rYCc1LEbMdHbQEHzCJ5HR3keuU2pka/cNPxDz5LE0mFz1KcS4E29lrT9cYxKpJZqfpi7EdaPlNGk
H/p5HLqcH90E79ddH396CRXjf0jvspIpsKBd2Be24GAJRS9u3Ke79Vav3eBCx2Lf1pijNITMNECS
6xFiWpnQCycU9UUAmiXhSRjVjztFRSRaSXUEYZU/vniiQwPP5hG0Wo0cEmkx21sJUhKJqz9Wek+r
toBDHcpthlxf4lbTV17/rPIks34TxFfh8uQFKiUjnRjbdIB5SXp9nJ90QkBcgRBDXBu/llGeFh4A
X/smSBf20Ud4wKZHXtSgSqM0lUFragdmCeRlL8PAVXTzPaZPMwInZxtqeElFE2I7uuxmwclJJsaf
Ei+tA8aBC/VTKtBjIcTmyU4dIQLO60Gr6R9TmFxnjjmXOpHMI3l4bVXBCYDeOH+KB5Oj4PifW4t4
ThgweXBZKzpUMghPdu090MYFqM9y2pZmmZCmFrurxMyxV/38u557kgroOAsu9LCFN0jUnbAQZq2/
NwQK0OzgUFAVg3ye7V+8h/NaJn9RRSkjRh8DYxndNy6AR9mR9upRJIktWc5Jlx5TlFnB7Ogw8XRX
dYJCl8MZop5LBW0ZOhENsM7hoRpoeIVdyIpQNpsme498G2zt4T4TJis9S1jQnABhqQTgwf6MizBj
iFtks7tXYHLWFVKz56zQLNTffsAOwlWzWEiuvb8xRdc5Ll7yurvBrj+kDTclxBSDjNJmwnvDH1lk
jPhGNy52Dp0wWU+SVK0setSX9QwPgBaTwxXvxiaGEE/pgQ4vy3dcTZ5OhXMuVFLkcwJVr0m3EfoA
3rXd837fpFP80c/FgaWyS+DZx9S5F8CiQTOeyYBiup5CxUa5NtV47bZnKiSY/NR2urjQGcCuBBqT
M/Cw+t2lZJEATtXbfxjadj4Y658PS3AxkEo2NtVr13Pjmjlu2Iq9FLlewlGgNm2nZFD5VGz/wjz5
XuABr5xEUM8A1z9lsdEhuTsv986u1iu3h8E0aGn3EPeIJ1rjaqEfTOSdZR20I4ejQQXyGlCv8502
EzpOoE3u4oNv1+4Y7yfp1hg8wXDN16T2nwWA7ApP6DxuW8fkX+QEBJiITqF5qQPFnIC3Ms4tWx23
UPtutJhGa2T2U3eOFZr7e0FzVYpAszCN9qa/RJGepR6MuJpxAJzu/4i64xCF1aGbFwImZ9H4TTm4
Hzeb3prFJMqLWo4cpq/xU2ZAAHiJJ06h0HuJUY7yPjVie0nQe8DwXC2k+4xXmPZdT+vseZne/nnq
bcQCui6eyHaOrNW4k0hD5TztDvO90+R+FODD8FV9HJvHGgtyJcLTYclHFZlSlsvAFw1cgnSUSaw1
1dvrAALZ3BXO5+nvGEh6yhwbBMUetyedN+VueDW0aAcDIKklV3pZ4G9a2GDcZz5arG6IVeMmsDEC
db9PTcE2udPqxUMsTlcPGgrH0HFTiNKFvqBeouANtPHDbYECM9o4SDRS9pwZEf5sW1whO0cPf6Ot
1KmxpEyfrhAAdzEgq+CHOT/AyE6oCNIwURL9nskejZwMv9m0u2giAlChMPQLnkCWX/DQz5RiMm9Q
ooSsSqpUX/FRPfXLDEUfT65bVvYs9PAYWmSJxmtuNnY5ZIhAfAQsibQI636D77axkfQMRHk5gQ16
Byx3U1bOhLmtu5l9wHpkNJ0vZjO/+9JjQkFCDoRtQJGVBbRJ7wWnGKnxZdvEANBXhFQp4dRmV2VN
Npl49TZdEGETuyO6s4svP2Xd9zJwEOuF0K7WdwwZNxOgEXOjlUkto8JOOx6TP8s9nH2Xyaow1yRK
pI87Xu0rWApt7BT3kJmZIQL46vlk44cHHmV5E6dt8swjfuXsqmMd91o4dpopPPh1zbi0VrsGzT10
gzZce82egaLuEDP2JshazCBcj6ImFBwovWAHkLm1vWeLfJgf6UXFqmxhOtRQdnqYOPS/6dB8qSnq
7A/aEdy8ujIyLaASqpTSnD5+PopX5ZM2ENu9ijT2xzMxbgLhBoHqgvV0Gjn094zrC/WnscYd/9Ib
XO2FpjBqI97SOgimatPREOqOIpX/7tlT+kPlL3oRzjslTb5CHWhZelgZeCYlu2lvD4QL7KoHCeze
RNlpweYKMv9uu9hKyoM428WTAoSV/nnpMxpOWzPyXCwRPysEr7iz4xhw+r2QQdPnJ4qYZ+Od5P0l
yazU1ARDUa6zX/bQtUWeIkeXn3KDZRZKjOi5Ju9ZRIYa/gY9ljobqEpvBvuWq5ZPETKotYZjPvMC
eTPIg1z+I+8X1/heFmxkLKCMHfaTnvyvjq7ji+NAK/17CZfxzhDvveQpanddGH1XQe7ZuhN1pH4b
NK4WeXmC79NJpdy6vXaNbDAr56pm3FK4schLUKNDH3km1r83YcpV5cJfYh5dlLZor6D0000ZUZRs
ZnLYBLTWK4P5catn5Up9mt+wxyEQfE6OXzemBOpCNyFDwgOwMGw1GinroBS7Uo63VmJp1Tnu6+0k
4ObW/OSCN49i2oaVXEyPG6rh6/H0ly/rY47IExZZav4P4rTtIyzF69WBk3kv0XpdN06DzCWqu2/8
HbZoqAeDoy8iuh7G5ruMREn7+5K7WAfb8jtZdnBZuVprP3N0uCV5AyR5L/y7LXG4Lu1YmBmDoPqu
yaXQrBWo2ub7rl2EcEJDuifXoEH8TTfhFDlWLrlouu2PWnuzhjTy/m9VM5DBqgQ0ktSArowtdybl
V+r2FIlwq4wbbIgyGwYDILZVUn1/+Wfo7R3ZWJryZl428YcX0lOsxz26JVb/gyZeU6PF/K0FRWVZ
F5Dil0gJILK9/jN3ztKQ2J8kOKlCA5IUAmUULd0UNAEUlMZRpakGNP4I5cfij9fHn7ZxdrkjQODQ
zvbcGLC8/RxJtBTUyUmCQ4yFZksmK4ARAPWLGs/bQdKMPrhx5nptkCLfAejL5iLw5rn9zNc76Dwr
6HrFysGI1mZEsEhJIH2zvb54p/oLoKZbrOH9+hneYnrR7MJ6W3ghE5j9DB5sNBmoJq1vB5lC271u
Vwbflijh8jugiHWKjSO2io/eZIJ9eLICFYZOqH57/cy3YphYqWSYWtRmoJACyt+FmonFM3+PD2/P
xE8IPe1S5sBPRklae93QbEkATHdgOdl2hGpWEGY2xbsndGNMOaIpv32aN2Zc+6Y/RsyoL/sdv9e6
qfZftEfccdh4Gtd9RR8FIwlDRgdhyvrkEproG7BDzXc7f1hZyw8Fr9WP+n8mVI1qrVGWg/YqX0hp
JMniYFNOXZPdtzHL2rddXummy5vgDoj7orfOrbgwt8M9B24Q0hys23rBKZt9NMWyTZASgkuxnOsb
caWe7OWPs7gBZp6wwkQab5Crnzj+L5cUdFcgZ91np7P5Txpoe4E9xjE2D5z3HaVte3tPCBzMq1qq
ve3m8sL1TJSjBZx1AWWlQT05/zfSTs2/Gztg9CpGOCL2v/66LmcZg3Wvk/6xxCa+mLJpHzYJg/Wv
nok8kb91EbA294waP3ZKon5cQxeq+I38H/TF8nhIj5pc4Lff76wMcwE4N3efAsn6JvWRYVak3Qr0
x96NKtK+bTGNHEOjmHytk6AdwVWZ6XZHzCq5bcpU8rXkZSAydwIjKa4YJmXOvaalEt+UesI8D6ON
ruHYDCf9OpxPEi88/IpE8mmeanqS1n/IoLIyYTcwoWHLmieGlt6BcnJ/xgrvT26ZImEsc4VS7Y5s
CrARWI0Wdy5sWe/l2Lbl3FgBXBVsTW/RqusYGHIA4dUbMHrRmVzGfUaxNat+KwMaZmcGMR32HY4g
o6eUe+4xdI1v5rSg1X0XyXh8omF3Q5ohox1vhdWzTK6NdP1sbiTfh54y1P4/nm0frrutLGlh1wTZ
C3SdQYNvSW3RAlZz2957N70aG4xh0Ual9ojYT8oQi42/pZekb0XjlxM8Uw3iRzveeSbYdhBfzbmW
x2BRI5teMSrLBcQ1au0qEtkAO/qh5HSTzLZ3GUHodDqytzieiZ3NqHmOf9LR73/1QBlISVxDDGIN
AN8UqklVnSJMqBXQ4z1KACQqDKz97S+4MWCjDys7zh2Fmsa6n0oq8h36RnUFPnXJY9ZG8s0Qh7r6
D/BldIEXZOwWlFVo+hBwS59gHnboPttD7abLQm+iznuyucZ7X2T6eFj1DS5tgvEs06ZboduTKCCH
WpTwkLF6COwi+gqKGNj6H74anACgCxidWj+7i6YdQvdzZjhC3cIf+G/qtvea9NlPQaHC/k14BbBf
APF59El/danqeMhLoKqX6/fcJ2eB82UlG1gQ38aAS0qvDXBZCwQTRwIGiiBZqiKgKg1whF1mMPib
Rk/xqyP7x0ANxyN25vZJ80W4MsWTP0+VwmKASQLFXWoFT8uqc1yXf0c9lZyZeVO4dYgiQsNUJqbB
jknMqKmiRv/FRkEfnL4F0hUC/XTWhjNv3NqeDY2XlVbjz+NIxTtnbRUTRtx8gtN15TvGTmOcrWhX
EF8yCjgH5kJKJHGe0+HHoixj8103annKCJ4dKi68nfYeCO4G+/fXs6vFtCOGOwPPTg3tc0bCwGnm
UU0b5x2tRkQfDhBL5HfX55WHOUnRSWWT8cNjZkMM6gDyHT+W33TCJXwasFJbVMzHZBAo+t2hn8LC
XdWFYkqxUInn8t6eBGYan8bmOPMNYDuNmX1vO3sMZ5clF1NHvxLwGlR6V41+4x1V8iU7heGGwvWD
b5IsFE46DICRAl5uUkF6wVmtBTCDT4ZLf0EkC7pajIAks4H/XxOhLlWE2XJScmHrsgFbvNpNinom
YMHHTukUBrAIJQ8OLyFQkW1TVQ1N0zYErzJKSdMUBIRVh7Flr3BsZA8YK9dsrNRqVTfBr7BHxiet
wHLWzdZD5Pvkf5r98aLNi3XLUK6p0g0NL3Pey+N24LjISKYZQq65Q4uhcBUMNi6kcs9hyL8uSMp0
/GGOnsYkMwWsAepJPC4aXaGy0ySHOj8avtdwa/qyFezPQMuyzFysrGfbkkuEGite31JPSy1Lweef
9R5ZdNoRMg3nSsceRl0+DgpgDpoJqJKexBhzlOW0LvbCuYhk5L7GTJQx1HzSErMXRzSyx+TtWN0+
bQG6rKqScvVx4GuVQ4ZqqLcXPfyIzF/Z2cHdySXlBcO2Im3L56m4SKOlGaFWqcnOLQkaiB93gxHn
Xf7EY/CGbwW7zgXa7nmmf7tQfbXVKuhUr1IhrS0+XCimAqRQxUf6ewTydCOk8abj5bblXze1qjGh
+peFWfHRWDAhzbfWk+1mRx9mlOxxAN2mIgwi3PcHxPDYwpwVoLiJgDeKjwswmumsPDSMZhoX37JZ
tm7pYYOKGE6Wgq9iH7mFYZKDDn1rjip53ZStI3faefYQMDkt7a0YVly2cPpBJ+WIBAwrOXYpsAgr
rHDsDMldXOkwaJWtIA3nqixCx22Wqe4xiPRTrobqx82wTUe2g7WfC1dFp7j2a5Dh0x3/YpRfkSzG
jOKG7YbtGcjaWjjUPFVKdjEd5hBuqYm2yF5p6uOnVhNQqB1q/MBj6o2gnyMlPXJrqTa3pfzwGTtO
VYYW1hGTod5pB9QS8Tb7JJ9bOGjAP644iXf/aPi3rYcEP+N26O5lr31DYkhwZEAHnoXcUyf48Hu7
gMzjWX2VTwAGrDXCN04JKeSVcVG7YGqCAa2p5CzkJ6H2wuLcBF5cYk/nSntH7eNtjAM9ZLR5WhrF
GGf5YTz6cmALnlVsbYuzfM8118nujkSjRyNpwyHc2SBDp23Sx/dCO4jegwoDd19rWE2TAjPBTwXn
y+LdCXzWBpvgOEpbu8wdaA+VXwhPCn2fBu900RtC12zUybfA0jPvg97+ye4j/2F16eKjSeTmz8u7
j5qqaCo8wBlmLOmJV+PAhoF0ehwW4grIT+NFeix7tfaX5KFht48PZ4Sn7IsFsmy0YEVlvCMf59ao
gq3IDHaRQGzu+aywPXihoRHA5dudQX3cZ/DGs2NsVaqtcM7hdFPERP9WtNq23+avEiXMx7bhz2jG
MAq8iB9/jttAfrJpXNwxzj1QuzfbFPPPcFY9R3AdSbpNAmMbdbGiA3svcTCgXRFS4HOV8FHVjonM
rmpBclUAMSKmC5LtTBpaCDD8CEpu6pqTjUjLsRquFKJaImXc3ynmQBMKKXRlkNd5k4f6TyuHgFQC
ngcuXJ5Nj/aRR9rtTjAzy/bCXGEKGPqHxq6ginPP/nZlNRCA9bSBWq+AKaaPP07JfqEU2J8Kctu6
izmmB7HiN2beNWpUtmiec054rnt/t9/1YBZ2Rj68RKQTG5pHxljt4nGZIV7pAndemLnZho4wKkgh
P42zOmCmAeJWVTxhzWPiZzWlQWCCG+51/Unj5Fx5ClPf2GnJES7pMlu8QlV9QMFXaYyru7c92JUG
/ZgYsjjD5TujhqAYNu/xItt4bFwBrQ0H/Obp0bngMQI2BYuGJxh5EK1t4WMUsV+wViUXFirPKB8Z
87YkuZS4sqojHN7EAUzvd+OmWKQs7rvyBbZV8aHsC2FRseDJ4zSs9RO/JiqKQOQKI0bV3uB9cRRk
/1YJ6zor6D5zra6sDE5z0gVDgrsjs1Ta0mai6yYu9KI3H5fXSaeMqGwj4QgjxtzhahVU6sfMeJ8o
YQ+gIkkzVfsOXABHRNhzBuGAZhrFzJkTlAbIHgWPuNhQCpOcJCXjUz3p8lA6TcH9yAk8RMx1eHTU
2H6HPKOr/b6iUODDnHD9MUOMgaZK7bMT3MtJMk3ChPMknllvsOXEpkaXmdh614u2ATlvkYM5io/B
rB5yDvFg+zziTRrB1Z06Kx0bNDT3DPrMY2OQLw0UibkY5LAp/qq5c88We+V4Er7y6ZKw7l1PhcRb
mWKHO7SCiGsn2NOnqiAmdYJeIooir65mHsUxazxKdrP+5Ib+qgNxtnjSKsnRjFBl7gDV5wrN5YIi
VxijL7eoNo3Mqf7IuiisMZdJ1ukI+iL0m8r5Nn+Zv6IEuVABMeIMmg1HRoopkg5+EXX5Hu5SI72w
KTvf9MI3U4oDYH0MnZqusXbnZnr76mXhmo2EEVSGhhSvoyD3aJy68xFYwGhjaBdyrQh+lXq39dAP
CsdmvNsaoLvMp1EmQxYixOYVM0MDsWyBa8wk0BRpHl/snkn/XjgKmSYa29PiBH4mVR0ObXZ73DPU
ltBil7tAKVOidLQytN76rbhiyLXjgA7uBuf9BU5EP70S2K4NMq/5+NdoFWUGLzA+FlbM3/ocD+zv
9cBNNgF4Il7f7KSdqHMw5jipqpWh+NAgp5OZweMkS0Dt7qlFQ1of23rCqiUSmZpL5NyO7V0mok2N
riHG0SqOS4xGQYFsV7yf7QWkjt7C6sIbdmD7Nttm2U+gqa/NeGZZr6LxsLfvFvKNAQ/nl5SwBDTM
IS3SiKZ5hG37U+Y846m76u7pz/lS0kE+TqHAF+tcBO16jBqOnL5d5uSwZbwZlS1G51Y9gGscLTqe
dlDex49jOMKbp2ad5d93VTj40c/K/99iV/vgaVrGr2CwQ50zIgscoeIRKGh7T2Rj2X2mfoaJ89BZ
ZMLAQPFSYz1AgvlMfkKNKtsESI74lFp97RDn29AkN3svDJJAG3cozU071Rmu0haf9KiKyB1Fc9wP
m0ABdBAdr68TTsfhrc3/0mW8+LCVQNvuBwUSLwVW4n6vU7IOD07+JeTmSeo8H6IEsv+QL6rq/2fJ
DfVBUaHjhi4+Wlnh1rJPn124AfqFeQEEiC+uNWXzpvX5KyUEEMeT6N84g0RnWhrzS9ClsPxXFY+Y
VYsv978jz8CZj5g+BYZChdZFbXJXaE+X2hfml17zzAYbfMvWytBQSA9mpHmJKoErjdbKA99sNkPc
s1k2EHfQRbRGt1xO3WKfLcviLbv2TS6HT4NOMobtNDdxXpS7io+0JZgXMdVuaSNqMQhVv1g+vyfe
x4lc3Q7NpYnMONupWuFMLX46uvaS7OuryF+VHsoSuTUojeG+osKflQh0dq1vB+4KJw0JqUvtXt3s
BkNkKNH4QUftmCfF2d+NeP3nyaLDVHGBLxlLK36cT2IzCt0gr7CqP+hgi6CseMVhfv6abraizvCs
2CXQaNYwfAzs8BjQoxYhRIHdhN4eywvbCnA29hc/6VG02BdMzKEsm+2dv5ysTHwakD/D0+uBedFs
9mPijn5LSgO2UrvWRjAF+j2+SxCDTnoSgYOMG7cLagvyNaxzpBtAvXIx88xeOwpzXaebSXcu50rq
084xH+dqexAupOnYNLLgWMthJecuW+CkRQl81DjWmbXFpnaq7xWCcEe40ixtzS7egWIvuz0NoP+q
S5XdDpmA9wT15o7UCE/Jpik/GTkSzx0Mrex0Qf9GB6D7W3kh0F+oCGm2n/MAfOz2REs1nLireffI
CyXg5RwXL3NEsz6mWYIWeCq8opgT7EDbkRxDtHpdYjQGzDswgBI5kJgJo2xZ9pSA5pilAqq5FJbW
jOuV9n7hd2jIF026ujAMscmHgDZP/GCiBF0048hGASDycL0YvswPnT2iNQgXX9wbTCIsXEAwPLI8
xJipoR8XxL+vfxX6ukZvtt237vsDfMxUxO98eo486sNrvO1qn2luiGsctx1LdUk/dinzBEJBdjde
ghy9o3fbxWwzpSjzsmoEnAqwgMGVjI0q+AIISXVJKiMQoQAjhqgVUKqh0aNtxJGhnnQY4ky5YFhQ
Zo6usoAtEp6KPCxrVj0r3wSVV1uraHUCAf8A/fZ3x5yijZoyMu5LAB1KAtBdyJnSjJ5U0XcCb6VG
Tl7kZQnOvR7ijA0I6TtoLPL1lEQpPbYpwe/ilmA0uNlqLoPRJrU2NIS66H9F5VIwG+pnJcMfQuYu
wSts603C9Wnh5hIffy5rMu2e32yKnzloN/AGiMs5vcWnz2Ryd1wmQzLTrxgoTIDlMZwvO8XkLRZO
HifJXm0lzzsYvg3J3oJZL+K5zBCf7E2ZfS1RsCAriyVKiKSgyxf1VQvKfqlM4ZXZLEeQtIC5Bz0i
XxNGH9F0+dNe2GaMYTn9wynLenbPtT+MdK2dsUKRwzqblQTwqh3L7grXsBCnlYcFLYZQcSVKxiPl
ttPaOUrjs7ZPf7IdtqnUiCtLin0ccJTyywJZHQXRjJBDl8MfHEUeExrK+WacTU1lp69OZkR0VGJm
KrEkqbtnkltnesHT2GKXP/x+ih/IahKxzqPfldXn07uEpEwhM/BrMWY/mgsXSDSpKjng8hBJindk
GjUxj6nL7lYCQZxSBZC8IIpupqsLRY5bS3eVq2YFM04/uRyyHqvahws6UNv3B+dWPNhg9YnsULgu
IWrjIE5JXt4IxWCW+8ctkIMkuYW0Cj3MdueBwZX+b7VZ8h6i3pM8Oz5O1EZnjiMfgoM9Q2GtVMpS
a8VTp7/v3BA4JIyPLcA6hIcyrUZcglxtZ4FACrwn3GdWfvW1nakvUcETijNYk8rvXWldbHZb4KaY
5UcOr/AodBfe7zM/JsrFEHU9c+NMdfBn4jypoVgsuFiiKDLEowJ1cyVETwYTZnIUuS6sc6PkuL8V
Ml/k7xV2Gg3u3w2RczAnCFG2OTIJO2oE69O00bfWvRM5NWD50cUuMn76+iUGKN4++Ggy8NkisDk5
27/k07BokgZ9mayCARASw42Jv/BPVip0Ahq4t+vu52k4Ml/mCfbC6BWw5tQlaIs8GwMyNNXsegq0
CCcwqB7uD+07h2o/+cMIJR39cFNJa1zmtxr6V4rGpq1Q7ps19Mi43+aVXvzautnA3ZqXvtu50RFq
5U6G2mrPCz7Y9T8JhxnKVV1iDS23YDUwdhSIMllUhwGaHizztYxdHKM3OoJgtJfdU2y0Ur3BFdCq
KBT7hOqsl/huI96pIywxkEfP4TDemizjnhu7UoI7/HMsTJOf+nOnW7oljVo+wlobzImSGhYeu9n3
qaggLiOOxX249NwqwqSlaN9Ya8yZN73/fOp2paNrgq60fR6R0rpaD2I03j628U1b9JE7byN/ZbMZ
ieug97qqw1il2Ws0K37Q5FqcVDCNXC0o2/CADHWnnhsytOebX7aL0LIrXpZtai32QVk6QRE1gijL
KJto5/C628ptnohXrBFJ0zoQ3oj0/xezGCWlX4hq/yG9IM+/4l0IATrXDEmTSBqTRWRDYiI0P+/o
auPlg1FWCgVVIkxuOoDIzLS05g30L/5si86rzxz4mJBBIfF1xZJLmR7Pj1H7R0geAMUBhtGnyAl5
A6nFL7kE/DMGfZahzahQefyTKQZ4SGfqs9bbEwBdelebIbOYCK8HrGgKZz9C4qzf1TkgiGrSGADc
vAcxIxBaTVrJhh7+nQJwTu6jQXn+HrSCE+ohD9vzeL2LG8M6udMRv7aGI+8tV8E/7+zPGAQTuYNn
o2SA7HzhTY25C2weemAVjDnzUkyv9il5D2GeJ5pgPSSEywLQB+14oQNzf8GCbyEF1hcSCJv1Eh7E
9GFQT8JSQFWxcMD1WPEG4+vCi4scUw09tS2Z1Nt5np5sWjEInX82YYtO1k+xXppT2nuxwCwf8kAB
zvwrE4GfnU5fzw7/kOCDC0Uc1BGsYiDFJpXv/0lo/prJyuB1n2+FSzG5kv9Itnu4G82xbLz5uLMS
RZGXioBMCsxBTLDfrSeMk9qusHCgNX4vKZFuZ6ry5y8TGhZqlnTT0j+A/a8vVmB1ra7QE5OzoBvl
k2TewlYXK0EfvZcxgOXdNgury2T95pN9oSDraT0sbsh2iNtdGwROvX+jRpswMuC5Io9/OSa+of9X
t56//XTBzCTy0BQ55SoQsg27l1O7Ft4yLzf+uRMgr3mMcafjaLonuMOgMO7k4YDOjj5rVG1p8ccH
t5a1sv/CJC/i2xnDESScRDi8UT0tUqNbdCRI5pEylG6d1dknh7phhnLxaHgaWR1ZZPN2HstN+wAY
cxNmbUcT3dVbxKnBalUppieA3E0hoPB+9/ZIAM14dYeyNhIwHBVAa6g8bgJ0FVgIaqNx1WhIFMJJ
B//BKQzbn+Mlj/QeKgUyEJ+9GZYdqQXtaqtJDfMulS/4ilaZ6MsHb9k5dPv/tP1TBrLAYIMC7WjM
9/O6fhASW5+1rfI7EcBFC8USQKJbXsbR+Ju+LH+Wc9PBzblkvy15h0QZKjuF49tScwIzv1oGg0vj
gpYgp+JCsHtr2HdoHkDpDTSiESFegLjAstt7vf8qCYZrCxA09DK3u7orwJmD923uTCuBR4j+uJ2R
TZ/ZQZYWWMR3yu6lKdNHTXIrZbJlk3W7dkyPcv9YeaRDamyydNh3zswN2aEhE7ng0D+hJkCywBL5
2iy6t0naZ+M+Hm4gNlCIErezRuA/gFfpDbDR2KDwwlUKLvt00mCfOHgVd+nU6EuUszPPtQvc3BA+
ytGl7T8UfnBBI1lx+tREVQIct7pNNiywsDFbSVBO2TbYHtqGGVfdLLQhwQTobbCevZKK7muKG+yT
8hfB2EWL3i9Uuu710jR1YuIi/iQ1xFoyyfHE6ty9wVpoS3syocPco+Uexe18DCwj8GahpQ/CIY02
fZ29AMboWJUa6BUG87KVBKlrpQwvgaw/wnWLCkEgYCA7h7jXd2MZpzeawX16zH9ximcZ7wFaAvLp
CQ0eleEfIzRhUjcGwqZFI1lU7rjeDzvB6J/9bR+VOanQKaQJCbQOrEAnW5juHNubv3BhhIum0+dv
lM2l5L+wKFG4fbM6s9qkKm/AchhOWRG+uvjn1jiAFhKebAjLr959fMhHjLrioxCphAZ6fYVIpM6v
j88HoXGeNSzbndr+2q89/E8El72Sy3osgnJVtEjK/g8fX4th1U2AztLxgeNOKTfibBRZE4zfmfZe
wHJG2+o8aDeNqlJh7XMq1SWDLX6Biq2L/11Q+FErHsrQEQV2bv6rPrQgW4ofza58nPcYHv6lCxaD
055UadYvhDDfUd+BWCLwW8RXti2Bbk5kAzTKoBso/C69tQV2kRdczmz3+aiGR0RD9t/ZLALrAcYN
COyQo1i/hUtIxWoGRtnTKIzbS1cNj8KAlitLtMcDY5cmetYukZx3D2ZT1+YDN8/4t+qJDBWElwuF
SBBB715Bc19huse7Rkz3g5xlle7DPN6E4oP6PyDYMwl8V8M12pjukd69LwWT3ih53H9410VJfHYz
JlBxrmSladzXqEl89F9BvB/fblGbbSMwexHMzAVJpVPfaefcAAreURXXAnkT6uXLezi/U1geO+NW
1igP37BGx4uzwcWZ40u+YQdK3UgO6/jPweSrd6JIOohGQfkwpjs6qZ1BaEYlyGUxLNBdXKCC4Xi9
nmzJ2ciUmOlZNcpf3l9HMER3W4MxtonitDE4lSzVtC/sIDvr6SsieLfxz889soI4oBU/3M4dkN3X
8LxspIQwjOVLvxJeTqSspbE6aAqbRnhy2yYJP8aFs+eTg1kMcYE1fUy7TpkmVo6WJzdfhjZyUiWO
4Mqlw+EdjpWEMLJ89zO5YAadxLah/iUHhLcb118HVTHM8I2FMEGbZgPYl7+kWqDZw5pWw5WTlvNh
gRbLQj1e/zyqvpqaFACJ/dFTjaYTmW7p00jdisnG5xOM/02qAYd0cnqTC+js37KpxrvJ8WkoWahN
2BUHQkTecid6cTTfdSZuVVDAIov1874ef5VeNPvwsunPwCcRao6uc9VFOsTy7LtfK9HevbUeYSUl
jJvkVA+zq0BZvyl0po8TUv+9Gkk48bvMFtfULRROvUkOBkXTzsRywMngyQTkr6Q0YagARzr+gVvp
1aVwqzEI3NaEUYdU4Hpvpbopab82PT+B6jm41qtrwQQTNyWzAC9ORpm+y3NLOjfxKxYcWNXYqg3K
ZgsTCrtkdBel+MysfsnsghF2D1w8ScRqc6l6fupjEDFUZYxor+C/jSPmrkK7Fr6dAC4B0jY8mYEC
N/aSgIKwzwesgxuVPWQ/2jM0zxOKqnPwyuBrCi2OG6kxkQd2NDU56n5xX2n3wNgVkYheP2nnlLdM
P/VXkDRUGvdpio9MW72EVYfG0MkWqsQR41N4hn2Ze62yj6MnvjqWFYBadPWY0j2v051Ela7iJrx/
1mWE2piAacnttsQQnucCTX/c+iFpV7j5JVlyREszbjRKOakuvrN3PKW1JNx0BB5bY46//95L7zDK
bZczphOVfI+Bt3WNEAKB7ux2KydT5DxdqAi8mhSzx8fNmc8amASwexoyzl1J6T5kcMxyseYFnDZx
xNWYixJsD3e6YLe/CfebDDQaWUQssEsg1bUU7bHknTEvbhAjhGMQ2owJXRpZHo5WWkEHYNagjBpJ
nOJG3E7y+UGhcu+QO2hfnKzdPmBQyzwEMnefqvIcXwF8Y6kYTSjAvSCXY9C7TGFWmgad+lFXeUJ8
J/wj8Ol0lkSc1tNyqt8gSyXSDIlHYjCv0pz5aYp4Xxg43kZzvtuQk0R3IiyGbLI1/3nbeWcy2MHX
djDnAc1Ob2FKo5fUqKODq8w3cwW3uBKtdLQMLApml2XWTu72kCTBvCm6xaQPfC+EXU38el82fojc
yGou9QX9kmNRsLTnsj6enQ6/W/ISEGQdjf0NrKrp3RI0pxCNIbEj/h2h0DMO6/nryNFB0DBSyufu
gcFOtIbveC34njKvMed0ELunx0oqxTP3IrDRUKvoqaDTmM2ret1HnwFQXo+NqYyPf/23EF+kSiuR
Lrmel/c2vPcJiZtDsHNNfUzOZdkeMfZ5jIvxkadz4p53xFf2S8aX0x74slM74hyWy1/Z4fT3j0TR
fY3LrUDwJJsOrI/Hxm0tR9rxTYAjcSvZ3I8h6CYEEyFg5jccAWttj36mUOS+eTixqk9tL9WjkIWP
2N+GkowzG3+9/XtD6LZ9mn5OgHnCDPC54PMY15Jbjn+ha3pvJ7DSVkFWAGyzb6S0TtapnGFmICFM
tnSglulkpEwAGWggQiK/MyAPczPGrswbBfRLmlSsjIfnmJJDhEQHkwrNY7t2mf8R7NCgDccvadCf
YH3kAGALRXlqvGf5ma2a9OlRETAzM45I9KNgRZodkwoz3T2nCZKQpcVsoskI3UYxUIhB3woPZ72u
AtOBuKl/r4oPmn5GId5P1+W9xAX8gOuzqfwmhKSLdyqeZQxJnqIylECG7iVc4pJGdk4QTyP1FTCY
7fQpQCidxPr/Sj+9tl7mqBw+xHdqRtU8/PhcoyL70wVcFV2TFUR21TEmR0ztLo6EGjCwN/TmZHsP
gkJ5eo49P0XaFsvPI0/1nydFvcPQQluZ+5H7YWnfGIcxH74/QrNfS34RoxsPryYrJQZF0FYXNQ5u
UV1RHN2B5cMiSpRXxUJCboGaG2fOf2ZcanK/12+7+Y6Oe32gEZiO7zdy2SZLDtKz3oUZ4sEFoxmS
hL2XqGjAT7P+DpQGn4jkB9/2ndDYbLx933ZNMCUZj9QVH+UXu3qeoKLY3oZfVd0aXHTo9GviVudW
L5rhZ6EgcglXpt3ByM6ZZVlxXHeG0H4M1MM5Rm8ZPA6v83F43FS6jspEhfe68wN2//NkchR7EZ0H
8D124r3zXOQRWj8oqPfSXf6ih6VL8YN8knFwF1Sx9oFHJW1oM7kNXubjOAobPJqrgy0dVSpFsBmK
VEHsqKq3ItxzdIM5qIu4nf1rZH5KGubQ/ZQiDpSM7VDyiRuQO5B81Ij77Ejidf4Np2e5z2orQagZ
mr26zQNd0nI/8ue3JYl4DAhAyLDp6860Vkv2sPbTWLEY+5JiDZkF5MFiN0528o5nqMdo6ciTXG3B
wsX5dWjDk1C2GxEY38dBTLkrEM1gItaMVIbzCeEL+MGfUkEWVPu5/VtiocGLUaR8qCBITU2hWwWa
fbJpEkuY8+KGNebKga2M4oIw5ZCX+b5ngKsKnY7JuMCkjbEozx/I9BHLxeGk/0owi1QuS7AoJYR1
qFg2FeK3P9E+rzTUqL+S7cKICqaDZloL3N4ua4PSeeOOQDkQlhq4Kk5EWQmNhMfZ0nJio8EmXh+w
gBG17GsZHHuDp5pA7R7vrYIxDq0KvnTUcDMZxsI/lg6tMX/CE0H1tc6l2FbJH0f0/JtQIVQUwNTh
IY7nrMUiqWKliPdV1d7VtG5x4J2ZdDGifGmP21g7d/Zk3hI5BXiJp0aqr6IMQ70R38jsVD9TvOPU
+QXSMs1sHArcvT/Vv5BC4x1o9y9KznJBTNigik8fBIRht0DkL+VsFa676b7G6m8IqZtf4cjOdjbe
do6IzKtjJsc9c7mJrM2PI1e0En19IL37wYqS92M1Adp4/hTuJBLoo/pVd83Bn6l4wW0ZJ2IPFEkU
PXRKZBZwnVSQZGRCW72CKm6rUh6lZbEBwRgeJFlLPijORSBdlJ/FiTHs0LzxgJQs8jz5hewixr/o
iGlA5r6l0ZtSd49hjXzO4tqjSg80NEExu+Wie9Z1U4l26z7TGzob5Uwpo92dbDxl1K36T1bdS6g4
87TODm7BW5OUGHuKPqE0ujLTcMoC1gpLEneIybBtCJCTiS4DY9ydTgupEzjaY+kwQUN9euOZi/+1
/12RtmAkdsvN+vwd8KeM1JBsp43v9/An6uB0FSRThjBZOiAwghFCxVT2By1UMkI1o/ZIXnFz0hIP
RIkXEgSF0tJU1y/gHZJOQvJjJMHgX79Swr90o6axLD5R4YixGRPoTqZSJhYIL3pO4qAtj4EQ7k5S
Uc8ThQda4gtyVxPOMexQe87m5dedHRNeehL1NsmYYVBrwesIYdnHcsbSWR4UlUufAMGsos6+LySO
Ncz5TYtVR+OkMG7ZYMri7m5M2N37Xfz5jTvWcdNSXgeSddG+YdmkKZfZzwkazrcrsprx+44ouqdO
V7EO+6CQ/pcyjN8vVW8eizzQYNWO27jqZ73n6/je42OGOfhlm6oQdf8+ULQw0iCvmNXVe/d0A+Pv
EIqIq8TrWNSgb+Zu3gaNS+XXcQcIwmDFNbkiBDECwD8QF1A+6tu6TOCus8TkGIOsssUfdVD4ro0Y
PZk3FJu3Woe7NgLeaOGZN9bVCbDgXnk3ShtdsoXpr+gt4ZgohbNOmKuRZlE4gunSGrnmUo8tSvVm
3hdTsTSDv+iQPe41yMmgLSGjSbpOwR6I30YqMf2GLYgpFe7mtoKLe3DgU4OZiggXjhnCqi/+++lE
hp1uHB7KoXLQZK64GRYRQ+gTmW0LxQPi2Fy6kBwL1wpCuCjX4dVqGJ/EDcs8KPkH86SBcAEdxPs/
5srben9YSxUsQnpP87cDN/a2RoF+W6hEHwFvHzG1B1EXcoHRxo+A/qId6f/K6z/bkjZvapqR6MhK
CZj1wQsZ7K+trdYSoc1dAakSoigFARabiiaqnm6kY2RvFgBl3tgZo6ikwyeZH08U76n5W/fwPOCl
gwyw0srrNueMDxhK/WuVEZf9Ri9aZVIyDT9fqI0hFSUqCn3a71MZLZnH/7o31DEwWKeD7UsiOVD9
RLHQRXhvTsYSfrrXrvsQcBWcfowbttrHs2yj4Wz7WH3nVxBc95SSLYYfnJE70B+1xSQVjXRKe7V9
+nRqhLWbFLwMxJTiDw6HeVQ9M6VMs0JdDroYX88aBzCykrxeObrv1n2bMpAJmDhKufD7nvJTDzZd
/B4Tzy+HQ+akUUqpf90kIqbjd3619hBMTcqgBMEThAQ5SLsxhMgnDWBh5fZKr49CPDxb9STkjUhA
LP+STGMFXuZIQEbA9XY1n3Gupvu/+SAp/audjIz6NYJeNg0PsqGovD574US9IYzDr1oUCCgCOayB
Zb1S+Xbowsu2+Rea3+TNGumNMDG/IAPxSx4NQTbbMnAklqsEn6qsYNsp3v8Xj0KJvouzQlG83d7O
oTD9qfeEqF3hZg2vCVcxdLI7AktJ0IReP+juznEKtcixwheDTwSqYBCgl9SQjG9G4ovvnkD9QAv8
KkEfrKpaBuenoSRZVo7Wq800BGFaJiGSqJuNtR1TKZuY6uisI1RfYiuh+BycFXkDvh/95i4fdP93
vtdo2NpzFzjZ1oX4cC9mv8MrtqvZiS3mZuxMgiJMG0OLS5ok5XF1/y4AQ7qpUe3E+kdhjkb0Va7M
AKlBxc8uSQ0SFbN59zD4Lw4RzgbhDj/K+rZZ+YuWYFhHEoqOo+qvuEi9mvfYm+898vfNLR5A4Ggs
7mz1mbooCRewaZ4B3t7rafSEvCBDzjjYI9ABYz9fbW2kRVw38EPQMlUSlJ7P2o7hqsdring2V+mR
3rqF+h7iuPDbTLcu4qltOMYrb5qGUYH5x1uZl2XPtSndQ7Ovgbp9CmIbVPyfUwh/jNvg4YVkd/mf
SQ9gvN0P5QHHomzEzmYKFYjO4yQ5ppqXN0By18u6D4lrhLugCv5T39Pb6qkWsVdHmtQ2U11kTVCU
NuxuuNCi69FxKrZR/Iy/Al/4vfznxjFG/xhv+KMTu7NXuKKe21BGT9QIzKCR6S9JWXWqRUhP4Ukj
aZRM3b5UV4Xpg5chwwVUBVGZQz5nvrtWXd3RdBu3Qa8e/hYxFcDXuxx20bfM5+4d1Z6p7+MxxOt8
XXf2pf1NCO5jYaoKZ4HTvQyoQyt2CBp/y8Z2fld41a9mwirOb9r5w0LH9WGHm3ckFwfmJWk9btL+
J8MB+vmkzVJufOuQe6YfsdpDk/6UxJTbrztPpu9gIstIvbyBu70IM9rPO6Tal3+zJbfgTv49u/sO
NYW75P+32xMKe0MOJRQtZvaKV7fGwgqKXfIXsWnI1urx+ofoMgsrY+krtzwiTjlhatgmd9LEX2Qk
19dVUcMkBs9vuJepx2EcduAXHtrzrUcTp0tNnaY6EQGI9ya/qtKCdgfG/kKFzrjHoABSFOuFiWPe
0+COulkfafgLH4bakJBAhedqbugub433glSATnrcBrddtsSgEAPaSX9KfhumD3hGXFngsfk7TCRw
iLlTzvCgHQ1PF1XTDQlIEIU61V7tsbA8R8HGRydvr43zuxFcFuEcxMHdiONgg7IkA0I8kg464Ljx
FYZayAxpetvteaYKCIKc0fDcz0R/usBcixc83BYJJq2U08Vru0D382YcfzTL3yhwMkiblqVWrWgX
94pTxbQoUiACWl9hqxsOh+a2E+vlfmHMek+NflbK2jgcsf3BUmUwte2lLdREkWyNNc5sUX7CIbz7
qlEXNjbkqI8HNvtNeAsdMqUSqRt09nH2BaqNAh0RIiaflVRrH4qPwg5/2ukLmoZ53FPlt356KOAB
fA87SpUg4iNasV/MONWJ3RUP+agOk9l0wDLthR4K0fsJS/4pqfuO0fzsZLJmCtTms8ONi9uqFg3z
wFbqb4mHMWZnjac2Imla1XW6E5Jo8tAt2G2XkSLHFVHBp9N1fyiXQvm8hBR69O0sqPkiKYlPMLwY
BI6Mf8mrfe0Q5lapd2a6HrTlSR4B57SduPOImzm+vdj577qF9kBLepzLOSDO9IbyNltIgGCZn5ms
WARjfhmqwdJJuN7tgoo/G8Qb6dKEcH2w2xiGYG8wFW3K9VihCOJuydwI4YWrn2BiHyC4m9tiLEkg
RKji8EVZ0W9zml9b3XCClDA/2qm47O1JleN1ZkUczMlBMkz1gtLngYP4VvhvOV/crNnoqktdiNSJ
WHTaF309TuI4bV61WWmWhDZZSM/1XaP+L5Lby+JIKAtrJnybF43m2TjPTEHDoxEP4JgNXetrEtrd
gVGtuea5TAWEgZcKuyFzqwlSTnTf3o2C7zKDDaOfMWc2gljYK3YK8E+pgl+PbL0EdjDqscWvoifw
lrxywvr5EHx6Su8FIfOijlGo/Prx87ZwxtVez3oBwFhqbp8SSS01nSlOwnDEohzO6ppGrl/MT6kZ
dhhsSKtx3d2N9FA5N7bJ1PqcrZd4eQiOUNDf2CDzfOESvnr5qulyuGbvcohCJ0c+0SWw2T12Io/n
xuIgxPWbCaTbDa5rRWkD4L3r3gwigTLbtLGIjU3t/IYBRK5UYGrCqZoHXPlNqQ7OkIpg2q1h/Nba
uHG+3Tvgv2kLdieKJgAgZ0uNp/hzfmupDn4tx2gPTM5st/ZdyffjYnjsr4vwjNJujplXuu/gAOQR
FnhsHD6gp3esYt3/0IdXhGCCSj7PxgFHC9QSHrlZvoW3cvb8yRq42n7npYjRd2g3MqlTkaarxOsy
wcWjv3O42iT5n628GDc2ch6JD/iefyr4vdEZKOBIBpRsKWxgX2549qan5TN8p/D6cBInbvj8pfXc
v6UvKNRRuiqRV9FAChsMicFhhFglrCXd8WxU1+WoUOYmkhexGF4zgUgqdsjjqGwzmtr+6xqjgVZQ
GvqSwdGPtXKmmk1X3c69Hesg467INd1FXeDlkKcC7w4mbo3gFTCPTsEwLeScdPBzd4SPlyhCbJzG
ytidSFRRmrOqkCQ4qtJRGyXi5oR784dgFA1WTH16kwHW0uJ1MDJvW15ly8e7i/f9HhtckFouhmUw
nKuKRym42zJu1mAqyEOwIimdLcZNGKcxT8cnjauCgOVcILAq5S12KEPpbOBg3p4giVwoR5hVZD03
D9p4JE5kUzJjJrVlGx0NMUzNoL3tABc1ljpBr6nNZrjYA3O5PXvH17RWVgpdRL5KODEGz0xAsMWZ
aPZgkoojxF8b7vSaPxVV3Re2u1JGvVuSRy+16I7GYZc1rpgkCt9JNKqmSbyvdqQTz7cV3Opu8bM/
VfY64CWgTypuiqu8kPfXekqhfs87pkvr1XC9AqtyY3WTdX4EYvb8SW94+sSgRgmboyRFRlHYv6Tt
EupIoahMfFpt52F/tEhooEBKn1LHm6xIHk0Gv+X580dw97k2WI6v55Z7ksUnCpcZc4vOpy22aoe8
+/luhkl6j3bKVUeFZqMVFsAcsbvzd2uFXs0AmWKhSc46Kwz48GLhhGDt80BYbrNO5iXR9OkyB2Up
W6Pypt4ciQDx/vukrx/KL4kgmL7MN7zwWKouBNMqCn90njbz6U7mx1usaH6z7pKf6aE6YEQockIz
Zihv3IA0v+P+lud2PdM4+I3A/PU09a0dN41qM6aiAk2varMyYJsL7Ga6ao7SedHqriec6CoptgHC
UNzOm54eYPmE+OmDJs1HyaSNUWlaW1+H2EzUEE9pBnZYHiwycJ0EQaVS84NpUhmX0HGHnZucKsvz
uGgSd5irwvvdmy/0NrCp2HlLTvmbSmx4IqBmG8gZbYPG2NCasLSDNZRxWH1k/Oq1EjDyeUfoHJKl
3C/RcjAxtt6EfbB2EbAUs9nsEPS4WDNKoG2IyGzIXWHW3MbIEwpusMX25VnfMiabDF8lp2ucUXzl
vAhboPpMUCg7fj8kSu5oSKTCEfgWFis8vXsrHZKmqrfHjzjp8V6CXMKBvXoTy6VLsWCYtU7I3rFz
3Egsv6Wv1OslvzHQn3iZ1L8HEriXCZV6Iviw2JHHfi4RH2+mcRBYryz3A/iW7QGV5uHME7pyu+zf
nwqQrc6xa79OMNZTAD6gtb7aZw9MxAnDifArr6b0lOoLRcej+cPF00+wfmOwtzYxIzeMcU7JWCW1
eIBI8GJAifJGxRcXxY/SQnkl9+/etypiSOkC+84KksEnnRGog7V9fTAtK0yC4D+QM97mHlukx6jG
b3tVR/mATwKfTityy6Kvk4DrJcpqYQbvbI9StV7ETIvx0e0kKyeORSjs/ddg1wXPoFgENAialSfL
2223v7paSlaXIPOfZ5eVG33UjriPsSCN6LEcYrx9nQn4r41lJXEMQSPxOp09dH+yjCYrSYUvlcwe
aPkNS+6gtOqeA509zDtnj9TcMkFWeTS61kGOTHKXetJXu8wySGDeicwuE5EETBDFZKGXjBjPislw
D/eiJkgLcC6cos79z+cplSpujPP21J237JNLkx/QkYlb6r1Hwm6Xxq+pv1LjYit5yxijoyk3w2wY
sf+5rw5saJnEYmjB040i1QpoNKbFVGz6DVooNIyLVT10rA86QYdxWeQQTGNzH/afEs7VJk1pNGJu
CDl6gL/gSvgwOp62GntOhV6VxLxXW4NfOBo19AQEhlJSfXrKHi+0EjCXe0R1UH0fsc+ccG7qPmPj
GnP9aMcqPMVLUxdhk4pG799a2XEaXCzEwUUPZv/rshqcmIUtuxF5BaeIB5mGx1SLA2SXwotzfpnU
9PkiXKaqcu29lM/nTAnXoVGSKVhV+CFm6+pOdKphY/vACDIj/dynbwLjEROxcH/z6DmMKxEHO5SH
mz0YzQdDZy/1PTdaapeigfSaNP6RhXr+xrTNSohWeXtXGZSuAx4R78MSK5VjmhumVlN+5it7zQAn
P2tOJVdCWOQRuYzQt2efVmKDBVJlhRYb0y0zNe9oZZtLaRtirY66V/IO2xPA/VsYLtDdjbVX6h6v
f+jVVB+G+FE9eHqfVpHkV+4gBbqs1VFqmDE9/p3mx2CcfCxveRqi01Rg8l2qmnNxdFtljzytNX22
zAWNQ3nA6ixXdaxEzYXNmRbZM0QUt+JMFEKuMkcQqQ1stGDhu0E0lrGcxrccM1Mc1wRfAX9ept7Q
CafW+0z8Xz0kSZaqGh8i7yaWPTrBrcHspzHMVoJ6DFraGhAxYhCVMtePY0oBnFmvNCMm10sVKoE+
FU4fHFvmQfnZa7gvTSdUITpMkCeih51UFDLaQ1H/mQ8g0LcX5ei8btRKHW9BrF7TsCDAuNEAo5eL
63sOOIENLeKE1dl6iPFlKYFJETOLcMfRV3eRbIRZzH+MZRHYbbIE+csDmoBqEnwcp9eO1j6Zi85T
64JzPG3ixrld/E5+u9G1ITZULjipg5k0UzU1LyNeqP+XRG0omzXnjKHEPSvkWXp+mLOenx+YhMo6
EzUQSdKBPASxAord0wXbyqYj1EitEL3YUlgfS5/TXTjfeGjKuyxQ5XzPmu3MdO0+CswZDCFDl/yX
444cNTDAiFvIvQhq7xHZFLhWQuzyjw7QKsbi3j/ejw9Q5cMfnJfSDYHPbT5bitXdlnJxDnRrZcIp
xIJdq83AtUVk+GF4bgV7Y8riNwtoZym/bPhCbLJ5DAjDhHL+JVb5dHSLdPKRDoBVlveWzdG/yLQ3
MfGKgYZCHmpJcCxkakXFRials8kcO7QsTcnR6CTxdxoDS2wIeEwPrAqotv1oBcIAaQ/d2dZf6jL0
Ev3JnEjuVxqHp5Su9RDzRtckuLhTioj+NgTsywr1EVjfWso3pxq9DwDLbsF/yxv1z8Av4KcdogjB
JEzvKq6Jy8w0esASo+MxvcdRXlKmwvaYASLTDrnBe8K6bluANE+YCCkiS5C7D8sQzlPcTXTjLuO1
vM4ecia4yjcKGhm7y/YytvW3Y5XE1oUkVpfbWByVIQGQ3sS7NTQKqrGg2H/GzLtDGp2X24irHef1
mFne9xatMAb3vJ0HkZzNQ5bJeVm5vTq4bm89kExPFjeNfC03fZ6N8t4y3Al094+HJ6Tzz8hwOdFS
ptqavqoLtSYoVcziYBz6ScLWeEwah9ANsukO8r6B/361PvRZb80iiclW+aS7d5r2VfZTHhW27vEa
RL8SxgkmfShWhrNHgEuV2IiJ8nbfjZ0IvDtLkP/Lp8yo5Y4welhvBqYibxEIIEvT9gejTR4Pm9VO
ZpU2AetcImN0YZkq32iSal3GTjS0w1vMuuY0PHWGhtPy4Cwffpt/gChEoN9bfTJ0BXLGV/yY/We0
R8aflSsv8jK64Jv6CHfCbvzqrpkzW5iRrOdyB44T1xG6Ri/Kh/KwTAz12gYkmzPo+/un7TXTdDGD
mvXGtwYBXBXZ/5RQxolxVJmDSqpdO0ZEcECAUvqJT1KD6xRK0jxPP0vX6JY+BRwaWybANBbzeaWC
zbEe5Knh0PqHGAHy64D/ie00syLUF01lilc2UitnFBZZOQCXJab0Ji6lh5fniKuOYTPaYh5RKGkp
Hi/GBandSSEYe+JbIvuVG35D2pqWK8IL0e3LgIODlYf6YflwTUir7LhPJbJD2qISw584Ywb2zKny
oh0Uqxz2ITR9sBWb++eqBUdR/CNfSC8y0vPbXNil1D+8D4iaMAotNkQ9T7ufkhQ7yZA7Md4SeYn5
k+wn1gDcZIRr6cFCCIX9BR1CHGqAk+0jz/J+9o7padtpykJXr2OSZ/TEaBk4hTHS6AEnbdR2KZhR
vkciOE0nb1Du2ewAmiIcQYava5rBbYnavGYNDeg1l1kR/uNFpfD1e8p80i2TdBJTKxIm39Mvcez7
ZSbX6SylsnkfqtqN/QnvsgApWQEOD8JF+7ZXYHP819+k3iN6G3/HrCeXroZcLXhUi2sDVIhDXclA
5vth6tBB49N9lqadc5kMa2JPeOmCFLQw6fX+xYNRw9D6fldu2FPnotOugWNAigKLJcF2xrHDefkJ
IcopvA788yUUWU/NM5Twx7bLerYVaTgnIcFJMV/uIUYIhKPzJIHUzXAUW5+nZiRZ71phPaIxsAiQ
4E9Pq6J3vAvxsdW2XrAPyealn9rIMra8sL+k5joGgl3BUuMKmbRcgJiC/YOQ/XhtUDr2Ks/Fdxab
qusjYtcAgGEBHf//BIm0Eq0qCwmIhQAAEx6qo+AngS/hkDjHy8NoLK8sJXAoIaAIlLJPhxyhzhLw
gveJ2Ot2Xy+nqREDZ6UwEkpByN1QJYxy1WSYVybm8IOy+ndliQZdyuM+l9nx8U6GV0PrSsSXLvjP
tgf7mdLd07bPn6WDDyvs4NjERZ/JRlEfMakbSowOILfp+rM//6964CEG9DsMlL86l4u8sBdiQR94
D7laU9lXkuHHuD/4h7PNXJGgQhexV0mkZ47MKmOE81RM0Z0Bs49TVGXUyeAXyRryoiCMnD4OX3SK
jwXAroG1rGi5QJ2o/5Ny+Qo7L2IFcdSqmTysoI6RkdWNv7RPXnJXDxX494b0DJRPTcfGgnBmAb12
56ybcgFMlhBPi7nswhucgkaNiifmqiGmyTzVPcHpZUkaBeq3TuiBe0Cfv8B5dhgKcg6TT5E+VR6u
HiJ7qdGskaElk85VoAb17JVsVUbLEy2kdGrzSgtSCdPyWry3wN3eDOb9yb8OqDZSIm9zEvpF6ffM
A3CVKhVDVhVQfOpCcRf8sghCyk7MhRC8eBW5gDaIfXBlbrWqcVFbstOLl6XGs7u2wIVPbHdHjPfQ
u858ds4s60/NH5+7NLONZWHwsEbXJ6zqJguP0PZ9O1uYGURYgNeED99p0J6SBG+ZEfYjxIohBOxI
552C3A2N7qWrp7WG+8z31N0HtPaMH0IYCZl1RMfp9Bu0AR9N2zfNwIff+u9XDhLNCn47VFtvcDcF
ZfHV8pj7BZFz32p+ofi4H2FD28P2dvHadqASsO6LGGvopbx810Hobw0kXo6hxM2ZkM9AivJ0g9n+
VXge0LraQwjYC2TRkqqrtq9UNS6x883dqzKftV8kZ3PQvln7rwugM2hMD6EaUokjXCr2iQrgKtJp
S/xhETG/JTmiLFqZb3m4vqEfQJwUo5G1ClL9qz+VgByKgJEAUFVsFU8Kx+/36qsWgH6ZYZ702Mpx
HTgmDB5wW84aLwtHlcUYKaacKDQorytDzllHmnwMZQ8AWRkqX5N52HmgWxYrwIyp6m3JjRvdopWs
VnVkEKWbzlKLruc2TgGK1NY19zC2Ynv5XPaeW6xz31KwQ2sKfhP57Ltk3sl0WYqnzGI640uvYU+Q
1hb9F7Ot+/wTSl+fGquTfiJ9g2votSqKCVHWS7Cqzx3L5ofl0y4yUKkq/e501w4unJmHcMG28oJH
4ICS9uuMW28HQP1nEIW1c1bX3rRa3VWxi4+9vzWgwfZ/lYFv7BkG7OF+hntGPTEztd8Rz8PSnPTz
VITXAazRLAmPxP+Bif6R+sIk+Jia996n0Vi0VaMx21ng938fKsULzJ3S8Yf48QuL9cnJ1KeA0Wlr
k+Xqj6IzBwKXPyNeHz8DkQsXwnDhAq6xgLl1lwRypb5OV66AxUXyC1kjPP3tGykz95y42NWSawjZ
mU++CdE5LIe3mXfHGFkJPkZZeSEKNy0VH18ZlL8dJjuXYnHRuBEsqsEe/g4IR7EQRPMDgzLfzp41
z9oPU0O2FoBy4Fz91dn2YejcT+/SPuPJxQtxdTsa6RAnUH4G0QXUDPoBxOF/cO2QRJ3B0BuArs0U
5Vcyc3y4lMTAPJrNdrv7JgAsFmpBaTbfAIDq5xqrM7zNrvdNziytNaKK9O8/4D3WSUqO+7cQ9g1w
VauJyQ6l7QTvMDY3zK0AxEd75J1gHIqih1iGF7aNJkIpYQN7GM20Osb3ggeLxiUhYruZLE6UXwwt
ciZtdAiG1wnJlpOkwDTmjaqWfpsoBhl6aM0iqUuR21rTAtte2P2GCrAZPtma0hQmCciuO9K1k6to
BlpzMV7wwY9NONEpqhShueN2z224u6QNqb7Q1G7KmSwarAz3MWNiZ498n/ySyhaixLehyPYSRXKT
/bzLXORnsJfqgXfx9HwbipNUZz0uUSkR9vGMRRsGZvL7zvEEAZ640sS7QYqXRbpvpf/7KXyRFjt5
dPGswdtbVXS0ofy+iyYPb+98CO7tz9GY9Tuf0PZJYEtUiMe6vknT27uXWAP+uaB9S/yauST39Gh6
QvHdZQQosYBSy9d2b7cr4XtQtQM0dQYlAEN6C++xyHceUllMMYxTr8/lpMpFwoNNnbIVw5S2kuXU
rJEA5X8SkGUZlToR203nyAIn2WP2YfBdjGtM7l3O4o4lOnZBtslhlvqmKcm2XY0i7PuXLYOW/cyV
hsCPW5hI9znN/FinR0bURgJSsHp3bbqX5bTO4fVNC8ZqtNEfjR8SqylU7KuTVPYXuz0AWE16AZBo
/OLSVF49GlaV2nsoKDc3RPBfRUZ1VJv2HWUi1776Psv+6TAVcnyQoqRKkjn/Ly81hTvstfRg+w0W
2q1E1wV4vPWyARXbhQ4SlLXzsJ6jss3z/cx4cAX1SSxvVNY3NNqQB3wDVPVreWfPljjrnH/AY+dz
URyCeI1RsWw31/T6erY98HO3o3TYjmTSjtuXytZSyO/5Zlu0zD+Yg2guQQxIYeo3D53cwmEL0vTD
NEL7S2sxz/c2urnQUst3ZnH1Q7l3ffagHoeZADSxTKvdjquXGAHMipsIQaZSVEyZnv5OY8Mpwujo
Jh9AHAYqEKbHlBJDH2NU4RlqGo1sx0LyNBtdRbyblC00QRQmBNiJ+HLOTIuS/TXWyVDiiWqtj9w8
Agd3UKyCsOfYrGBJam0T22b4l0RgS499tWWwAz3JWeMJ/HjvKLTnmqSs6eCP5akVBWUXXl39zRFe
orgMdkYCMRS1vqZtLpSyCckdEHqXqXHwKzEveMXDP9L/JRBIte0lZjpB+ab7waNv8WzOKcF/xx/S
ta+hOc9EQ5kPZNp4+AupQEfHm057HBrIZ19xFRL0Sw3BtPM7OY1b68eQEelV55RK6RaP7FWdWgpv
7b4wPIsuJJTj1/bJugaEGb/LxvTblEZihkIfsuLULZlH6z9EZh70G7Q8IlHP2P4gS21GMWzIktZD
dU5G+62qiNfqvxp+yLcxH1Bn1FNDK33/sxAaQmTart59TsW7Ngd9G0XzF5542W0i2YPTmI0jCqrt
+JF2/L3g5+prLDl5fBq7/o1jRyvDi4ZMG8OlJSPQLRBlwEP3VpcP+We2P6bD9snI9Q8JH2AGTuTh
4E+45bB5WjibZyNj8yFkdwsjZrKWvYGfl8UCBlN+PZNlgl800XZfIZXZ+m3m1hp3Ag8mvytZWfWP
CfuKd22LDGeLjR/n6VWzFsKdNvWM/ScHA9RcgTZx/WQ/XwwYjRSTmNyvlDtYnVnxY91Y8psfCQlJ
pZS1ws2No1jXu2jKzyAB7R3FeIT7HYsCuhWGBPRuWmd7jrHnd59HpmP2quiuyDMybiFNnQFkFs8J
ZV1ArQPUmh3k+E/4II9Whv9561dMCYqA4OMQQVGFBmYIa0DI+EV7iSnR+SuamwJ3ECU3GKeUMxUv
uS7wXFdPIVaag3wdFzpUvBGtKWEaRKPfAqMk++xHShyH5JZnN95YV9VDBprKi895KcKpPtNLmUBk
jlDGHGy95gAYIsDfIHlZ/OK+ztti9iqWPyIauqSSVmXYsJaDOB1sGOdJ7zGN2LrftSWGguNoZYgs
NfHMLBOD9FgJDGJ3OKU0jws73V+SRlpA/Fju2DZslOW2vhmjXoyUHCfAx8UutXZ5HnXDPx+r0GVc
nFTOtulRXVTAFJaTvicbNCkxlZvewhwhbgqeVPd5cKgqG08Uzc1jVkQ2hOwA2BSk0DVXCbP/aHJj
H6amDLrgwyw53cR9jx4/PnNqjHDECE+zc7HpZQr1TSwpWRDDSP6WScSN2EHFEbEUNzE1kbMuBqF6
g72c+rTM8Mh6aJbdgk9D+k3cKsuSakTvSl+Qd8rZdr2rKW8seN2yjfrV7xbaQ071kajmq+4iiVjN
cDFHtckx+tK6rkISS6tzAJkEDPasnQwjthF+hDr3QfT+Po78iAV3MmjDKjQ2W1nstTdbSV1TMqv/
2YeoXvYKcpeXqy3LHSFDDlKrs7RTzSRUS2ashG0hOUayHZqtS/tiH7BxMgwT4G8deYW+qPiQaIkv
j7HHNlxgJN0JO0JgMhy2pzDlPnZ7sMd+4c9N6MlP2CO1DKUXdKP4cwQiC/PGESJ7KlVKoYcuU7if
X8TtsiAGuw7QiItNKqSUdRbCqC6HgtfCfGJGMVUkcWuOWdurO4uuXKD6sni092nfnldbWS/Ri1Ye
+s1yBcAJkCo0TjdmtR31vdPEdA1D27H59Cf+sDyUDzwpUA63L42dgtqfJzfUolSN/MZHYI3FT8uG
/FgT+QfGRKe0B7J60zORRkxWWkDul2fFATV0ccUYKRXH3XsHzaUV/SIoknFTdNQpiK/NOiNa7imC
o4l+l/VLp8dn2BYr+vdKIKMoF6A+WQBshNoM/byo8vfeheMkERShhCbDMgPspL3XmkTecQE5MsV0
+ACGDteUH2mZwjMoO+ZrhMsHk9Y1ShYrEc1oQ81sWTeXhkWz/Zr0T1rucVx1BLrjmpJRGyQIC01H
/GG+tSV1f3AeJMkSV+nkYG83eR1TZAsVP6IopgsoQShFN1cJK54EIEk4tuQsR8WXisjPm3QrvydS
6VxAxKsbg+8mofx8tRsxA+grV6rpaTqcj5s6xqVBRvAjf4XADjjureENse5MEPnWjZVJ2ycinIVY
9rWp74n2XVm9NsOXpmUx5/u8PznDCx/EWyX5jKC3S6u6KymbKWWJu7MpBVhORMrclekb9GChgpTd
lnV465KGeAIaqNdDz68tOkM6jzOZHqI2c42IDcQDvsqQDUq3Z4Ay9Z2Uej3vo2xef6my6nB0BYOG
uwKHjChHOcwsf06r7ZRWuiLYKc3/edLIqkqj5ZNpkEFrpt98osHfP8o2z7jrkS2LlGpgXolIrj0J
DSzTEPmy0TTAHQflzDtPY83g4lQHnYHhpOYyDKeGpRYcurYH9sFOWmhD84C1SjJDL0kzPWpOBjOZ
IKz7cDlllRNmCalY78rCmsJvAWQJYfzi4wV93EFdlbSd5npdLVbU9T0uXDaBnK0dSndWairynINY
YnlB/obuS0JxdSb0rz5Ucqb2ib60jQmCUfS2PyWPG4owleKlXKcT7jdudziTCrolkIFthm3/bHmZ
tgNfr8a3k+Vyx4K0uAYSex5Kb1cRByqVzQD4jiXVCZ3z3zca+Hj19WwYnn76dNufVOCb4bye+L5t
HOjK6pdob3K6vFPJGzjhWH9bQROgqh5oFykVKADUQl8q2lGolEh5uJ2hZ/GQM546oytegEiXtNH4
HIHYtDIKX2UjrCPfmzmOHmAR9uX+wa5iMQnWXGUSVpfjJIG4CmLZicKQXpHcHdKkPNuxZ4AceP61
R1P/7K7NRzIz6W69HPkQSB5ElIkXLm3Y2LRCIwTYtbnfBr0V29ggpryqFvUMVcuff88p1RKiuKvX
dNRW9CmNpO7/E8+VdQ44lZ/iYypICyXSzzSqxTseML5z9Xtncv7rL0d2XlFErwR/ihZ0L/9sxVah
DV0eBp1hAtT72qZ0qFd6g2Yqfri0aRnK6MfSIUfjFgALpyA8oNu69GbHQ8RA1x/GhrJ+ELmm2Ltl
RitG7OrqRY5hrnBQeXXV2a897tVF6s1gSREB8NVnL8pnVUoVJ8ab1vnedrDrUvSPDbC+6T4oiwga
BWn3CWTeeC3hnUScs3uOKTZcWnJpGU+eCQQP1tHMW11zNKlqkws7Y/V4aWuy4tYnGiWl0y6a0vv2
N+1U1brn1TJ5fLpqSmXj9ZmpdDvdm3JUccpZXILAd/s3tMiNdVKQCRgbp0NVzfbiQapUDT2AlaQp
3ltv0kBt7zKsuJdLmor0pxJJl7YdBZcDBLA9BSbzAlTWDvwB5bpgwLjWl+IQ6U2BHjKDWg4543AP
GQxVg3ouRD4CBwXKWg8RcmFHTVwfvj9J2gwKRBigA0e2R54tyY3w1+hgAZxvQiUeb6RLbF83/RrK
iTGZey1wS6csRXlNw+hvEtZDIZO9OLj/l8rgtidwytzw7U55e6wrdQCT8labWRyOPFqewDK6/Upg
n2ZGvNs5nxibDqmFqQeCOSK/LsABD5TDLaBKPDMHBIvSL9QYUCYJYeSYuLQCwUFaQkKqHt+PM0HF
2A7AHvzoFvd3hMZSa1C66fpQNUhE8KTaAookVTUzCz+x0CUBIYHTQE+dimrpt411DUZPLWNHLRCF
xEpKrb1Htj4CQSTg6jL7DyLzrDR8HWBGGzB1ezLjM29OnN0LDLoh/mx1F7uK98ha7JocItLcULov
sPjJyBvLX+bbSDRtM7SUtvS9jQ8cY7IhqQ069/Xp6U9mcqnK9lD156Jp2eX2g3rcrAH9XL4O4F8J
8e2NQLuNiyR78CbsQ32k0SAtYrLc5ZG4oZOPQb51QZNfgrWbIY4s8j82aH9QYI+vZY3OlZK3Uolj
gbdNcpVDeNi1Jc7gZCteBHUVh4gGLgb+Jr3HWYfJllmNCtDnbO74cZHGwtV4e8Lqjjl2ddvx4ZF9
Es7MoxjTbjIqyF0KMMOzy7riFSBypxb60yzY7G6SWgoJA/gCnc7VCyz9nAcPX166g9TMVulp1G4a
bLzxEqceorm3AiKgy1nX7SzW7nroISKHH5FbLxIUUqTMZjpf/r/oqd7SWeHkQbY+rhwD96cMzNb5
3D2xfuRd1477APLqt1lEADQiyETSlbniZZBIyuX7rnB6LVBvCD0bsL3oDlHzsGUuqIR8V4aMPzSz
8jE5MoHrHCs4cBS4xuQZn+6DK1vdwf/OHZ93d/uM/fvQzR2KKAJxkmK4n7QzjGrLyEqAqdjBBBVI
0MJ809tNZsmUB2jwjEiKKr4DeIjR7VJGHMY9YBl1IxtYSRT3PZy384Bv+ct2CxHBNNv/TahYhVFG
LOxG91N62F4X8iBSYKQ/sgKXF7pfvTXLFhRzEM44UAQgLQYkqeYwsaHwq1qLZK1/JEHMTX3ALgqb
QiX9MN0vYLZg0NhQBxpFBJ+Tr35vGeHZAI+pIV1VN/5iXXy93GvwFI46wc6sIGjqDF6FU5JaM7kv
iR0qcM1Rm0wnY+n8n0V4d6cyfxqcbrOvBZzE9+x55r3IHqZ0vqTPBuJWqfPJWmRWl25tmOvSd0gE
2xQdYsWNEbf2pm5SGpWJZ3HCOB/7FXSxDK3aUHRzF9tdpdCbUcGMbMVlw3wOeQYKJeIAtvsu5hpi
3UazLnSC+02/skMy2ePrvFgjtP61dxJuKug1xQgrtSth7Lnz/1SvaeNkVMO1/oMigrikJ9JauBYx
Pd7cU5AnFr0Xkf8QOaG8pp6e3KHvNuBjek9/q99tuCW4HH9bJC1AzMhRpWr+g5APiXiGFr1UJvqv
IF3qZdAgiZE5QpEx5Tj4AZD+ulypxdrWu5mkD0UQrz+AEBIRdsbA0E52I+AIrbm/CXHNj4AV/Qnj
y+pP7wKO3XN+YhKRGmJ27VN/YXtjbabcWbUr6eg/ZFWgoxKToXX7eLq4IvKVe5K26iXZ9W3oDkw3
+l4RjeFaWY2P0rQANhTV7ykUkoWrYGrA9X5h/Kz9ipYv2X0U7pgs61qsEjvjrq679ZCU+ai6XsYf
oJfbKgOofXkqLV7NPHTLxR21cp9QtpqAoHiaqsrtBYM/LDusu46R43lXjyYhijYFGa+gxCmCoCs4
Fg77EEgkYMtafivc7xwtQ1ypqN5XYCSjyOmrkq93tyBrfJfmtQQ51rEDp0QUGWloQB88sOho8Viq
xDoi0jfp5hL4o1FgApKt7k5h6VDhlP9hwluluwdzrlnjUnKcq2XqdGmn654TfYPgN2VNJmGUg/YZ
7aga2hx6N/K5mjBt55dCni396rSR4ZSX9MW0whY5t6F8cc7hy29z0U3qQ7qJNAbNu3BkB8VKJ5DJ
hjmCjFSQjjz5z46foDirKE8OSYMek8EvV5/1fIv/FKPr0zlgww/SuNTk6h7qYUeb00utEvB9CwMi
bNIKLHwqJHMFh1Hex9x2blsG/n2LsVqA/RBHCd5Rdnbe4b55QK1pDvS7oJXk9+ydg8+HMXS2HPKy
ooYdKWCSqSM1dm2YBy4uWgohxdC5oR7A4x4XzVWdBOT186TAMbT0JhqM7esg3RKKTZhTqgEfOk58
oxhQYX4sEGqJDTvtJQL693T3GzGWOeNEWZupI3VNKR7NEUf5+L6S/fJ2dg6toQYxShe/m0LoGhq/
0Lk4wQpXYw16kBq2FA/b+1CrNFEcarEJorwStoeBOt+qWdrXpqsgz2Dka3r0YDakywUHlhP3f8L5
kZr0+S/dqLN9mWvTsFV3CqlkoWV6lpjq8FWkP626uLdjsK+lxqNmtAPSdQEA45R+nGKo2kuvrURf
Ywp5NDnIEv/Qyt764cpHWe2MlxQeFHuftOUucdxTz1bY/5zIASCGv4HpYEMTgPIMKeXxvZYjC3hf
m5UrDY1IEC5GibSy98cijdvcLb8sQXBCZxG3wbc6mUaubrdvrY+8r8DUBHikcdwEQUJRdXE+EvhQ
eO2ePrMheszdIcWXyYq/eVPcBJwk6Y1LA5cWDlvergl0hman3x2n8Qqgi0JzSOr/kP0/RZOu6jZF
UbXGAiQnZtSDR1t3/hXpItXsgSATwRekVYIC8+9wreppQkFs8EwKycSiJBJ7PEyzW97IQcv3Otx5
bzOuntfjxrMap3VVR1YtJoYTLEN0R96YDWoxayX//glQUD2wP4oWCuGiERqFAYz/ZJqLkOaiglG7
ktJG+dADwt1z5biZI85W86OJEkMte3PGsAfcx/PcotnZE9yekoz0ZXbw8r98Ebq2GSgJ+zWnIsdp
sgrpfh0hDvKM8HQATCH0aYK/THtXalnXIcwEN90edcf56uRIH5Aexglwu+4jdZjYchCpRHrTD805
zH7bKmDCV5gXQ/gZ8GscXvHHafXaHS+9ULVmU91cezL4PPjsNRFSxphxdaSDjszuocoqCKupggel
y/Kh67NOZuu4k+DZ6sZvqcXU8TL0938Bt6WhtIaZPTXIj9AJMhxN5W3yTcofYOfQldA2mYCiVD6m
epqImo5EpVJDwvkrdG6smA3fyenL93DZZNegxZZjCYmFy63D/xUtNXHnnt6LUw4lDdaKSTedTyBF
aQpW5Ceek1bmeIyXIa+ykXsU+6MWvul8cEAUaz8q6EmrXD8vhWl0Mvuns0IOfgEu6QZWcVeOaqlY
o9sm1eTTCCFW2G+9/Oa9HgtIxMUJHSKZjA6C+6EUdU1mo+KOXP/dA5hXFqHvgtx9sjyUIktWZA4F
kZCXsY5yTdL52WX0CncWWVa1SLHAnzDbyv2Z12llSteZQvvqbrxUGoU2kwWkkMtHKU2qSkFFfhGg
4+0gmWQTAGUNi4F/KGTgUwigH4zmzUvFZd9wFFpv7SPp3DOhrQpz+fJHwxTMnVJ5fFz6FE9eGzj0
YWVdO7ONtg43Z2oPJRAkt3n18bx2LM+wC/hXdvvr0pGQmGKP8TIN8F5VZJRWqSlrC3QyGCeA0DdS
lF0BD5HGoMcllj7IkspfBpv07tINXOGqIxhct0Aa2nPun3JmRUHQpcODPmdkaWK4JAWvU9oAUMcK
XYYKw0KDSZea9rGtwBmNPHCGVo50L4EjtYbtwWodQRaJ5uY4wy5kKXrNOx26geOlQRI8Je2rc6hq
+3vo5p6c2CAj6qdUSMw+gMJ0uPEEIZRksZTDkfTes0SnMmw4VOPZtiV8Anct2ryQ5hGyS7pEJPcY
2oHB1gCmDlrrkFdMCDmswEajt2pXxXTO02itg9IKZgD3RRmcCxU3Lh+oCxJgc6ZfqsYixbxs6spf
HPneRFh6Q8LiXalZ5403BzMHiAppTeZkmD8qkxQ0WuL3U3GVQbS295Yyrht3fN508jNZYa+A6/b+
nxEiLpSsR6/vUSvxPo2rBgjlYsuuWbfdiKNQGU+Q+BriNU0eQEISMsYo+G8gy2Kur4o6iSH+8EFK
tfnafq08PEulvmjZZfvc7fuqflTVWeMMqh4Ru3OiVbVmhtE+VkIB/tW9wpboldl/7XrqUvDkqjUm
Y7tdBAjEO30/J5PPtjrq4ElNKq+Z9xR1duY35sHcyOkkKsJxFIyS8kuoIMte3IvaNH7btX1dIex1
46m5olz1mIV4BQm3Q4HLa1LRncDzVHT0iwWxVdF0zeZBJG9YMEQ5YSNTvXAjTDwS59JHLGNjxleg
gn5dz9yyra7Gt/ljGzKTa/pjO9/KoIm1C0uBor4WNi3GYmZlzf6aH3NpXILfXjvP6ipRTrw/ZLLp
ZPZHn8pub7mN/ljEVnqCiS+psKQTCWTXUz2Y+b20ofrTubm1+/xYBLdoK/PrnlUbihPvpYYTP1E5
bJPQvy9bkhvVrayrlkK2nzD5IuGTxGwBgpeA9V21rYvlUMJYdnho/yRtdNpXsGBvAqJneP0gUvEd
Obw14+WpkdZh94OViLWB5p3h5BwdkZ0/uRvKQ8srlGrLgtdS2GrCv4lmvM49dNA84nDOmr4fO2ct
ostdi2fntARYiP8hsaZK+dAS4sAwF0Av3PdK2POgkbBFo9rEKVmBb2Vv9Q0CT2Azyp2OmwjiGlbE
/AVr61WpBK7cvtmLifh+EzB6u3jGIIur8l7JXCUNU47X1WYfJHV2QS2DNDuqCxQ8h3nQIGYnVk6I
O2e735iaing50V+w+eJRGZhPA/ap+PJ/erJrphgKptakvnMVvmHzUOsxtL4ne60o5GRBdLVJv3Vi
OwXx1IoI0WG3/YXFQGW2879zABExPPyqnhLHgfERFb3g23m5djUpv/hJZYCPM719EVq2WFxSqrqH
TAeqcMnlUb+JHKM01ZocnmtzBA9CQ7R6KILpUl/CUyPwuAxau4ZhRccN/FRACYUFddRnkg9LXmoz
+awUEirF6w05Aev/a2LjfI9yIlVDogQG/N591SsT8zXiPyGAHjE2eYu8ZNEpk8Xw/fAvuDy1oH5v
BOujE4/fPannlI6oEt2tkQ1F9Nh0CpsKs45Zi6mpdDUNwIyYMJoPBWnFpmN4YGyFeCtm4pul3UgA
z8HajczpFTQtfchyBh5cojk9mmmzPDqzuLD+vVQe7J60v+6nAhIC2G95ILP/ulzzaAm9j3b0jT+k
Bz8o9v1XnxaxkUHPHvl3Cz55HPQE6VCa6d9ansRM0QnOJShT7XCfi/nvwGiIqKmAlxeUZ3uGo69g
rSh74v/TO8q9g/XfVSKcRJXE8EU+0HbnTz3Ifh2W++ITRJYjcW+gVORae6suzc0RfvaLiD1HdOGV
0OCf68PbblcgRPbwYcPFLujongy3jLvm3a7OPkbX2ob315eVsuWT9Yq2atIpAXkHWzEbzNjRvvbf
AZxqga5ccQRSnW7rjYTVkBiI5vnbvpohePnuudFxI5fYsjTA8E1LzmuZIR0Lukx5A3uI3awxPuo1
uJYTZJ5riSbJTXjtKJ1TKsNxP9lWYgeMvT0qYxGqHxyMGu4VneszwJ5LpluGs4zdPw1YNmIOhLwR
tUFKxCOfjRYQXByszsS87Gy7a3Ug7J9pNpNXg5v0quas3eV9esEL8Rcvy4R+m2Db36rzKWUNr8YY
Co6HSYv14FlT9xAbc3yI9NFXUO3hQrZbNOpLVvAbbjajF4Mfk1jBRkcCHX8SgEqY14roMf3H9GWU
XPciWvYLgBdEYL8rDYgci0aooePMFFR94IixB/W7V7jhqm2RKzNwBTX7Un0GFpRbTIPRz3xxIciF
HQWZT3Nl2s7S9bC3kXec/BS1WzgSmytSnMN8WfdC4dkl7CsoO2SyuiZou/xMqyur0T5qEjLlxcxI
eAg7ZiJc1tK/cULb8s5LmVIcSIqjuCIE4iArocAMv7HR/IwqE4kRJKRFREqbi60WlZKMGIC5f0Pf
CplpILjku4SbbYY/+YWKQgS/MDeTVRAPuCqL9zLjmXlo/5GqroDEN6cikHVWLyG7lpx57+PWP2ei
/tnHPpWLj///RSORsoRipWXL3e8IdOxZeu3jjAyKMJsEYMf1tAEOpuOf5pB52lSwgxr5IR8IRWu4
+3G+3qCgMUGerSz2YbpZUFDgO695SmXuUmz+q1u4IISd7gDpxgIiW45gtPxRzpCMgTuGuIXsV7Vo
+1k4BWx8AAJQNAVv3fvr1pdYjOZb5ahD/Russze1D0HES6RtIXmLe1LRKqXhAwbpZrUmQwRhsWIn
muMFv14oTJ/ysLpxwWiIl9CUHnPPAa92CTjUaPkFY1mste7KKW35kNBkd8HCiQT+bcclhEZPWbfR
IDz6AGo8TJslqfKQzDwmYYKYRohmvE9eCXgAFcc0h84y7InldSYEBSejkknJ7Y7Ob5DLSmEjZK0z
iVp8n/RK1Ygsoam1HLNiwqFDA+HD7V99kq5p0gMRVJqInA3RIvQFS+yjsZ/msdY5NzdZSJVJe8Ft
ALLWdmd2XtByNQ9vzmuYGHu3H0ITRhhIxhO0NUVg99WenxK4wmgHAmevJzPBgEUS8kQeQ8U+G5IT
6Nt8l/C1M+InF6CPevo10zaPl7SEQYE/M8Jnb+lmSx5iIe1VU1soIFYemXTCn5rg8zZJwvTgK8U3
Pymy8B20m4i7g0EqbeOp8P1OIXzRsEuQAgnCE7j4XNyrNRUIKDza1rMnFhI/8U35zacEnY8VgWKi
1yn+mzNG9bOzcr3jzql762gwhbv+VoF530elpXnyg2N5ME3/A2JX/3fAP2IhnUHUJJVFv+MkF0+6
o9JcpZhGrdF8P8O5y+dWktPXjuP7vY63b1ixSfvBhwXJ7kYwFsErwZi0Jje8i5qmFgC8PdYluwDA
TwouoGIN2cNTQRxQItH1vLBi6o3mYTI9UeL2dcF59pRhlXATGpcPp/5ykA9hAnt9bb14wPfBxgCw
B76Y8OPilbM97yKUhASJMnM4uK8TEpJnqwx9VGyh5Jk0/qKJvcOqOPquxBenmrRTEAUJOVXpEKlM
+ia6xUZwy9CWtu3+huXu0gHj34El4yY5tuM62EF7iilIyJ6A36IEgzz5QKYrHKdRPDWqbQEn0fov
OVs9vKaidCLeIpqMP3D6Xpk90J25y0kzXn7ePr6dX/7il2b7rNAudPwfeDO0BI4UXcq3OtSWXg4F
pQIRWemCeqq+QGdJBwePqlp46uVVcvjwpWTQw69IHOH98ZMCJb3eWeUzOuSZiAlgxNzO75wknau5
YWSyzy3FdCSoV/0H8SGd22sykStKjRK+oFAnTnKhULxupkJ52mMks/u0d9KkZsMMUiVAdSOVkHM5
buyRDUiYfnouhGiMcknAouzSlseBZdAfvGtyDejddk/yrrGTfoAmxaYD1AgVQQN8R0YrIAirAV8j
A6p+sukuR76ku6W2JgS1s+Ki62VtzsFWCduDByXDiP30zybM6eWtVZAJkOoM1DvYJMyMB/Sma/TU
EQXosaf6A7YQwV6/baFnAS4Dux88d96PzOsD7P1w7RXrEYqql+hz5GMVMrqCISf585FJHFqIwVtp
/XOHdQAxJd4Sz5AQfJmcHtYWivcbaUsZF708tWRT2GXBJlrKyYZRQTAp2g20bpYzncwzVvGxEXw2
AohFsyvLgfpLF+Ufokfl2uP7ei0rXUZdZbYSPnrOcfAU7dnzfdcXQ6Jid0I5H/eeOZvlR8mgA279
xvKleye2gAkpOZvAYqBRsngxL4Yyn5zFbtcpXH6GQaMZobSn+GpbJ3BoTJiIvZvmlMHdq0HkoC8r
5PSNq3WJmhglbtuPuS/kCqL2RntOf1noQLM4asMfXdvVKEDULlVvzhEQBYbvWUwlmrDUHHBx4Vm4
zlvyLomjLr6gYay6PS8Tgk2gPiHwNF823Lgl29SnyMHU5ZuKoAKmxXnBKZseMJrlBsCmhnbhSZPN
tF2pZdbNuZ+UJEHB+vhbqpj30zxeiXsJOTxfl0nGSNSlJLm46pKJCNg25ITOxBVTNflhut2CgBhR
B3EUMDpK4OurJhjiYX0/RrGeWaRJmXij96qizKvKee9wFezrOQ0sKEwKl3q7sUmCLHjGN1J0wh8+
XXViyHpLuW5HecnoweTm6kzfEg/l06Hor7wcneS4kSMm4gCXZwLXRCyTolMh0Sr0fgEMaU+Q19SF
u6lGf/69jeLHw/8PEDvI0x7GudYAB2tbJVyXY073DOgsQVfx1goVk60hCWd0ejIsGwvnAkHuJDhr
bpF5DOP2azRw3kMiK53wXxZ9Wbe2zXS0qfcxb+zUKDZ/7ETlj3mN1+OPSjXKHXJ5b/sD/ve05XIA
vnCWSMY3mO5y3/3F4sR+SWasfu3wAf4JMHqICHmKbxBU6ehymrk2T/oKw2Pnm+1waE/bW8UgnWYh
6csAvBvmewL+IjD38hxKXQIFeTSjs9393xVC3JKVOZqUzYWMVzbHtVBehdncUGdbBiUtwAs3Kx0R
16LpALCe66DC7hY5O0PjEMYJ6DviGw4rjheGhnf8RqEnL9x01Hc4sB2azBbmjMihVNJhrPivS3Oh
6WOaNr2zaU5Tt+EYc68as1Px0fGLP5Ik9rEUxcxpYSpCHX4gEewrz1fZ4miHi4HswZkc425QJze7
jpbKoi1nmN4vgU6ThzT6sJcCEGCz2mbjHNFF2fOqSJfjM3wCJO3pchXN9ymAHJ2Zqxmw4cijbKH7
EyeKaegIx3k5cCwMlrLR/aB6nxRXhvfnlvGVaa4OcjZxM3sFas1n1WABP45OLim3mAu0W64sT1B7
dQg+RkIYAaQaiQK190dVseESs3WTOoiqRhWaG3G5kjFXchhRuOTUWJCrJ8YdXHhDZerhwLvMiNil
OcWS1kc3xYj2cyk15wdhZ/UTsnLyTOcEuxz69xcvmn7dMFkEoQ7m0Fj2oev/97BVqiUow27wHPBb
uQg8Vck8sx8li1GTqAWp8uTlr3CIUBmaGBxYEKNRSb2Su7CM14Bd09b8b/cERppbFMALhpFKZRCI
PcV4siYXWy8V57y0pamZYM66N2un+yHI1jJ+rkOKeR/mnpw8NwNApofn0jvt8Hg8IJlnONT0nnNN
pP5V6aHbzdvJ4bB1iKcOI9T+LzCMPIkAx2AeD2iKx1NgM6DIuC20uHSY/Z6cPaa7kzJx3MwOAixg
QN6WvaoGtxOJp8hgBiIwhDDkCYUTTHu2win4wuM4FC0LJ7yorPbN3xLd3DpC2NiP7u1HcNPu4ewr
aOLBXSvyViTtEYTEbD5DaXHawstS4vvhD/gmnNVWwFDmA9otqjBf6ss/uM+taWjCE6Q4fLm+4kqz
QNFS79EN8JTSlpUvFWHqaW8n+qp8nN7tGX7XTzyRdRbMHNDWF/t8WiOifH9y17eqA2USIj1MLv0S
WUnvgnQMtP+bN0rJNtsWPXZv2rXAsLAM1rEPWUbPS++Izy358pK/iDYlU5Zval2cQagD5+BPA3QL
uEpNfQzmD+TOGU1I1+TTiM4ko6py7d/V1QLrhAZ3Pv+t0dOFs643I762bSNtH5sMWNRkFCayYKuq
jTFRtMAc/pIN2Q1vtDXllr8OCW+mJUwtnRoySSg4XngcSMVWojiYK3cLuaPMyZlLIqPhsRgiUoQL
lU05R2uwhM1mkximanlh/pCbHfQq439DJiRryrSil6wEfds9QLypNv5U+TE16voVHSkST9zEMbLV
sgCiExUMzh7VJJwtMwGDMSiLsE2bsmlv7oGxH26QQl7wiQFdkpDxmNNC5R55I9F3yX1wkq7Su5gu
pKS1g4ofLwZrVOk3CIXN3f3laO877F/+s3WkO4qowgOaVROiUYUvvSsx7Pw5RzSf4i0KEer1lIBc
tDB6AfgXx+V2uHnJEVMTINVq3c6EnkZFp8atq8cfUos8xycNZ9Y0ul0bUeN4iM6f0cTfmBRxF2DJ
bKai6gQKDGJE9t2Hj5up27FWkDd18FOZf+EEXlUl4S0tXwT1rFXYThPK9+vSgMNrOQfxlM4CGeR9
s2Co9ujHOyiC+GoXgucQ7YYvrLT2vfk/l6tZOov9RdQfLQ05Kp/f4ddPY8gPg2l6sg4dEXMZy1FS
zHs0DGrnMkdTXOyCNR4wh66gZCX6XKQdC4JnttN90HUhI8W2wphYaI5nOIzY991kvn5aqGSIph7u
kOTv5bVK50rU/o+0Tj/W1x3oqq4MVjpT9j+ZbyRH0GRIjiO6A5zr+9kAfPWXNB9mG/OyuCN+COY/
B1hdqTiuInLA473Dd6lHBFxqsjf3zQVGeY0Von6VxNshDL6pIad00/cV+18BJhlbGexeSF+6RxMY
fbDsva1KL7P3ZfIbwQMWm9NAXHFxn9fS5zWnYnlVCsKycHOGs59wAQIM41zrRZsM7VTMw+v68S8z
j2kdtYw1cOqhePO/V0wXsgi3SCI0Of51B5K+bv5OH8d/IsSHL1xs75LNmm/xfeBlnLEay9jyk88V
1pLIkyKx/z1wPnVvUfAjJzh4hVDxxGRghSQJlhaEcJUNfhvhgE7rr1/MOJsSybQNAdBTXeMtZytU
O6pEP1GFwRSbYv1Eo5te9sDwv3lmsx2VUgulh0U/AmBvVGV4KNe0afPkHoG8CZOMSZ/8IJq+KfcB
StVJkZpsgxkNIcyJq9vV+GZJ2s7uxl4lRHKt8Wgae2DjZZLn/HMH385Jtj+NR381OYZU+Joripo6
PA5KowU+RJWf3bgDaSARmNz9iU2ugC6RmS85wEDBRgQkbMVSltQYnxivotwfBPfyeaeGwghxsbVL
G1bV/KWyoLf5GueqglOM8dpR0bu+sk9vhnb+xzvO/smTUhk2k36hhf+WQ2l8FBJ7gtcIlktPJw4Y
C4O7/PbNib/vEWqBVStZ1lUIcmkxSvQSYM6kX38VksX5T+8p2nLbkQoCVHK8RVrtdrFjIXeWcEEY
3z9pW1xGcE3QdO9CN8nkbFf7zEagFpxEZgsf0XOJyUIAEOWtkYEHQB+CzSZJQz9vBjTPlRYzKH7+
oFvDLe4GEiDHy+5th/7yMSot2yT99vLnWFXZwg5tZB1RlVnp2ts0GQXNL47wNxEnP94F+nUf70Oj
jMIv0jkjTlGiMuVqsi8+GmIHnQJKL5MDaXN1gQu3/8uj2AWyvb7awpAiVsubxNqyo+rC0jN/MDnz
s/oECEm8RNbzy8lFx70VYtpv20/RLTPz20yoX7KTHZ4dAUkwiSU0Ii5PP/3PYqW4Tlwp2blK9J4c
+pXJTAbWaEKFWZtBv0EBzISuvo2ggQ3SiQ5JemOOF7HJ4pqId4KlMmtV3LijX8UJS4ozT3lK4SxK
nbg9T8/81vxWRv2mLy417Hl3nwPfyckHvXvlzb7QMejnfg1d9ExFAyzpUdSA/B3zAflGLVWID/yA
BGJlm8MT3FFhPZwPq8PD+X0HkK1TFMmkCJsbXgk7fgjBGPNE3fldD9JBIPI1FVypXOlvgYtCAp2L
PT+tmaR0E8Iut0tjLgLg69gJzoc45ZCNlcUbN3YlCe1L5zQKga84M5vO53R3WJDML9udkRBk6yPK
82zerKH0srFYxgb/9DzXvx1EBJ2H2s4KJcr5hYQulG3P9eMBtVKsdR+jB3PSe+b2CK6/5/CS3QCF
xHyWWXlUoC3sBq6bZlaFnYIf97UjFtdhx/we+ZHUs+K4TipzfI1iBN7ZdYkp7giJWGzzY4tJXvUL
Qahu2bfskRqDKCp8/bq4PsuZ817mmukPkpg99zcso3ZzfSq2N/kZEMclqRkmQ8qPsykVg+Ht7415
noDaJQwq0YcchsKX4xzIvnc+LaLeYWwiDBM3GiV+QvHzFIA7+Gzu8sUtLH1HNY3KpxUNr5xhxW8I
Dr8egWwUz5uBJMtvYtMVYm1kMqTQuiI26Pg1/xiBjMOJNUaTw+vIcduzBW3BHHnmSQLwbdvD9sGY
/PWm6uyCOkjlsk+p1jaipN2+nmhfO8Yx/vn2zAQRWHPqZ0h68iJTUBaROTHAMn0lQ8iKW22yv/dH
CMuHVHQKli3G8aYwA0DxqFnHzmfgbaYn4m+KAtDyLRLsEXVGVYbVZ9NH0YcHQAE6tMbZYlNb/nXs
nx2izGpcPFNrAL4gcFfK9i8mgU8C0OaioDe/3KqOmFSjCa+9ZupHbrZvQfVTdzP6kEu2UWWOARyG
ZKEfEstTaLC7W5ko5utWHg2TyX1P5jHzsYuS3kLxsFUJJ6C9+vbMjjWNHgERVtKLCLj653jzA4gJ
mEMReBpMBzilEF3jvQITp2LLJISOCSNXsJVjVcDJvQ3Yp2VQY74x8K0omp1hzSA7x4fp47wKE5AN
p7OrUIhC2AnNluexoJTVpWyPeU+XQrZPaPBjetbMDoTzRqttAfgD+fEmOYJGFxznr7/47FRqEWoS
2TaZWoYUEJZxVT6YLCNpCw6JjiFY9VAZKcRittGIG+IxeIe25It3WImrI40tv1MFY8jQF76F7U7S
qBjHtkA8f2SSKvLshDVPf1RuIW2kDBPXnzeLOVnk9Z0Cj7VK3W07jBOxOlxWPZzAqtgiB7cdI1Rs
IGbTYkGl6MQdHWV6mgCpxaeN3otOoqg4yBONufDbYzQ+Wm7NrxNXg0otrXEW75ISjRkq31YDm/Bk
iMg+wuj29sMr5u/8BUSTXGNWzdZWZm0o7SAkq/bWpdX4BW3ZHRS38xf7HL5ImMPNB65KTsst8ct7
Hn62K+Xc94pHbxA6WQlhmAzVuOQIQVcFN4kw03GA0PigoP+LpWFC/h/e3R5KzSIXO10+eabwMNf9
ChGQG/eo8FdUcHZiU5R4Z7I2TEDsJAV4eD2lJzLiMcm3zsT5BCOOPigtMFS66KGCx2QBxcGL8Nor
dstihsFRk/vLwqdJZ92Z/wIq8mlywc83c2urvkURVwwCnjy4PCwwe3hE2sRNQe057C/4vo9Sp6WQ
NCS33PSJUBAl8fkJEpx+ek7Aygv7AIHJmiaMHe9zOgelfGExJuz55cOAEFPtNVJHUrg22bJKyhFV
A+3iRFEcw9+Oa/G1vYCBMXH2KeyrtLFEdxkXYEPBMzXmqmnWVFqy0Yz0Kz/2YiSFjEQ82misvoJH
MmN/XSijtrTUYpYl7tRDj+1boCoKV//kuYUavV99A7YPEeBujbIpUohVYBSDfgcScDIrSlwRj5XH
Ap4YwuK3R3IoVuSg8tVbrXIYuIK8ds2PBiAggsnHq707XMuKt0iJapV+ksAc69d5wiLI7W7E/ZVg
EM6TJN1nZuD0iIQr/fRaRNzIVA8ZdDcMzeBAzIsgxYKnN6NWkBqgPJ3PXAi0Gf2vCvxEef6rpq6X
PoM5e2/Rv6uN6g/8iPQPZ1AAQpRm/mItbxdeMX1oPU2hmFBZ938xRnszMu5gWYRQWnvjbo9346c+
hzTHc9VZfE4COqDV+K/wJY2YSy7OsK1juV3lOBsaoD1/y6itdWL9tLZqvA1HaCGyKEGKWEi7PnDt
zm9D5YhMLQf4lVBGkxYbIyYNqEfGHcyvFboZdZunZxhfJBYvdu8nv8+skFscvo2TlhQxqOvL4Bp1
vf5OhH/7Fv2nbRxijIMICabDXt716LdV4j1Jj8MJNUljPLyrCYhz2reQfwVlbUzwZJzr9enStfTF
XahrL7QdSIzSvXiZZiayNWwwIpvwI1HfIEZHwhGEoeKWdiNST80tn+vA2TsOzhMnuX/HiuIiLyO7
12OAXWqx7ibImcz+RSx8HslUugr2LNkA0A11YjX+WtDgayCFSLWyV6GPe86QMP6HVVn0cvG3X1fJ
F7DGyvd55rv1/pBSyMtoAh27M5FbZE2GhVzDqrIli+ZR3wC2Kfn9VWagbtOgrueNeB+n6V0+sIx3
QqH5gnMJIN/MpD5CBxHEFh/4yB6+eP0DjDm/+3QDPk38lpDBiR/1MJf2WUftjJM3U1P45GOP2QsH
lZvv/WleecZ6kExvK7WVRm70p32oIi1V9YYT1TTEvj0pTmJskv+yUDhCe2Rnv9I47IrYSPTZaKez
L+g7Ubjk+XWr/v2nTLgg8Dga58CaqWyM1V7Csg3Tje5TMNh69Ls1BBw34MJkk3pmUoXSUmlI6ya5
OSVmp3LizPLxXPGZiao3kRfXrp1v9HaCkDsiTW//oZpmNKmoMgwwJNonNddFPK6nONJIHiCX3gGq
ZrTj5kXdXf0eGHUvvgctYm29XSrgNbT9L6ntB9ZdHRFnkoB2sdVgg0R9ma8HGvP0gZdG04URMN60
nL00Y3wW/sbSmwsUgv1dZCVVjSp1VBXwOqdqx3y90aMoKVv5uRENgn7TfwUAI0hjCvijl4CN/+r+
3NDj3/EGOI7wgZd2VQ0fTcSgysxi5K89ExVo7y1FSMvNjTEQcmSOSUq+Sa6f/HgTaGgju68o5zYD
oS0UjZJMa2mkJOIb6nDcmocM5cQbrmacFhCZu8ZfO7B3H6QsKDjrby8nWZQW4wO+o3tr8FqnCQ7Q
pkpzLzT2mVq9Peq3MGbMG2wjk0spkmSt+jn7m3EySwUxYLRlC5OhRg71wNgRhLONLpfomKpZJPtL
zdOcY7bXdro8fM3tfy7r0GSOIwE1pzzDD+LDeeFFh6wC9PqVwowH0BVSeLxDAe3seaEe+WxoQMyM
ethpcJtVuPDgUN6gZsqs7o0/dwSm6NXCd5mHxSFHrKs08bN+VmneuiPanVHrMuTPrwxex2mKnCXM
dq7xeaePmp7oapGh0Jz+HN+4HJUMPaZ2w4RchzieyTph+oaO6vfbsx2Vbdz2P4N0Gen9+BomkxHr
JfersNCNmXZe+KKOnZxIJMgqwILW/0J2EEWXzhfSFLaNavZ85rMTU2fvx6tprbxAZeRfCwBBRI+g
JaENT77HjUYYDqjBALvH80W+BQJ7oNaQCkI/ysB+YPsYMhJH3JBSJPFKsIpX5F+SL160osrW92eN
dEp2xVHxEPAuy18gQ4w/+REYfdAvWbzaGKFnLXZRpJcxvnmHSGYVxBq540pRC8UCX83P+aQ/WvnC
IVr6l1e6aPb0kmJL05SQAqXfYZXAJcrn6nB/G7HDVZaHDJsOz6cTzqq/y3fO3ljrkxiyH3buqnzE
TlhSjNrpCbxPnXAb4Ztw6o1C92InodvcgJn0VrcjBjPPJaaDsu1WvXFQjFo97XCZsFP/X1nvFeoW
iK4x6NRQ+NOnkTyeyEn90pAbaLNo7aRr/dxUWqK/Jj2gCYa//yO+uet0gDFpSQWZ/cb6TIlOkWxE
80fSTs6oJzfRxIrZAenTUiUvaIOyxQfIllPI+FviEHrtas3W3bxTgh3JCKwGtTMQyVR2aEnR/8RS
ZOMolhUs69st0zKPRHlDyoDQv+QVV4T4n0e3ns17dr/XG4alPu5vQvg5y/zHsF3zzGHeG3PL85ce
ETMTjwgqKCZtPCxc7XfoGR29V8fVkBpjleI3R8BcQtfImGsQmCtfs/dZ0LELVMo2VScsV3gGZSIK
pOGqzfJaP43uGFbY8anUKd48peIWjmJqSu1shYdToPiowSOdaj26eK4LUyNAdPcNaglCtI16Y0Dp
mLbcNXcyhopR3rJyZuZp4Zrg4h/scENcmXdkYsMdqG0vkZ36JRSI+D+TAGtaI3EteIyCTFmXdcpI
2+IVWi99PSBDaaSvZzo6flkopHDWAWty7Ab/YQ5s/XHfHbNM/Ixc2UNlyfMWro7WZDhpeO62EKX+
uxMm3G9mIcZdzT7u+UxlWT+JElV/LMgrtFg1mlHgOtzEHYSMypttUHHsp21uEXmkKnhRr5k+fS4s
sZ8gPeMBG842ZzKrUCASPBbH3DSkvi7e7B+FieqwGF73PhsLf4o1N+EeJK40HNZ/jRMqjIvIZBqy
70dVYnxD8hScbh7GaAh+CREzvxCQGyb/FHZ+3UxoVBvW6IzeN6Rqh4cz/TGT5YAB+la11UBY8T3i
tNkywX08JLuPJ/XsjLcXMeygdqz5wl+poLODCIfLVvUeiQ63ZVDjTzAjVr2yw/2nEGp027kv9DGM
NWAdtm6JxW/z00FUiLxoR8+uo/9cuKBkeVu69yQfY+7gqt9sqHV6OLNH5RbeAeoWky3LV6n8h9qE
T8OO4pvJyLRe0wOUhHTJIiypk0RWgW1TqZL1PmjFhx5I1Wmuzd9e0b2p6Y8v+4xeApz+SJDbiYXG
WM5Ehosc2RaYeDpvKLzhJnTt2k9x+Co1J30ee64CgUN4Rh01bAVXiYymQacCqBhuVVAgr8J2CM1W
uVnBGullAPUDYNi4NyVCrqyEi6kLrboKqIDiPQrTNLeG3tINK738u3+bxS1MZ+m3yQCF/3IJvYGl
MUxspBJnDYHTEI5ii8LugpwENWuqdScjf1JfM0cJemx3Gk/e1StcZFcfmUQYIowwIn6QFPUHqAzt
vEXUJ6cBaFFBBXPnmOrCNHoslr3M7XPUwaoaT9B8Grvs3HmActAKRwZDS/9YGug582H8Qww0NLS7
+s2lS7Oq4uiZOsYthcu1J4W6xqBd76oc6drPiEvZPFnUiN92RFUlOLbTDVh+5Q5nM7peqg5MHobX
IQNw1WVJhiGCIa2AdSQjfvLZMIpi1gOtfqBiQW0NOruBKjWXaW9YVxVhUCtSDQUBHgYAYpta57TK
pInJKia+i7lu/uV4HnXJ4xqKMqN2RGmgH4y2TKIBxBvzjy68zuHG9ZDJxFnaauR5z3N2AQdsO5qS
borDFHRF+1KtMohXPiUjtCSwfPlOLYQCtOyBJqAv2gvxyBvh0f+C7jeunh2sxInwA2NQmqYmPgWX
/YPXliiuRMzahMEDDBVaQrF/x5+NpjsVw8AN3oz6nWfMBxgEWNsqZtnrQe+i4OBBYt/ZMQSHCM1C
toIWnKz2DSpT8+0F0Ds1cXpBin7EdKM0m6/ZqpKomq3wAKmCDhsJdaoqGtHcfCFJYuAOc6Kv60J9
Zisz15UKmHGHsLX3RDowTbW+ORagLunrrmj/XeclZFaeC/VtmW00zEGmq//9Dkby+A6L883xorKz
j2P+nlzI8Y1kKnOD9cY37TAo1aIvf6Vj5zuwLAkaUUbD6VHLIt7DVUWlvI93MlGEVjtosqSG4KkN
9eW+H486Ny6UcwnD+SWMO7oIjVva7XymSdhCiByy/YLMgI2MuxluILtdoOTX656QFEkI0xtj3SHz
fnOB3xoAz4MEehS5XCD/PMHhTaezcjudHjc5Tf7fkTbAFXkO2xk4Css2aA7tt8tTLkqdUDOEy5QR
MUqrrAGltzTsPONxW9XcUWKeQmoarou5+xUoAc7tncwoajSZTuTgNUXbxtPO6XH0SXyK0k271axc
g3DFSka5W9FX+KZzuEMjG3Q3RpUcHS1Dd2DKgYjkvm8wDFLSladetWNYsTrV1dxh01VeWdvgxZk1
ugVy/M8Z3vQcxxq1gniwDwBFFdGS0vT4nqYvwJV44fCkUzJmdccNM4HDc0rBO6GqiQvswKLih43u
w1crRi1DBOgC7S+FpxypY8CGp7s74oK2kw29zoD1N2Gs2EmKz6tlm/n+nA8/Zqm8+/tswnFCvOPW
qpJBesJ106OggB9nnj/oOFWmlfEwgLsZUKxV6gT78n9mF6G8auuLh9W0t0r7D82RnVFnDKUv46pb
v/BN/E/Ng8UmAkSK2GCacOf6koShp3E0hH/2oSwaZ4XNAkY2GBJ3e13g6yZsFUQzR7op99vOt6qR
cm6yb73rtQGXASbRwrbMfTNJGOJXZKaoa3Bxre4NmrZXhoqZnQktYfY0nndGfWuYbFOoyQnhVKF1
d6DLuTStn2C8d/cMpEkT/U073bVPzUFfysyN/EWNOX8eE4yYrYJmnhwQgZCwY7CEWzvFg0gabDq5
Sscr5LWIQk3uIbLvAhumbyNVEbtJCB5l0LgaAtf/no7d1ueaeRxHBx9ROhXPhJXfvZe62O18hRNh
7vom+l9nnRUFGA564Mu6z1zxrPlL2NR0SpYFL2DRDSgws10D+JeM0zDgWdgV+UZWC6Ly7hJzKWs7
LrS4pkjvwZrIAwKrfRwNsKu6LT2bI4pC1wUuv/tN9JruKISzkGJml9DPYDhJv9GOy9oPKIWEXomG
tjALZhFrVW0jIdUN2KloLt59Oenc9LrajS1ZkfQMHIL8YH7KuBdfvtcSUHIjugJyLBdoW6NM16+K
Kq9gxpwawrGsbmtHIJBopGJyRkEpP1lOLVlG2hbG9KYDLFr17gPdKg+p7orsEddsi/72WowCnh7Q
/WktJFssvNvrKjBMeWhqISqODGMFkX6rAK20vgPsPURDGktibcJkM9oUZLXWYnMHUXl7D7JULpdZ
0dh6uC3kreF5u+1ObgTYbMglWlKOjVNwFLPnas03ut1U78a2BLysKGybT7MiAe1YBD5EdOSi7b9g
MWqd/qeqwwERCT1SYJwi1DREnZa/o8GrVGtQI8YSOT4l68WiGdLl8XWYv7VMB+bk/L/AeOzj77rV
joJk7nmEFaUNo6ghN8Q52DIbWw8uinxKXKaZTOLbnJtEHcvmyJ87RxRgfzgcMSmLYt5lPHUc85JN
Djq9KSDJRAjCMajiv5uXKG6mUzSc5L6nUCVYLcpbBwNuobqUbedCbDA2MrW5CwEhPBFox6H3xwBe
jCQ5nVSf9LLvhCExksn96jGTCkUm84gJedP35jKv5VNmYlAvfrjokKD7k27nZkciXY3Q4LM5HlMl
atduacn2SW9QavyqVAsNwaAO3DhLwkLCViPl3nQVA3yn4KOZva3AjCjsaa1/cGgmM+cfqO9FtsBU
jQMHsva8EPVBwMjO9Mzu2ll3CmnZST0dgHAf32HA/bYwiWlgNwR37IwZdvEkbj/prj2TQIceyp+W
YWd20Ba2nRvM3RRpF784xo4fRAYJ/qOLf/9fRozTlhe/XZQjVfIClNwYVI3hBbCZCFuc2XaImtQP
L8cImJX+M1NeqVofWdtM2LviJ/+w2ovf2cWrnoy+bQV7doljmpJG3JCn6fu4X2ER8Uww7iaZq3z5
e3z9nenEvkeJwvJBK8zJJGw4fFXrHYWXD0ohBFUWpdnTx/J3xurMXihBhmQnkKx0rUK/m8I+/N+r
4DPhmP4rSaVcgAWT6hU0GcA/tx3ukwIcYXyu+Qv5AP790pMT5EvEiLhk3NvtceRyZ8axDVWLRuD/
mgKpIHafJ94i1vGBW3tgAE2URk+jjApM0xAus3Sf1E+kRZT93W36dO3vLk8rC4S2oM6FqAxZLpO5
LNjG02vAbwguue+YFNA0ZbyaMm9UIglK6JgoFYf1PcU8q+Qg0ytzfzW10jG0vImviRBoDb6tnJcI
QEQNAl5Tj0wlu9a0I86Sl8IgIflqt9ajUVwyKn36HswkFgPrvCGwF4cYWbgWlbyj/2nrqAf1Ea9R
0ZG5WO1I3L0Nt4b/81Bb3hmYNmn0N8GwCKG0FViD/ihJPOgcAEIbWWs76FmNUfJMsPPXtiYFu3YS
rMXIW/QLMAeY+7guM9EKXYsdY9JuwnjnXRwc6uPGlTQ9FjZyflkJ5zFpUpyTIkEJtG31Wl8YFbo9
ZIJl4HwbhCsRwYHY49w6HIgT6BX3jlHcCb0bJeirGNSL0K7e/mEdMDuKMqf4O+WszrmviLQcgO2H
GEq25kXoT1YeE+zZ9dEkiShG9EiN5tBjiNdL5mMzU1+9LTHjj3b0L6WSfpG474vNaZVYsqA5auFb
So1DUoWX0M5kXG/hFlUCCqLU8Xuz3L2VLZFRBdcqAMItFa6Gfw15zkQnqo4UJ3kuRIcHU5rZbjxw
5R6yp15I8sKGw/S87/Ugq4hYUSt+vP4lKy7yFn4Pm31h3kI1HM6AcQKVgy87XtD/Umk+Babv2cCj
H2F2eQVNk+Fbcgtt+c4uofs6PiywIH3BJP+FX7k/EU4V2L2fFuBgRbpmyF4AyifhmqO+r6rIJIRp
+g91XMjVhXC8hc/K752uzH9eHRdnAJiVRbQ8AAwO6JsuQw+B7AILnzJjZMfQnl8MfVYQCDXNWTKj
D35+ldchHIco0tiXFLsSWGcp16+RYWoLXvHr+R22kkK4SYsOov8abP4FId6WH9QJJ2oBvdEicru0
XpSK6MVnDCICrbvoTOcqPp00q3K1Ax+xqh8wPUFScwDtaOktDcekNaC/F6QB7Klw6rZ+CVwm7ous
jEYJhqyyVHXI8++F/XRSurA7yfQM3wPkPsTZwCDiGAvO+IWZZIZAil3VW4D9bBuR5lJ8diYkU1ro
KVnSnSYlXE7ctdZj2lWdXtwHJThYFtU2FrsuJHUYxJ/T/hGWqJ7RT37VH0xO7dZMszjZ8Kuvg9hp
Ij6SykIGVxsDlPqc24g2bzMI4NrhrtxRN+vCgOLhXoGWtZHv9Rb5y3/KREC1SKmCjDOFC2LV0rYg
cSrM/SqNc9dv7s/DLEJTxNjiZF8GjggKWK9u8Cp9oAPdpya2fBuXwBni9m39ccY0+0r89ZDWXpNa
5Pzwe/ytSjjlfQcfefoLM1LrWi5rH079wQ+aJ6+cyDHdCxxQNSlpUP+8S+KrjRbvIsd4lnNv8L87
9UNBEhRvTzWleb1Lm0kPLdBPsn9UyniDYCqcwvx8s4Qqon7UY3Dbyr1a2M95+YYhTgVkHyB9v93r
ATetLRNtkNiBIdK1nMO2b3+zwHxN2H3r2Fxs4/OWuVh4G6paYptDzr4nN81VFCFKRxdD3kU1qXih
ABXANlhs0PZKKq7EIsTKhhxy3UYL+qU9NqlCfe8sqGTD5QoZd8HtgcIKAcWFhmEwfZFa2wFFiH2r
uQoOsAp/DMvazKbcDfSSVUc3eg/zqV0+FfoTObC0Ex7vieXk709xwFKEYlNE1dCJHEkC6DelSNlm
0L/4KTJQJIWFdxkxkDrLApgjHcFCCOFUilW6iNOAmM6pB328pT0E1Knu7lyy1nn8NKdcIb4wOA/E
BNaN8Nn64lrvG/FIeWtGIE1OTxqVO1B/8SC+37bBv6sQ91teqNJN20smn1fvsdZX5oR21RJKOiss
aUR+4LFna1Is4WeYKEhAdE8tXJplC/vsaU7z8yQRXHpjvoYYw32EN8gajjYeEDESMSQdr5k8PbWW
CbSY4I5R4GjMWyeXG82U2OuTdU1EsqyZV5JS/B9l30yHKZRcn+4kl+W7joNcedJrL6kwywKoiWya
1L2yX0pIK5xGIZKV5p0JpNsd6j+4ebVnaojdEVs9qvnvBExUdoPg1xz/SR3QOAMNkzOi21JLvAkd
qNoyAU6KXt4pTa2Ps4IbVBInNBAm8hrTp7MRa/a9sMQDTuiQ0/qv5E5Xlnx6D4HO49pxckDksI+w
fQpcY+llJ/Gr3Mf2xRfUfy/1H2uV5zV+f4EKD+AvYqXQG7j7EyCoQMz5wzo90ddC/SSq528L8mMB
g+XzsbhsHWDa7/LFN1dPgEGway378/5IkPXUFP+WQk52kFMqH9BuZrKDp8qmRFMIH5g954w0oH2g
r08b7k2OAfTYuaipPg2PTTxh4lCdJsKxkFNrgLjio1AtZtCnzp3DFF/o3CjF0sWOPPyJ4OBk+FFl
hrGzOCvYRtlfCmcKTXNdERLzOWyqGHcS+/QTtac+nvRmOj4t/cyu8G56doLIrGbjIPZeseSyhQa2
LGGv3FSgW7zwIYeANg6v7MKVmNBxG7YOUNv4D0xDUEF4G5L/53rGW2Te1an7jJ1ZUUoMxpu8ePkS
WXHj7kLmIl1WQM8t2c0Z46Q7/uSZQptTvq8zRgF8/kcf6I/EqkbMA0dwE9YlDITDRBKOuvnckXAJ
7bZxkpNJXCx71eWUeSerwKRv38EmIgXh6RSP7gdZlwssoAeF9I1SHkmV7Ik85vsfzMjcdOz+wdhg
qbgGe9RJZCdXHtEqQVz9Xw8uEcyeYlZLP00bwLV8CTd/2YPzeQK9UlUOw+BZOZUiS1cwPLOwNlLX
pBxzQKVlkomT30x+B47VyBESXgtGus92gdeQzVdQv0svGhUPs44kdCbeqqC2sab5e0kg4zauFyfV
z/LPuWTSCWQ4bDqb3aBiW64ic1Oazikb4BCHlYQ0gfAW3eXGKtawIjBXSgir6hbKaQdsjLsBnnb7
nFyr49zkvWIb5vjecOyjS3p9jnu1EX7MX331jLZXRFNLvf6yBPL8jL1I+S5HVvY3ae2S/dh1nOaS
5VUks11gBZrSTE2O9S83z+LQ8+FWOKTp0ooG7Rj+lNRCvxJ6RigsLDHuJL2t0JGxesxeWEQuNBMm
QVNfueZY3UGhaRK3o6+Q6bT9bhfWW2SIeg6MY3F3ma00gIRG9NJ93CThWoeDB1lEOCQ5LwShvjrl
qrZvTrPeknMrotd1xXIj2rgDImg8TmQDHe769noebL05WXsvDx4QgEkskxhzzvmmIlcuyeqUVIcA
APjFwwgmosIn6/iLI2V0ImxobLSrMyl78bjyBQ+0fJkFdaEvEHL4nGmjOiyjwHEn/PlzIQ2yTWrS
v6bpm6rFI6WtO0Zh5ecQ0fpcDKs9iUIqDq/9nIYGzWXPswO75nL6+2twqKrePY7QAsbBTYn1EV8w
+/OZIMU4rivLUrb/2O7ATo04c0zR0IW/98ZlzOHQ3qP/iZRgnQwn+99ieI1qs6ckmJfxOOJJJe3r
l+mIeWIuU05JHhi6yfnV1+FZ5/FqTKpA+lVxAdhLx9zLzRZ0XV7gSVU1DxuiUwdYbyOneu8Nf9lI
u+bsE2SbeKarfY4WMOzgSvz4dIo01PcFR3Ixozi/9RGO5M2CthqW11JjOEW9KlFouMaM4QfOVxhe
pRT6fWzY6/MNxDfYiP0E7Pnji3PeJp8XK5qh1zkrtLNEKYq35rnA+DPAr0Y9QYXN8Av4QRiHOMQs
xNiDQ21IazvxDalPE7Hc4x8Miik3+H3Ay9PWoY5f8s2YwqTfHVTMYc9g9CLKgMAAEgm4gy+kDsEP
ZFEtJdWAqwBa3sJcUIBtctwDCwaf9dSmu9tWZLbd7NDQawXjrMNFclFC1gtK9OrWv0eDbwjezClm
fxQvtdW01K1pV0qnobXgmcyvSnKflW4io0Sf+zgoj2MdbZ5reUk9YYWIChKUZfGwli0NhQAVCm4W
/UJts6Cmy0TE6Z70mnkC8TBWyIxzvdC1YUKoOZ7GrcImOTIqiLnnlLQNzLqtWR+bijUTFy5h3LO6
MqvJ6UtYl9IMJnWH9tUqQjSIFHibC661YY4NeXCZz2hXmbE9H6pd/MC77k+lnUferfy6wrlHLuNS
gbLANGO3WIJpoRs7K9jTFy+0HuXir63qWl1nRlrc+qagEf82ERbat7VuTSEfBipq/aAAJWSOxWdW
wKlswPHP7LlG5Rvcj8p1gEq4c+H/8TjefwymEfbuNTXOyikSjlkOly1jsddHm8Q5fskUwd2pNmk6
V1rQann/MD7RMw3RNV8+6htFlQwHqbnIt03PiEsgXbfWcQKikRe1lQ8jXF8zCcbd6ZoBUm3bFu5s
hA+OsJtH9reZAtoEsxSGy7zDSqqBPXz5txTzY1DssO/G7/aOUO635W0kWHXTS3qggJd7VfXCQRA5
2X0zRNwr6pT6ze/dToOeRwLvujJioU3frObMvRXziA7+ilJWCNUdPzlGio7rIkkHXM2QfSrWe5jg
2fL3rpNylf//CrEBNFBbLMBWSW6kpPfp0hIboBKO0Gt/tlCZOh3vevwllFeBz/VcEI/fQk1EQjx3
LjPjgtm4NvDcNKisz5/5+QiZ5I+rYpnm5hLCRpYdO5kL3hQGC6PNykHEXW5ZCffIhOgNlDZRJsrj
apiliU4mi1E+veBt3S/Pg8Ed/P0otp/HABInzq/jSQkdVHE+0rovZGJA6dpXkQ2YZUT96CYjAiWX
W/UP2VvLMQBQhJI4wOp4Q5EvHtFsy8DU6MKilSUoZdCi+D5V11bkA7CQEE7JYdLecC3BU+1birkv
X5zMRzUZ/KsOD5kIf4GUZX9Kg1bYoFcEZTsacj4IUaqXLHA3ESmAL+tOStpg1R8Oz+WpJ4RaUG25
AXJkR7+K2gq4F4r2Q+OF8XruLWIF3F3Fe7B7Bl9Bw8YPdPUv9gUSikLibwrT+kWxa405+aXK/uta
9QI9aV9C66W6An6zcvqRKT7MaNen6jaaJEuZZ+T4ADegQNx3bO3m7/cpJidpQu35uAzF0rs0fL3Z
/ayAYBxQ5JeMdsyqZvm/mByQTY0kCdr2jjTswVmRZ8mrhWHry99NIJwHorsjG0o7SWRu25BnIwNN
TM/7YrbzAPTvteDrPUVJ92ymI6qFTnbLAH+EWAxbpHyJ257+u5Upn+SVIKr+jLnGWzj0AxgW5Xfn
7uddXJg4MCqco0M/HNIVLQjoTbXLoZLEHgq/UjJxrOh9RXcjqfagrWtIY9/AfftHWhM9Og4Xfd7V
f9d+Xd8iZKImzVSbifzEEQHLhLBbFbtR6MxtrHNshHZDNJafBsTxSam/zKUwh/5L/hV6pBXL8mgk
RnW8LUuBxJ22+7KEbcZZFfAZ1MulhlH/V+uB0kj+W+9J97URrlwq6syTzOUzdySs27fJYacrqE+Q
NiXOwNhruhiM2TEBz7LffVY3ueQHOTrxRh+hMZgLy9yBrXqInnXbbl2dYYtzffXezkBIGwYytYUf
e8TnpI3svqv7Q+sAWbX1rpKilOEuBfXameXeZY01MKPaNMt6WONQc9u5hdfGvmv3jcFug7RPT6Gw
S6ZdNve5GrKPWVJdBAiVXqlMzofZCEsazVwTUmo7v1hTBKOf3E1aF4i5E/y2VfLVfopfEMbceE09
TtIGKk+T2TPsyVDaOPimkTMkycZgdX2pWQr7udnjVsWi7B+SyTEKwXcZQsrT5X9Zc4MQdoxwqQAN
LC9cEwrKZ9cmOWieDeb5ZMPqnjTOh/CMDvXERLkizGl9NcCFXoBSBipDVi6a0OwKMsBtMT4ItF/R
42dmVmHKRr9Bor6KoElZGi3ZFOmoNDrwaO5ETs+1eBH42pVNSP+A69nGWViobD6rmmsIzLaHSO/T
zI1FDujqkZ11bhOOJi8q4FOo58V2QKqJr8nmGovO2oZHJmhwtnMQdb00xtWV9mDBcRjzLcnlE/Mv
GXR5/Uhl/jHi7ZHPaRntqc7REI7Jw/hYEKuKkTHa8tptqOZWy2lU1AdbIdnUwh8v961xyzFLybUX
jmL+wC0rdEHP9+Pv6UZrn0FJFW077Py8w2W5gNiuBi2dnor6Hq+U9N46u5o/taK/5igzV3EvonGH
hVzqVlntjIHzcql4zVn+maH+/KBgBuJZX3Slj4smdiOSjRcyqQrkZDaeDN4uRyXSj/KYLFxHvTKL
iTrVNoLKFSxs+LtwZyVIj4VknjiiEmnkqo2rl9nHi+6VDTI02i2NjTFodWhxXcOOtXBLplH+KGP6
TttvWa9jluDYVKDztUnOWqkG9rujfqeZpoYZ4bSLjn3ONQ1O0szdbUesU0+2zmiRppou1dDJcY/r
C18Qe87QEsJIpPzpRgD+RnzkEuewH6sFQ/mL4nfphocZSYPSJIV8d0TtJXa2opDGMUrU7TkIQ6Yt
UhKNsSIF3V4KOovnMTn8HJOe2NClgaFkGCPNx/uIqpq98iS80O2+upHK6GISKBIBQYt0p+DGkys+
8mz9GP67M9EG6/Pp3T05TAT0KoV6mZsABHcp8cUFAQ4+SkFuFsAoUZoTcZDQvsNiF3fFUjcZMjm4
MNKxt6hbYQvFBsp3Srm7XbEYYK47JO3uefgm4j+A4vzZ28HmY8iENdqH4v+YAIZAWJcUF2F4tckt
paKR0XtlHLtTGz5veLIp39Slwg9JjbABjFsd2kWnNySP/E5W9E2cpm9GJcJlYrLMJSM4od/xRw8B
e4G7sAc9e/k9AQVtZ47eJ1+XqehZBC8FHGn+Qos1piSExcKIyMEVD+tRXKcCkA6g0+o53QgZMsRh
aJHHokiblNS/O7v//2XUoEse4Qkq33XOsTbymN7Dr+mtVFAroOGVgPcDzuLNrr9lxouK533+Lfh3
9zpTvV88aYllyZeeO/KN++Ehf57Eh4pFFLRyZR12K+Ui8JyG4VS1ssvdXib2AYyKs+DxsHOFKsYN
NVXIEC67xgLQlwZAskzgTJZfTnW0SR7kV0U8QaeRLEb8vqP/Dggj6YD1V2mRS740m+FUZV5iIsHY
mkLOcm9fgjDDJLLxzXyC/xMvbzq5wxjdS4a8B9pQQom1eIc0+7MjlO3Fed3oiPxPW6TLTGF+pXft
2AT3iNSA7t548AQwlV4cA0tCciEw4adCPiXC5P4mJ0j6eSocihA+QlrK/P66i0HxWrNGa7LODzS5
ZcLbO5hJ2A2Yo9C4DZVq7mc7Ud9lJSevQTLpGz8hK8eEMF713bxdMt8foIIZQ+m/nWIc9Hp9/OnR
IfX1MNJqyEN9+ONSJEtT7Y9lnRLGifgXStPUvSvG9WI03YZS1SfSOH91Yaa2/x1gK6gmwN6okZq0
rRoIKOe3UqKbZ6gkLUGlwnJwEI2MjHNqsRiEeerU29x2F+UStvLxBmxOEbdK8cGeUNC6GX30+Vd9
Ei9lioLryDfoqwWESbcpnBoZDBSHOHlm7vFIQm3ATP1pHVTG5ov5I4vmFNzsx5YQiwD9vIf8Wxhq
lxRczFTiD3Hh307599U3uHZ5tQhfkuwkGYIsgCYk3qGkDki3WrP0E4FlruHb8kb5c8Z4DFDjiauH
yC/8ycjxBHsLAJsUGza+krwfidOLLyh+xtm6S+ql/xHcf4gbfMR6NgtQalxcvOGHbJArNqqVa1Kj
8J/3tMFfA4NCB85lH327fi6Z+I3JcnjZP1u6VBWd1imAtYsKtz59WP/dmoQN9ZvyagsrI5LSbdNk
zkrvP4QHxN0vQY+WmPAz3PF/ttUpApF0m65Eko6CnDCBjeFy4N7h9/8PJ+LR7LcodHh05afdhilF
R6ppfTekNXvL/mqgme9S6VUgC0J+AIfEzB3j8QXz914pFP5puQwYFlY7enEgfRsVL8dz5HPj+y7t
FBUmkjuNhyoHfPdU+jog1kl8rOBjaPxAqdm+pekNiYCVQ3mkEcN9tWmtPXebq6DMUIP/KSulByw4
pfIalqeqHehNfiUdaAQ0qmHQbFFVkbFHf0MMHzZuRsXmpSYaGrWE0m//DFV05E3vGEbH/Nuso1UA
9cKOY1DGZbCV+qC/21mV6xku0qHkBUj73ImdKz/blsZkD3KIp00jP06Ddxk+HnIVyTAtM08CP1b0
uiSgKq5vEKzI7tT2qt52DFHR5/PsBb+8mmqNnSMZ/M316Hu0Y1Q3tBiUREn9KW++YbSeTPNoAtZR
E/lkQr1GD02NyBxbQfjYCOATZOIH85cQULt8/tMfDnneryTHbdCshBcXEp9gVot71mcwWl1RLULf
wZy6tGdGFuWuOeBqGyFQ8tP7quGSFeIulWfR4HyspUdw2fdQFn/mV8edcwkH8XtQrzgpz5hA/U6K
T1RmExvF0eUnCQnfK3HLnzmXk5DGCbFEog3gR7OuzsJNkYgvTLLtetP9gh1/j04qidOhNUC7Ge8A
ZYBPPj0v7O2ZuTaeVaJW9XREF3lEQw+EIFwmWvqnIAPc4ZARjkbQfEdx5M8SG0Jaoql+9mA/jTG2
I7uV1UVY1DwPYqBa3wBoYanDnBG3o1zFZS+rRHSIVWy4DZY075E1zCnjis593EJycVYxMxBBcoqS
/8Q1G9bJx4J5dAxPK0aSU/TxL1Vu8wUt2ppJ68/uZTaTgOCzUpPY0yi1JYFu/euXSjcWo8we0pT/
0gCbIkAfhJM0qNv690F6sL+5s1MLfawOK4eKwf535LHP6HOga7TIqsHM/sk5Ahg1WdDJKAYGr0YX
Twuxaefe29XlO8A+TFXhmNsmg2LSGV/7tQd0Q0Y1cOm0ZVAtYBBmEnLTo370i86vYIwprlFD1xSe
rok/9r6g3rs8OC+fwEpBJ3Vt2mfhHOOU0ICOTET0gVeJytv3U1+TTn9QbmgiJL7Phc50/WB3zQ38
s5amQRp80aLR7xo9tWdPR2zIr+ZVz+ekhztUyHQ/umcKT5tLRdIpFl470SA8Kp97RN8PhS2vXcp6
av4SFtI6Pm/T5+LcAO7svZ++lG0zQXTgCM2gfWRyNy/Rc9HzawuNir5ulX4+vi+DyH4ceUcOnPul
dBFCT6YL1O+DR2uzLIXY4t9HadmTqtwSf8u/t3m4SFDg57k1QemMLAtM1KfV1vqQQ4zObh4rEss4
BKXrMiT3El6yUGKrQsPDSvNKOACRFvCQYuFerNfbOXCN8r9diYiXO2Ax9bzhrkr2tgsgUbgkGJIV
BMUzovt2zPXv3f30wW7onSzudr+2TyydLJyNUv2NixaiJOnUiYHcrRCz0t0CNwYh8KHR8CDxOo+p
nygElgUqDmzifjJK7J2qip/hI2pOqrt8dJ9lwR7gVwGfNNg6YLyhQzn8983q3DmKyd8u/bHHRj69
wbHZ09hV976lpL7LawCHusapTrS2Jx/ZdF4hCn9Wr9T5Igwdi9oGogbTtPXiDuBbg2cEK7umBXtA
fyd6ubYRZQHtvTr8BwydN3LPYvrMpq3/wQn6b4o7aiuWXBHn5kCOviTetJ7XuT5ybeFpOCtvx5iZ
5qZfL4r5h47z4KspEAVEZu2McKwthXC50H3Bk2AwcVsHk1Tm4yyTilkjz8VFTZlxKga6AYR7lHGN
EosN0uNpowHUY0rviKJ8FJ+s0HQLnHMhT5HIa4VpP44IOA15XVH3EvgQYAGFc1P06PuGJRtq2Eka
D0SLpnBN1aJrnmvEDCivPvV+vxPuk6yuXi9EIBwgcZVYyfGA3nSv8qFVsA9oR2jOq3YyMC0TEE01
WkFnrFsA/pQ5iYNXhH7cU3aSrIcIKH8j04EGI7hmuEGE/7jWgnG/F57zroXCl4DhdNf1v8sQ95Y7
v3ePcgFN5xxYi17r3Aohn9TB6jNhdf4ic7LlOGOoKQm+keWgvALABxPLaXR1VryEHzYiDXtuTHAb
SufxIBEeLA3Yz6+upBLA6Y5hqCVn2h2TrTormrrAeE3/gz8WvlfhzshJXBzX3MlcEe4JPgKv1+lp
X+CAt2o7KIo3TBz+99EA1QCLsiXgmeJxQxAvnD80A6NIwOPPvck/7+EQMNE9lAfzgAWphsYQMvsO
G8x+rKTKmKt/ly8OupCxH+snZfZSHAX3gcr6+1aWyOuvi1xbZx37bqP40GqPUSU66mx+4DqFo4vV
P4PHdnXHn/slBrUcLWM+IjsNOc2lUKga4Pv7AVxWwMcFSmPHR7JDZd44bocaVMVnJKc4nMTV59Md
icnxIZoRy+jYTvdQafvfAnqWggfgC0P+g5QVJCj55aYqOYwzwvONbjeprioPKptrFhTrCRRv8gzW
Lr7WiiNEPQkACqMCIrV20ved8nKvJ2AAVSicw1YDe0KvvURTbh6PevxQHQNeA0Fy3BEdKsFs2j+9
VOGefNyzCF64evG1RHBxwjLZmh6U9xQFcwxD4wLY/8dq4ec14HCUnacVyeV5s+VQ+thnG0sRECmO
k5PJPFqJYsJAXsdFiofkZ1K75I1nZzCusnirGhbGWxi4ovI8E6T7/FHDr80O1rzcW9Uy7NJydymE
lLNp61my239Z3YAsKp+V3UBfCHaLau6Wc4t9QbTlUTj3TCopr7Jg8j37mla9mu/YFRkPLRGTByJx
psN28VzXNgZLZuvt0/leQBKhBaH1CPBrs4hp9Y5vvNstU9vi/Bdw8TOJPazo1LKy/WIR6UivcGDN
GZU4UPfQq09HhOXAyskE15orjFzw8FeLMUwiQeg9kdQSQuroIoo541ashN4LAGIFcUIOwjS580CX
MsIVaCCfA8OLvESRvQk8pM05+KKFJh5W/VuKOmmt1C4lfvYU4uau0FlDrZE8oFO6v8mA+urk+aP7
ClzHh2SItZtJ6QUiWsX37/28gJoeg7k3D4dCvNA14JTq2ttAughI7l1ZN+yH4nbE1OR8WS7A/LZi
hRI/WPjwcE7O/HyDaP0u0q9yTgsvolJKHSKX+Fxg6MNAs6jAHAy2R0J+AvVhvOBmAkClwj8XyzWw
sVLshEF87z0JYIZkDAkqQgCgBpMXpw4UsoCnDYipmuTd+hcaLMj/0Dxd5/QPPiVYwGzr61XZ10Jc
e1kHixgiwNk4J2ecfq3f8jmlHntyloOo8PBq5zJyC29rWNfDw/f2i5rPj0DPvU/xBwqYeiNi+Nw2
1AwWFMho+Q5m0YFOnek8Mj5/QUHnwc0lSwcex4/+R7siYR/wyVADAEJFzy2mQNNxqEJeWcPKHVm0
iHEg9Hjs3Q77VCCJwlf7dzfTpBElPYjbPqXfB9mCe56oxB8xXwWMv4GlMYZ/OimlsaG0V8vGsbzU
mcVMpJCPmv2La7eDmiDf2mQPhBv7sxofQHFRmjFpbK7uwFit9vOCGZZ5fB1NNmJIEtD22lfdAQiT
cu35bR9/IsGOn8yplJYx9q7pqMkSz/8LmLyJXoG9mAUtXRGfcwQqZJaKWA6OeI+VPw5T6YAa2R0i
zAgYQfE83AT+sOMXsQDfy4RVEsgx5F6l5KLHU1Kzynrp72Fsri/gz8OLnxPBbiDyoqXM0YfCJyPN
FEJc+qC7yjykMAT7nzblit0mnZ1z/kqmVusg/lpIU+5RbjybVB3KvNweUXduJwN90soP/8xZaPZN
+T5UgabPMHiynTR0mZIcvWx4wfhzzjv1vLb14GClpzGuxt8EqghU/5lPKDywwBjmS916OnJKUuF/
NtEikjf6GRTnd5JxideV1YkFs1kDp3J4yKm/5gS6jqQNwQCs75ERBtOkc31EFIvsOtkiHHAWjifa
pCyl0DgWubxTBDxvd8pjP8p+wYLPgDfnbgYeMnSJWscVtrAwdcREXDFUn+1Mnd01ezrtLWVa6JdC
nhjEcLZXrte2HBlsuYgiE1DgULdNqj9iTH1kLA8S6+OcpnpwWpVWZA84rmzUs9ZK3ZDi9AiT+GIt
kmH/MRhOOZgvOoepgo1EUZfYh4SW5+9z03k8KMAlcqTU8W7t1ZWcREzdKXxow5D4ALrlJ9KG66Bq
aVDDKpD1B5JJ52Yi5ONvDDdTIoXee7w8LFc9WTwmC1oU9bX5DS6iW/E4jscSt4UqIs6YFAbTNMdl
kbjtD7B+GZuUiqYAvlHtFd/4NXyTIwvtmS/um2Wr3XiTy3FKA6MgI/yza6S19xhS6M5aZgZWzLUn
DTBSh3KIeq3rhBASUeVqrNPWNS9+5ZNAtPs+Ndyv/hU/za8V+DXmFlmgP4A5zF7hey1SEcEhdbv4
jOXNoxrQEZK236QXSwbFQAqzaSCIR7H+dCChaUJygSkfHystFDWRgs3+rin0SkuF3JQWUf7Ufya6
taodcYNRG0jHhHqMipTPC7e7hXcAqltuoBrDljLFraO6GFFA9bDuOQVnWhOPm8cs1O+AUg++arZs
AMcszVYeyjlnRkWM+EgnJefJGW+x0kgnDRZ/OcwGG9HT92sxWm9J3p/LQzd0s+JZf6OCr97gAcKX
cRwFh4yCrDcYs8vkz5KtoJN4xDu9O3Dru6fAFO5J3+NuLNR4ZvRQ0bpooQMJeOoT5r2KgQjYse0g
B1JwIzsp/s3MUDOyrb7AqTciwGckXqVBCyf40g4IeKGxpYQSqbeFrh8L3VHJfD0NgvDSP4Lf251e
GDP3UIjxZ5NwqrCbfDl4BRZSUDMi4oblcSsz8jODrgcpEuAN6rsAZzKkMHzq1cwxK3Yb0qNHpDz0
a98zTMqXI5CS2HnXRCvXJwN8Zk1wxz5UZ8XSMzch1txssi3vsRbOY1TK2BwqshePJuzFfAu5bEtK
LmfmBt92JGut3hhMtgydeaOTzmk46b+FaDoQYdWsGSfPuss5Wd1admXySzuZl+x3jCkpMsLTQLId
8sWdl3WpoGkmHXi+ImvqhPK6++EcvgPWTL8W2Si89AIlTgJCG91wz73YSBAxi0J57tG7rqoQmFDG
EpDaksLlWbFRTHy/z10mUeJNYBmzVeZw9ywBaqhbDt2J2fZeGpJxjeSkt2HbRHjIes5oc32zaZN/
BGi2zaRhNFyoqQmpj+wIhQLesBWk0QTDaD3FRjj/Vkpk9Vav+Jbzcmg5hAUduc7s3KGaAnI6xt72
w1Y4mOoMmcfqZR82ITau9xnigTNkbRmqOB4kNYXFTIb2cjpfSxD4e7iUbXPrvO8YEXj7mTrUhnLz
hrNUL22gJiX2h0KYterbxkki1bQ8cq2nbPLzk+CxgO7fGSLMCz9uIJyqSP2RXUQDJ4PJKdrR+cBZ
KizewzokK1yOMh2lYKhIVx6WbLBe1YhlPCgHEeB9T7hZ1v7q1PAr1d8/nnNbPonRYw2NlDzhbaGL
URlVHJqBpiGiiLDatkGvDjVUEVHRXLjB6rN9Yn1Ux9eGKcE4v9xYIMQ2gP+oKF16+ng2dvs8Khkk
4eFF/ceELTT5ze+FVdD8xrJ2nQDADIFPzf1avD4Z+k7uDhAZSgwqrKbwplBFUBFdS6dco+dP7OgM
p+MeXfU8OO3bZl7qedaIZ6qATRTktvxDCrccwr/hBT//lJMQjcJ+qT71IAYN4uWGU5l5EDFnw4+A
GX6yCZKc0CRg/lAK1nTNUT9pO8x1DRy8iM7u4dWvphfV8izD9Sc4UR+M6ic1SDqNp/J327MnSHk6
32s8bSzsdOi+oLVFxw6wZ34SFuEJO8BJsLuDH0PRddMZ3pRFiE297kIYJhNiRO56dAhhnJqmvdYd
7hCK1a6G4Z3KhORQsd2WICO90ozC1dnnQEd7UgK72RFXH70Jdd59veKR1PKunSswwm4nlPWXoiQp
TSenqmJRZPbytXeJPisaqgZNP1NbdgzLSBtY3HhGmsOZKe9oR6yrldLqXeeYUXa1mVaYXG0i333v
iM0RxfLy/QZxih1q1oeHZWn/tUF1KAG3U8FaZnHVvhQZXlEGgfbHFOcuBCvucz0ZFYNbXEhEczbz
8ggjnI6ig0j3IhqOC3KP3cmV97CPPGPjGQiOemJxPhHYVQm8kYJMSoiMrOo5uejIlAXSmDFMmMtc
m7FrMBzvtFh1+iHNf3cXhZuJUqhYVmZ6Rpy5JkS6uwM37X2Fy6K7AbnWvHjdvjATQWuuJifEcYId
Ul0VZYrBSnJncogqfgOFQ6DWs5zPXr9KA0pBGR/aXy9TUa/FWhMxyxi498v5g4B0UFUazJ/lfQfJ
11P9POY/ohKIAR29ayVUao0CkTxGTm6VkHCr/0/URZ8AT9Zn9GGQDh8sGRTkyzxHbT9JrIWx32KG
A9ZxBuse4zjoHG3JGfy/PPy6uJQR5EIemJ22Hpbk6h1pOEXBLNlepoffjp0esLU3ConSEaIktmcH
yrmLad9DzIglwWVBecUQZsxvgmpKZfkqjmVcjfasz9owk9DZ/S9dr8NoKOR90TDNZKbxioDdcy2a
ImK+M/83Euoc4wbdsJVZ2aK1X/MSsY9GiFd/gV3XiX6R7566375JzUDWkKA7TLwhC1Ug5MhIBHpo
Zx9WhtTRM9DxzmHrDX5eOPvCeJIpTrYYC5DQOlI3dwQrp9FVDazkFHwhwXsHdj64L4AyFRvlXa6w
oZs8b6kpZlWKzzwoyXuq56lggbzwTs1Uwbdpaa7hu1MAirVerUVVpmkGzXX5m9J2KJeWmRUJLTqS
ZXK9yEtoP2eFg2v6272lBhCl66PklhoMZOBANBjfACFmIrOSHDwNa4IaY5fokGF8ONGasY40y+UK
ZiufiIDagl5hRkVbxCASjkRKN9cDNGepAhCMPbRTuE4a7BOWTCBi1JpVMgml0AjMX6030RYi1Xps
i5dV2Me+kgbMjP1R49FiOG9LRYQpak0Hvgawtv08QDiv2MXRRDhymtJDD2qHLcw8dObP8wAVBsxy
+dMFXdoPqPJKiJpJ+Qc7pvHWb9Ype25BnWRj0/pJfVz4zIDLadWMxp7xz5EM0ybJxw/0XC0CpyS2
ksJLg00f+CzXgQzOQ+cGHWK8tCWOqxk+lJ2LWMNy5AskMKn7QFtRx2tIXRsdN37i8uddpS3LLS/y
J8Od9zkLmGD+kQskQiYSixw0LW8tA1pI/kNTP+jHzcTaPyYmn43wnXTuD65QH1GxIkqPiDo4Bt1Y
7acJlukDVEmZEJxON91pcLInOgr9ikziiWh6GxIx049YV84II2QMppIkSy2RRXqtxo4rjFnIFRUN
U3GsQJW9NYBMLak3p1YCIbbPIfOk14Ov8QCIKDNOas4j6AzJcda6dBeJerC+p4M0yYYOZnkLjNlx
2PBNsElgREPQztnO2Q3kdvs1IQhJ4nVH6vdcsyCRBDWCSh7/Xt1PsYGdMisvTy609YvSpQ/n4AMj
ZeP3mbESvBCk//CGo48ZcDkAFsLRnP63Jba8d1/nKBF+mVn/wcRpjz4uURx4XbgUtE7Sa+42xMIi
IBY7bzL8lQAV8PsTvhL/TnP8oq2j2rPrXDb6rv/40TWwufe1M3WwdB2VXqTqz4Zs9CAbZJnXKIIy
XNgjR7cW+x/XJs6HpLCVV2OJvJd69qNi6OuTk8X6vcVU0HDQgCksY8hE1dhFQbeRmnTxIlscuHA/
KUDGyJCFU85GWaK/ZHoZsow7cWJREni+P+WYWFyBszd2V5v23J7gUGRmlabJz0pFpNOgcCYwkRny
zAK7YNxL/Higpr9EwSACWc2uC3zxMnKLEDNeRoUWnV8wdBr9jX8NP9sXBhJz1YEEuFuuCceu9oe8
mbPF/tzYsA7hl7atl2/wcj/PvCST3vDEj9QyfJ1wzIiAPkcNA7NTBAL7Eeo+UMQtV7GKEy5BtxY3
w0RkZ3sgWFgKWQpvOvnDLS080r1iSxSzPSLXINwSKP5O1wj14TfXsp4OARKiRjyKHPxDLinxAAFb
dfrV5UeiK0NhGwxRKd8cuq6T8MuZ4hrzJkGXQUWeYyk9AEyZP57J71Ukax9V1UBQ6uba/7+wrv2p
7z6l/NPI3EDYiRzOgbTMjbl0lzu6cxinaK3tyYn9GxjRpqftARjR0WqftqCYEfJkYB63wwdTpcZf
moKLgRTUZCrWpqu7Ku725XvlwAqA7rFI4VSvgWus0CRWe9n1ndLI+FYYNxx8nG6KocngIhtMPiWY
M+a8ctwk8yg3x0WyAiELAt6KaeGv8wjiPwdTyTIwt+JdyNxWKa2ARAqVEV0f6iuIVjVitd6ejNx+
tk36VZ3cZeaj/K1Vf77qcbl2HOocebqFoxNxVwI7aPNmPVZfsLiccUN2AKaL6gbLI7zCXKXlVrjI
lde8sSMvCS+2wUg+g6z8GK5/TiV6zyw96TgxUtq1tb8vmtOStmhwSu4pzxj3BLvm3OlQs26l/4Dz
tqfrsomeOs9+iZZoHLA8mAUVVfgVGbaxqPCaR/yzQ4m1YqjwL47FMn7Pt1nqyHfmsFsyj4E2jOdS
3PLmApD/UzJUluOH9eRJOrkfyJoVg0dliJ8PZssQzsz1HCO177qDUejQpGmTJQeRu4KJBcoyZfpz
gyVPGFqb+JzlUnokJPLl0jH7gPF39SnJhIQM3ZWRbV9+h1eAOWx6SMoxvKq/uv1kjOWDb7SDPelI
eAOz4fm4jwCeL9ZQ/TWXo88Uo8xwbXzwoIvJFI0uF7VxWss4pcQ9FF6fy5qmI8+u0rWqzjZ140Un
SoK8GiIq6w/YGTGxsZ4sy6JCk2ZzgMtTWu1MtzO/9Ea8rzeZOZ4s1YWGL3YBqNwPfJ2elhn/3fRh
H4wC3EGOhzn3KXQ+zXd35qpU2RmmozTZOXDwPWWwJNrHNFqv+CaB9XHKGahlflqNt5/sgfiXSMBd
xW8zI+bNAuwgVPmwbnK3eOMdVL++5HgZ7RokW2s0NSaJr4m2Byp5SqmT05YURP4KAzKlOTC0gJ/V
oGNUEVpJ4TqXXBIo/a2+o2mzi/1nEFmX91fBsJYA5JZCrwMO64ju9w5FHJxibVo+UOe9695pCUak
0P4b+kmwTPwgRuE6BQlQpGhj3ECehPThI0jQ4q3x52KjhjeJ8z5UA2dN9Z0+st0W/jJjuLd7oRKB
yL8+SDejVH9a4mfCZBDxbC0aT2YYYv4VusLPisY3+z99QUPH4jChq8OLvh0OzCUcA4xuf2YdcKK0
nmUXhasX0R2UydTGdfaYIbU4iAY0YEm6wKEvPrNaRGGV5hmAjYozDSY1vAwvAh+crG6ya44tGCvJ
2eNsqVLfeHqvmD/r09uH8FsR8V2qQ21tSXvriwnwftL9gKA/jQCE4y1ng51Oyv1CUijGxvb7y9cJ
cVZkiLAJS0dZopI0Ak2VIb69YFYPpt3Uvp+hmOGYpDXVIE18Lv/X7nHzUofWxlEEKlc/0JxNRFSO
qi1j6aHSuMgczRZc2ZYnHe1EEJfHUQ58IV68pOwI9RZwLXRS1AFdDkU0014/9iM6UAIoMPUKqdOJ
qtFubw7OaiqZ6/aDgxIB8KfeO53zoiN8397hyuSsRXD3RHXe2mBVI2pyH0CSfVb0kts7Uio+/x+b
1TE5ShrlvEra323zRg66euu2f93XuuJT1E2jNnbixwGVFt/H67IvBdzk8YHFS5bK50eWuaWAtqFd
jCDLKFjr0qOpdtGTttOjBDJ/TAVTSfC442Dm605QJ35Lrt+rcbEi6hfX91G+Y2hB6syhEOndC1lP
Cq8b5S0raz5nxpOd1D0QEvt9YP928USabgPukN6gGk3wxIPQBrcYxTQLZvW3ADvHzfLOJtk4nvdM
irDk1dlAnLidTu7aV75Pr+jGEOMYIbS0YOFMfbY0SwMWqK86e08jvD+ApLqHtckkszYXpXCzpnwF
Ad+p1xLANTlUgE3S5XLSV7p8LKPHeT8/6Yan2YvEjQ15j9v1YJ7m59jBRZoc9S1JDXMyWkx/A1HJ
nV/dfdFPmtm6uxp/80kxQzdjPa8L/7AgJ06HdVBbtHzgBZpHEmW6aaZhpCjtBkoUi7usw3ort12i
BnDzJ8fiV99qPDHyl6EINKucwnWiVxrbZimLIz/C+4xFgRXHCN+RsLGnEOZZsSvvs+JfOqCeROQg
VvZEGbNL8z3G1QP1Oe61Am/GIWCwYabjQcxO5HeTVTqlcqAyp9If1IZ5R1L5TxXJFrJznqPKj9oA
rw9JUuhXGddAg8fcZq1DKiXSieN56EUUg/Itqo4oQcDEM5Iled+sh5hzCVS/WKULVqqU3a2WQfXy
1U8IcjAdQSwntQzT9yKJ46MS/ZVZghEHIqkk2ImOTyVhCr8uhVjC2RHBeNBL7rtjLVY5Z8Ob/KOg
7q69MpqCYb+ZVcN7OX0+CLAzcACSu/kHvgsB8gIqVoDfJogVV/m6ngDQRC6AYbJneFVgnoqqLg0J
rs9hMYQcI8OPEv1VHJNn0l1dRgxz9UZAcToHdrHmorroknuSVQgB+MHfZfHmu1zoKWzL/b0c1jpN
kg8ZQTI4NDK+AVMbpPW6RC5eDjox4oM4+G6PdcpagEoPXKIdnV5+EQCt0Eb0eT3AMuJ3b9O3IU1N
BIO1LNeVJWd3pnKYxA2Bx6zWz8A/ve95HJFiTMNUAD7/wZ1Cgh4pDyCLriSPCmc7bvtljzaL/JsX
467LX2TnMESAXMifXWhmNV1ijifGcqCCq8Bx+bn2y42zfKP/tfmekTD0FikFoR4Sueanhv60BmZP
twz6aZH0dWWItEiStsqsCNOt9Chj3WOCJYkOl8vxNTjXlCXwrwFrXLwKR8XjP3gN13uPb6k1FzKO
sNzphvP6GVSGUs4i7ibTifpibPweWCND/bxe0kYRG20+6qv5PGK1rfITrlRFk7X8+ggfewnnNaPk
7mynTYcQ1iMLcHm54Mf5kdaWPSeL7Wv2BoquPOAr4gVvKQ4oFf7tcPLFMrcAuFRMYC+vRH2Xb0qc
oHqK9uvwrtXxcCm9C8SApRLdDDPqBn8Xpy7azEAc0PPYOlHB7zhBeCWXLo7TYQKLqv2GwSGwE6VB
jWMwTx9F6XVOHbD2e9asX1mvKqRuokysb28l2dIT7bE0BdMbz0poYb6hR6Pw85Z+zburR0PFBZ6b
C53cnufCaF5lDumg1eDAoah3GSUsF8vzebu58ikZP7P8ybDpL4iCKEPJD+63IwDW3cPVvKo3quse
bCsveqJjpwRqyFOj49jpwbSiS4UtkFPMALWOSgzxagKjS/W8Z2f7TyhpItN2yv5JlWApRF7GH4a7
dhmU2ISJyvXGtJLr+f86QET3TgQ7tZeJEq8FF2cD5yQ63G9qVeoc/4vqHPlemJnAL8flnPQmts1l
uCROBHfzKyBJx2cA1RqfvZD1J0b7/fL/kJ/3ZMixZCO6SF75pJIoUgQCCppD4nGdWE10BPZF1LU4
dg05+iLcyc3MHVfPAwQoREPf80agyJRPgYY2YfZZ37OVCMaljIba+PBahMvz8GOdSjzl4MIg5d5R
Ktam+8/CFdQ/8oMC8m1s2SXe3P2ia7Nk572Hpt4YeoDFUITRxx174si39PEoaQMAHBcCh6tt7Gqm
mxYoMxExrOj8wz6ki0RXsLQTzZd4S/ke+SprFiI8/ooHKTCJPQrVCu+XoICfyFjcMLwWQ08WUaiU
qUsNTswcjfoP/Pnh88eI00ftG+F3AREectV2f+7FAvTgviPasPR7iXab2Ruw/Xh1W6FWiGnKN4PZ
ccI1u+kBzar4E7JYm7N9DxnS2yh4UJCa0ArzGjctlhI40g/H6j5aJTTizWcdg/lSJShbptZINjE5
r8IUrhxRKokOv65AhZjZ3qxSr7/GRg0XcWNdN1GNq7DHlrUIXM5Pq1q4A1pzoeVA5gI5zspGUTTi
+ssQvDRRsSNLeHn2Pl4AtbdUw138P3JNOUwM1rsnWSNfMBiXE5vBm7TBGXnEHmTsob75/hpweU6R
qhZSV0cGOrWdSVTIxVLTcL6RRWVc18pd+nNyvHOQ+41X+YUWQbvtzbT7zOHfqDhX5kzZkqQL4ETR
7h6YbGdMTPIk8GObV/BHEKhUKYrYZJB82VnFiVq3y7TCD/U3iWLkSCsNq6BZDuASDt9T9uz+0ls0
kl2KiQlcV6NzpSCOSiu3wd3495hj+4xD8AopXRbY6ABro9ZbSD2qx8Wkkeib4dTtFdXHVKhK464w
5hdWJgaRYdMcl5lqEma9xPPHKEQV4MR/xMZMfVM8ZH0f2dCei5umcW5HSbIWhjYAQls2KA8NqEEC
VBqTqsnVAmXxghp8VMfXNAyuxOoB1ohjQmixI25t7kaOy7Wc+0ke+nPbe8cqwoY4lUZi+7A590Wg
usp1Jzeym281oYpt2vBZo3dekEmn0OpOMIRRpE25AMZTKbG1u5iKkFwDr10nRHt17BrhgaafXx57
vgNrnKzKVkzXxx2R+pj/IHJ5+q6n82gZrGKrgf37MMoT1euDwPXyJbcH10sQeVwzDdsgBO7R+f5U
Vwah+wosaezGxgeQ6KoYBu4vmi/UAidipAi2TCkUOKmff/q1Ss/mVRr8uomNN4mF6u+jq8wz6Gi5
w6orp16UWlkzOQ08coj/3FX5r8TXEZaSOZoeVzm4sjrJe2JqVlAhRqTVdoO/Ahpve4Ok4N/Br7dV
Jqabgs6YdeIXtQ5w8+2BCfjtZs6Pe1nrsOdhyxeQzyayYCx+NZv/PoSlTNKS4ce/o9z4YhjRy8rV
bGKysmaNr9u1eooAflaX7JDXKTV1LJ+KsSxb7YiRAr1mzgIDLkEdWAAV2F8AOp7DgPsEY5Z5yR0+
1V7eoy1xhsrIIkDTZqHu2CU+EyzEF3Gpaz0VMGTX56fPnrne3rXqt2Xn4g/OLJa/r99+oojeCvLB
YxQ3ct6Yw7f2/J0SM5HdNLYLBh5zndJRk+zI86XCHylxU9iRO4GtbUnYJ2nCQRYbvFbMqzuJMup3
o1nDjUz3ZSOfCDzQyQlXC8vwJzqEsMueq6rFiQcsYsyQUAxseb/DToXMGt0jKubaFD2bBuAIaJFZ
nr5VeeQbvJAZquB4NCkRCFvR8XVxETZa/SWHcQsKckh8jM+Q1ur8cb4c9MqmFRSPhiypPGUXc7a9
xqJKijlvxsgYx2oeFD4vt06lG+DeYyc34KsASpV/Q2zJHMbnB5I9IWjZsxVZq0frONKpadUQ216j
OlY2qQ9ibdC85iYsDk5hql+SkWcBipwUiomhGhVGVijBxkJx7EdZ8uJmSIeDiUPkgio/3aUWNK81
qouQIL4LYu5WcVhJY/IiS3qoD4D9a9h44FVckiJJZzSefsbqP6ukzCvgwt+BheCf4FvkuhWbLzJm
hp8Vyqn3ySOYtl6IlSneBQoRzOm30uYPbYuJfevF1iGfybKADvunFKCd0nnO3g6gc3yj3COGKhhm
hsh+04iz5TVaJrn0DXtrBxSicKYbfhTs860gXWsqAQMxGbk3+qedxtdiD5xffE8cjBOxVEYtviIH
jt+dvJr+CJPS/lgM9sL9wNWqY46oavZzRzbqqIjvuIVIodyjevbD7MJ2mdkJcAKGcptJ4Gxl55V/
dehVyQG00m0iyui/uwWEzhak6L26iL1t/bmnEx5dUuNUibdcqjXem3wx2sv2SE7JB9WbLUI6ICt2
6kXSqi1FN+lGcDVafhr0SszALq+VMZYZKk6rPyRu8L2C0VOEzXc+fw/LGOtSxUZDoybpNAiNt+Hj
y+HL58SsMfrrRHR/VFOVhy8IQ2aBg2Wx0WJpk68u2Qw5Y97BMd+9vYhwF2U8oJJKY0f+nfjXXs4k
zbWfdAmZ/cm/6oSqVpX3IYmH0Qu37Bkca72D+RUNtXGuX4c3TY86KwjSZkbDfw+83n4kTINXgRI6
n3u4wp/t8dpI/X4TUWGWBAHwHgyojh/FJhCClsIr4qsRGkAxNjNED3LKWRThyoL8xY0Fj/ZhgJwD
CB/XbHaIk08neNT5rXZeyjfpQZvXMyC4BXtBG161iAKmgmb8g/K02bFHzf8MQRCu0OllG1Kl2GER
cAMmp8vq0tTgIIudcTgrpmA30A60rwIi5NCIt49c7yVZU+kM8q04K1Sg7Xn3V82ANd0n4d+3jZW4
uVqncIdK3MczAU2S4VO6rwGp3VFdSd8cteicNDBrWBvL+pK7khxHfhRqy4dlOu//zURIEknmBcUh
QFeJzC5b5JWttTAydwLdfYm6W7wfFzDQU5xx1inhY5VI7oO6xSovRGnuxx5SdRS9SOYZLd33KObc
SVZyN51ZMJ06snqgmL/WMmAKvr1kGPH3uw+ArBjNwY3WFhkMSDagsIslUVZ6eQ1myee98+5Jhb+n
Xe4H2gg6K0MkAM0UfsZHZnJLMFL2Hu5BSyR85QQEMv3iA6YBVfge4Uh2SapynpoBJAMiY6Ho4649
1CsYmfu5qjYX8fkNnf/4CWDF9wrFUNrgNo9DdSwGkCQoGsB4zellTEBuqawNJ4aSCz56Vwpf/3PR
hUl1YfmWIIheMoLUiQC5pJKo8kMgDUz/XH5fBP56Tx3YrD1tZM7FdtnvLbOl9sbsg7ywyI9Em2gP
7EGDfY7FYfFGyraAbYv4/FjRmBJy/n2KuTGRUTuONfmVbft1DECpNDHr/MB6bLqDBjrfoqM+YRwM
obf23wY21z+sxvRccKQTL4ByDZKQi5lPWrW09Mmw4eeBRjbyzKuk2a8Pyyuh3JAHiFPnoq+e4fwW
cy66VJsmrC/g0tETzLJLs2idUIXd0rx4StRedGVDj/bQTYdtsnJGirZSIVDi1ck7YN+g5RvVfIOz
OFisPRxOBFmTQRRWSakfcl22mVrcYLjFjOYkrbZ1Oolr2MoUfyXV31DTknlv9QOuInW2J+giBvXh
/9n926BE5voulO4NAfdhGPHIHvxXqacImlBcb58ln+vMeiAnZ3/FUP2DExbK2OhStdJXOJgMkCjc
TrXJ66Iwr3sVFM/1tgW/35EIWfRAzvnPtPNrCa7GBBV/9i38RbFTpc192mbcSrGPaJwd+TEOWf4S
r06RLLRXVaANo+nZOjzj1cJyrwgDe4yB2TWuPbrTPlI4n+Pb+OhPwDS6Z9yGycs0vOGND2t4HKxk
Wp6lhm2IUf8phaYd9NC3f7Ty8koN/W+wZDpq5qChexZg722iaXIF4Cfe5AARkwz9yb2C3/3fM+kJ
tYfLGKmDJjSdBod/7sTwU1esgx2STsvpWHgAmhjk4TsVU0tOPqL/uHjq6obK+LhkajSEMmAHqvM4
t5asgNDtoE8jXgAvNGFGQu2y1gWbbSvN+/rqVDbhmmAh3BLLjWLc7jikfYAQ3jMHSUcaG4mBGZQ1
JFQZuc3ia+yPh3wJbB4yOBLBwOmcu6cm/MVixa/i1ZkvdFmzF/+bdcvkms1gc4ijybmcK4N74ob9
hKShYWt6pT87+lGx5dlQgd8tKwhklc4vb+eRBElunGrJNS/HLW77clJkWm+qU2JGY44wdah4f4VP
XkaihhaFv+rxGdFMp8qHe1M14+dFjykOpgJRh6TXA2g4TOcpT0IC/seL673Wa2r9i8iEB03ztmO+
YKAH4rkd1Tki4RaPIcRbdpFvQ3CfzAW879gH4jhRCS/1AM9drJVok0wXjQH1Ilxc9DXtzcSzYI0R
pOJ3JEF3dXGBQ0RG7sNtB0+0hXAeEpxjQ3wI0WMll54YUlyABHh1yiFmAT4uWnIXAc3fndvD6s6C
PEF8TqUKi+f2M2Mt0MpAdig0bNnNeTze3JZx/YJhop2I+YEqBzmtDykpYjMyDTfURW+iPQOV7l0o
+9cm5z0kicIY6VxJtoTwFMB5PElmJkyiVeL5wtmoy82EcoQ56AEiMst0B+LL4v5+mADW5OxyJKYb
4doQiiB4+yfg8aiU7RrKykukYUOJO1BFSgBjLDTPjM9njhfTz5xa460Yxdc0ekSgndMnHkYwoLCJ
twsdbxPI1BeYUucTP3bInFUkbFltZu88TO/SQRR6a7huSS02jX+KUuHaRQHf6gZYZUdrXXL6MqKs
mgIFwME4T9ZuHKVBbhzNKqnDMnc2Q450t7ri0sVCz/cw+jxWf2oEoqSYfRzcMptNICfLTT44jrUr
bzh3RcKdTQ62eSWGRbYzrKEBDmtEbBMxmNvdnIDfHtUjKSBSO6ps9HEfXss829fuCHpkF5mk+Pah
NI3J9ox6DbYUiR96gXCZ5ZhoX/MBGIjsbP6rcv15tDivJO5p1kyZ7+veMtWoDitxAgCR9TPL2uWy
HDos4hmQyN4JS8xfiapJuIPCp7BU/Nw0audvZSNE5MUM7jjNmIt/IpUEW8Kgdn100ASkvUmJ/RIg
zlv3/0s5qcWuWw9qHu+E0t8dZiUe2Fba7HREstoTZmO/l5AK3fmH/aL7vmYHdb1A5vhJGehsVb30
miveEcu20YRyhjNRBs09CT8VSmRzdhAKxSaTclFwOlHjSWvBuNRqjzPLdJL/UAhOQBHP9Xg5vjC6
k8szGKIS/V0dpgapO0buPIUKPWlyZ0SN+ID2ccMANFXOGU1liGnh4SNlsDaDf3vrrE4JsUx6+qln
lgGwAmL4ktvekzWUx2ishQneVf3oS4855tKYxbpc4Z/QzNTjaNlknn20BPN6NqawEKl+WcIf4X04
Aa/g8zisffJbqrTbitJEC2TBjD1IOR7Yf0bl/d6hEYropWIZcx39qa/H8bAygP+WkUXmEo7bK5kd
rVG/J+XwFITvBbfbo/YL+5N6bjpxK4i4uHOcLJ8zbFXYEUFDxwuceB9+Bhgw2gINx74JjTcT31i1
GX8XxNyFmifXzppZxpguWZIp+sOFDSw40xWc1jNr7Ni5IbMx31rLiz4I7AZonrF2nWjRYWNf73TR
Iot8W+NVRc2O4QPSAoxB+NtReMlpOlxElLd/qkwpVla4ZhdFs9uOJ0GFdQKguXZ0mZZiPA7W48k0
eDVNQTsXgu+Jg7UyYmMCzPCoNnjuLkCPeNgLPtzsbBJml4FdMqWvlu40UPTSNbJNvBlfnoAHv0QW
NyjetEMEYaNSWrnOguQ95RwE7ogK4/8HcMOo7SfFQ/maS420PklA7dbw69NY5ilxF7LM/fDzAllK
ttvAwJoEDmrIMIG8BVrsRDiPobHncyJGtRWRjzKZ7Hjucgv/XYwq10DOIcmgQt8txzhLHIj0kKE2
hoADS5em0ELjdlRbBh6ye+QGj7Rc2l5/fXTbJXkekGIaOSwZKizubvw0hIVqTCHtOuocQfYnfYNA
AprPlZX7bcQLk7ezjjTPf0UosRS/3YyYgFAVHpemcU/rD4ziMuLWWOeALT29Bte6FF1vEl7arLpm
vAaXTXshe4Rq7sTsEpU7AeSp0GaN3mB0gombA1Azn5P9MFzH9ECVDTJdm6i29bRALRAqLSOpAZIi
7W74LpapHO7hZtjQGc65S0cyDKVXOfzsLKD6a3iJh1m97BlUGqpkJ1s/hn912RJBM7o4xYGmqRKP
JTN6D5fpb0xT/UHA4RdgKV3xx4RP1+hf8f8yT9Vt/mJ8golUG9IuXlD+O2NQEE3pcrnMtgOo8LK1
B080dcjmnVdY1XzIhBRHCyJlpJj87XddzxzsCPeeIYkar7nrUgf7WdJunDaJBlW8BUyEpuqSLF6L
ur+/6A5amZuDs6isW+/XojacDE9XDfLlKQQn5uJaDJwNtOyPTe9m1U/arph8ybhwEZicAjQXp3bm
X8UqX9m552t3/UzdD/nK0I/MglY1tlXWGC3sUs5+Hl/f2EKBFNgCvLtO3jjQrXbfFsEWGe3dgvXq
ppuAcrY9vb/ZVXLt2wdtpQpP79KUmPWVuelk9rC/P2uZ2ZOL1FKZ5euzwRBXo6Tbgtie7N95ikSf
O6YmnIoNc28rGfKVuB63NWq6nPTIk5gbb7sljpfEut3+JplPV+3fx/xHqVhhZClcv+HKTQOel9Vb
HEpdbEqK0aN5mxRqEagTdYWwxHmGZ045M5c+ymNQwtOVtVD2IDpeStExANTly58NkMu2jUXRRZ2e
eq2ROT5NVt5cV7uYealR/KT36oRe12mB/g45GK+PAI3A95R9Ed6OTgzxRs9dIOdHOpmW+yTjFpeS
FFe/RNckQcxiCEJ5fU2jmExxmLm0bdKL3rmv5i5lF80P4S0WkmHi6rmEti7dlYFw5iINlGYaYeRY
7kcTctOkQAxFqURKEnikjuFfifwjEWT5j2JLNqsfXBG5nkpkT2SyNr3AFXxuV6DFdx9yN1If2+J8
ykySnPzNGyqWZUMusywXVOyQ9cE4AugvMqxYls438v7eOu1L7u3+IKU3+ec62qylqNXpmGqZY6Ks
LYJyCAgfwNCYOJu9iicoZhrGIIsoqlG9OigxhY+LUqGL+2BiMffcZcJLC0o3Z0VHNAYFOnmTCMbg
XwOxeJXcgDPuPZwBLXF47IskVRs6dInAZWzaQlmRWifPlp+SICMc7dPzwcW5FOjf9zS9XsCgmai5
mDSCz2dCie4sU1YP5Vn50jXeCCMjfTihawW/5rHh80zafyvxMV7qwQ21KC7l0rZVbln6gt/FLncV
/gzNXfkxxuq9RtLqiEoy6n75tZgd71FF1hpYLXVGkHDD8dZGDu3r170IzeNrzwe/hg6Nu8Y9A853
yMJVdoa52d4NhE9gueuim5jvw3xhnbpPlG5fPRF4rabBvFgIGCHoxOtfX4O+nYSmL600JfzUykoi
hmsA9Xu8BGpadhlhD3EW+x99Xysh2tilo5KKM3Vbm+WQ6rNHBJTsvzdR+O7FerxcM+D68+l1Xqjk
6Mt2CGP/cwqEIAyJDizpZBxTiIxqsMpbOCNGBg+bCgtDDNRr7WTkT88nIOEoYDAsDD/KAIhYnfGa
7KbssDsXuDxxB9wvH+5N6aoaugGkNLDE+CCxIPz/ilaz+anCzqSRApwrqY8zttwSIKB4bpID0fgW
6Q2t/qFxeT/rNXpKtOdayxMfIEhopyq+jJ46XMLpxKRvQ5spMZ9f72G2Q93ctJuWpVBjujrcTsM6
ZQDiyuC60eydXfON0n/xmi+KwaTQVSGgk7YYh7Zx2U3WmypCjJskKYXgABA7fiGCQRtLd3FhhzJh
COlexicPakrnL3fdeX0Ctnw6p4mNQPJgzOlW23/3C/7Rw05+GeIJP65oDuG/UWNG9veSxO504YWA
S1HPR0t4NljjNOOA4LTf3YygHi/AjFao8P9DhUxoL4aGcdPg/n4kkNN9hVFNyyttczPzsaq6rXET
uk4Df5I9IhWEGntWQG0dstJXMsXdPq88+dZBre0Fkyi7JhczT4pTy9/Rns0YU3M7XR7lAxdLXCH1
qlaEr2CTcnejIKinPL1jBOi4trmt1LDZpzMGTxoP+jM7SNe10zB3abynzI2xivrsNQuO38StNrp9
HO5sByQd9IpeXIYnCPrU4oeeRhysmo9yQ8pCFrrwnt9Ixsf+19BnFGXux7/Mt3k+ZXNHPXdC1CYN
ZZzGDwWN4CIWryBB9pHELSvdHKLtKeZvOEMaCEOK3Dy6+VKjrVyDTnMzZ2qdEJtOtl4oHj1mX+oq
GqTifT0ssj2wniuxNSOiLDkN+aklpq01rR/SIsMW3L6zgYntV19o/IWygauZzJvkTzAEoSdJjqfK
yRVlDUDOPnrJL3aq+/BG60+gpbqdh08boJK6WRfj8wBXNHY5A4rXhae5WsPPY/IsN5PCWX0z1gwh
Zb7/3cHbbE3bYBQG2SXZyiUu3d14PWGiGhPtZ08qsYPX3i5mj4sVGcYHCwLN1MFklSWoVpEMtlqp
Xijoh24af/pA3mvo8MV5EWS5e5V0kXigHSbhLIEnBwYVyg5VfCpAUHX9aMAfAVOUiIo4w7ChBt/b
vPFLD6xQFEyqY7xfBDMipKbirDDS7gjNMWeOcdDbrOEiKhXHHjs0fXUhwxEyNj7EhpY+l4XbWAwV
vJPjUqkPT+rK9gn7fSIFw8hdjvFhRyFHaRfwEOukiAW01QEVhT1W6mBwe0CVwnJQT39ICQgG5qfS
hJXrInSVrlx639u5afCV7eRt86hOCYPxP8yjRhe5gOiCG11tMKWw4V1dKJaw+2iUrjESWz3E96A2
OwM+blW0EB0hkgf3V6/yjrxMs531EWzizPNMw382ahzUinkSo7k1OVmP7Q139T/Z7auJ9P6lCDxp
inuaiBWm1XiZSkvxbbjjf1ku9TfKAsEFpZ/2h3LmQbDTWSccaoNyvX1AJkEcWqg6k13rrZ82846r
fFkzYMDAabT3oTxMXRFM1qFU+j4Keqnghdw3RrbZ+LoqbhaTwRFh9Xfq6ZFEv5Iwq2j5+8j7HTF4
pidKTl9+Q/3thX8KJQjvEZzJA6gclG3i/C5RY7YQDiC/KGxSu60UlbpdUAAjkWqcYsXzBgK5X35K
xxTbA/IOLvQAjlnYcSi8PyS1s/w1ZduLqt/YPk01hSZ+iG9S1jcAzqlzeGU8Kf7T5BNuvyaMIutc
VmL6hxJtzMczIvfxGpMx1PuVdcOsybvaZxZ18gCHyZ2+OGlQZ97AT/EJwFwczQZI67fcQKCLvS1K
qGEynU9X1tj6pL/F44E/Ty0W7AT4rD6SQ+krB+63ulOQJAF2G/kWto8HJU94NUNUoTB2oyKeGsud
RvSLc2qnalO1MyzoooLvR6Aj6djH0RuzkiGzxdkBTHtYGNAjivbhl3zVA7XzSdEvI5Wb2gLqggEg
1481VDSGi32TV+gl+p21yFVMkmQWj0/CZSlwNGW0skO496RJw57sWG+ipYrHMnz50Nw/nuje6Wy7
1EoIk5BXGgf+S35Gj4uiRVoy8jYRPctng6hW+Fl6xU4nPzFr0Qe0Kvm5Nhfqw0x5gcUGndKub2KA
L/wNQvcU3q9mLCcW5kWU+8rZK8g7XZkl6KWgL3jy6ZErEh8TGGO9tPzIshZiTz9Wcj2yyDCKdIp/
HrdKfAGR8gULwx+x+VjE5ummddB2iMgjoHL+CdAuNUO5qm6amQZ2GCQcoNT+VZ5zBxP733F6gc0s
up/0tDGpeJdiQ3wC1f6emV7D/+lXDiJD1sl+W8FnM7kViopWK3sUR7s54pM4jjABsyVEiAfNOEm5
4Ob7+AHW1LJYYC9FMGB+gCrI5eMlu8lwJ+gMoVf9Ne2+sPoYJpumvQSGz3R8Umg9YkAQkQQjZSkb
4H4mf9RijuYOzgFIqsI5kn8rVbUS8m0d4tEk/UmS8V3J6rFOitPP9GBp0EQOqbybVhZLsdsUmTf/
DDtMCPCnCvSjJ/jwbkl2TMBb9TMOHwKQEmzbEnAV89Q99mIQaw1QKquthEUt5cGSeOyXMncTHEVR
Qgf+6pOjwwJ+poWtvL7rtJ67Rre8Bv5ZzhuaomMKIoOdgMgczKbknVFXI2TJx/pdwWI9LBnxXA2R
d5GpCdDtKiN6TJGM9v+iKNM6hGUXcUfV5HTpA1wFUTfji28EPT7tXtC2QyQdR3m/D8Lx5+eKCO+I
/bQa93SZvegxeNlevIl75FWiP8GciT6CwhBszBUU62EQwuh6e1H1qVbefeTcWScPghKGKBCgTXKA
cV2FM2gPMPbfPLdnXxWXVs7yY4mV+5GZhlL1gCNivMFZMusaDTL4857qVOH0TEakHOnJqlzRHynX
qDpyEVIweshckjsrae9Mke1JX51Ls2OSpfs+ki+pAcHiwmyfOQC675GgaGLQihdxXiOa1OM5U6ZS
aWOHRcTFDvsGMgzqNsEYMZg41ZAr6OUkfl+syrwzbVB1HrJXMiM/7WnQvnB7drdifT+Fov/6ztyo
zxwOD5+7sZP+ZHBE35LsZw0F71uNIGQfX+6WUPnttV0Hwki3GvfZtwoWWVKJ79EFmyEbDk7Z/X0i
L39L72wkpiu+AJgu7HrUxp/CxJ1CjT0AjQkN31YrUZTn8iZ+sTbSYmsGa8LDcsBh+ZvTwW/htUM2
XodKSozROUy7oMdf86QPz+pKdXxgWimZGOOAko4seafqnmVysY0GG8TT7ghXE7JnN642tsqoQ2SI
EzrTX9EuGYd70MMOT9rUYzjhqVs0wvk7acjulzXm/irjzrD0dVZ07tbsa9W83M/WwjQV5t/rpJha
Il6CArr1VZGXqLuV1/fzDSdbNsy4iZ1yBVcc2FEkutqG5YZnahZhSujV6K/RVdVNEC6Iv0EC272w
YsP4rMxnh0FHgVjL2fduJA/vVCwm4impZ3VygaYoGerI6C2HPfDQoRlVKet/aYcs2TPqKsOaPOpX
5r6rMNH1DpAb6N31r8FBYzS1/t15HZJD9M/FjmfDJutVlfdEh7UG//tkeZsyKtHTL/zV6Vnz/bex
7WyWoOt0AqNXMj/DVZ8OyYIV2YAthKOn4DDVoFHLu6jnEMaokp/bXLeo4ocEfL6ymgwm+vAr8mDg
X2ERFGNnYjSFJGGvyoQeQvN64jbH/tDYPULVkGS/ZNlIa+uxelbhQ8QTSZqWY/6cUXtcFwFkt+ap
cZo68OA7czzxSAyaNYN5EL6+dRomvrFklcJUe7INNAZ3rCzDhJVY3X0b42aS6q+xNpHgehQ/hwd8
XDg2Yf6OIMuC35eX6W9iq1PCD9XVjHwFfgOwL16sndDbDpGLq4h1t/17sID6SKAnpTpYUWyIqRP1
Jmdgp3Um0GGwF7I2fZqyFuivq1/pd5Zwe23Jwgbf672R9H57fd7ClG/AdAPUXlgl5mG1iOWA+C/3
XT4faGdrG30rj2gczr8CzkP4VZbiiM94CSTXPJ/+mjQ2ECaZazl/elgl/xRTsx8qppshPgyWLgNb
fYYvaiVIFCqup7NPGZXRwWtg/Gj5kahpxAescVvMVOBzjctJc3wzMf63zNmqFxXE13ScZ5l5HFdQ
L9cdihBR6kwWduieSwJsOUYcSH119TB8j+O47jABH+ELViumK3ki3X3tLRTwkCIeWYOK/812ZE3x
2Qs5B2lS/nU8qiJ0vHyV6Um8FXgt11J7Gqa+pM4UK1CY+1yNa753lj1FaMG5s2FMealnu7xS/HH9
lqJxhKNBijhX/LD5OpZpr4pzVIvGXAyM6Ts8vgG0pla+O707Ly/hqsEc1fzM5TqS45kJRN0oPr5K
ca/pDPPNpR9qxkXhjLQ/VwgM6ZfVa34WUXay2DS2nbULiJdPCWRdjG6ru0TPZ2kdhxyJ6+AsB19O
h9pOwT2CkNY9Qe5WeLx7pxEb4sIrZr5g+tgzhAwTdGsOONOmJCDNyfHUV/T9U6ixL9qWd6p8EEmj
KpyoLGLSFImHjF77XRWAa/DLuaeoUZriCrc5FSJtqbjuWfWaMU8LQurO/qAX8Ux0m+rcKqmQsIzt
Q3zko3V1DGVLt+6nUfuEYpyIAtkRQLPO5iOsWZUn+i3bn66jt0t8brbsJWe6LRqe91OMfZwzgm/Q
j61GugFPlsmYHhpEtNyaCbZWLxh+BdxXQ6KzYhMGXbVJjkZDGidXbJvPvqeT5MqvjhKNpOYWuLxG
yQ3/VZl2ro21Z9PJlWYkd8xiANhcSshD9g1i86ZBixmIBCPiHDgDQtZZZn9i6uqDJwx1AJ0SDicN
ePkemQ1ljYlZRg0/ruGvvUqE5KUq82H3tozcqQaoxMiUCTjOChR2mqzppoiKDfaxkhTOZWA9rsAp
JgSQSRwIolKFZOuF+diDWL7cbrkDOLT0Sr/h6NqJ3WRReSI6TAFocmI8MWqf26A6dqmu91VJ6JBd
3QddeD7jEWzqXUVXrfET1p2KTOdZxE8U60WrXZJGUmGylV00p9h6B4C7BpSRQzqfUlIOeSEH06qB
7uP/x6onCdmnAujUoC75e9xE+rpc9o2sE+sNBg5p44JU5IMpDst3Lejr8vi3bhsNPqNGxGI2j6Na
vdX4rHTntia4IwRKHNrjmyzKsgr7jX/w+u1gbyKsptWYgscsqtnE2JA80+0QQwanrlHxnXSk6Lty
44C+kg+xe7d84V6fHd6hjKpJ9P9ZJ2jtZZHi+wXEi1wgY8j4t+3Bg3LEwF0xdHI025Z4Yxt1z4zh
i9HR6rwLC2Za1/PikaihUeiJimh8slyIy1H9I1MOsQ6nx7b7swQsh/KlMHY10zIbQVeUQdquJscF
5T9V9iy4iT5RqPhzmNJ8ENtHA9inDcnMfktAm1u/CaKr97fiNVy0Mi6ZxyG3NIjY/02xjq9SJHKP
46mN+6A4NcJ/68DL/Xukf/5knbiRjbO2eGwArZJ4fm7tWyoE9BWXDcd8Zp848ND2exQ806adgaEb
iHweJTGR4rw1S3DiPOAhNxoR0SUcXKPxhQRsyBeM+k/Y/GsZemOQlPS0dF27xbXUqZT/y3/O4JTj
eYRxaPuyChhH5+SV68sQ7RFkCIwXucqnyb9zHOexI+j+6P2hnpD7+8ZxKjT2peLrhI/CngS0l8WA
9XkDFH3QapeSmEFptq79Gyj3DKGfydxGvB88x9fVwa3C4KdVUtln72vMiFFnodlEUboKAAQ6z5/e
OVxWewBl1aMAVFO4dq3L4nEYSDK4Ho8MGLLQt48UxGTvN62hMUov69XBQbk6juVY+TLTVyyCrQEX
S6W+HDzoWdUoPXT+B/J95NpX3ywQ7nb3tgSSh2BfuHvts61WyRuWzvmRJbLYRP6A/oPDVr42jDDE
VK9nXYKZVAcAHCl0NhHySt+3RWYkO4c77Sc/oMN5P3XA1T2Zoi3Dpgb+0wuOqv+JINJUMcH+IMMM
cTKHEt8Vpqfd6xpsSQCE2omO+seMpQOmXNBqnNxHkv2FVdgu46CgNsQWcLjOlvPEaQp/7MuoTY0p
kxsx8UOBNcGJp6u8z5I3MEhtSiNsM+e4dodz2/ct9MV+r8YiXwy38YO+EB6fo5Cc4T9jZQ9jqUTT
8Ot4WUN/WaEo8KmYBKKt6n7o12Xi6FApSgN/58/RqnhfsgFA1bEDOn08FF0XsE7IbBMXn9cE95wc
SmRvAc7dkwGpiw+ZHgkzVNwOxGMUx4FdtWHUYo3mUYI6KRe4m03x53EJHjRbMTAwhkbIUajirvie
FCVTyvsMNunGw/Hx6HoXUcWjqMXe/eo6NjzBI1ICE0wBqfo6ZwhEQJtEVqb0LuePGcY+GclOnva/
ccu1+eFiWSxv1b4m8IsA1IYYezTJGFiWU+vSXmEDvNKZ6GkNWjHNza1KfOSHeATUXTSZxsu0k/av
kRgohC/MWsX0gBDI8+qp8XcWQbakLu952cSNNeHbE+YSAm5HDSWoJegQDTWk32vuzDbQ+aydG/iG
1vZvs9hMWoIdL2McKOCWxPGNDRhIeInAKMPaSDGXUJANsDNk1TBmhOahhhRSE6uo+shuVKksnxt4
MtulLmdK58rtuZxRGjfhnxuwIi47GSEITjsmdhifDUxncZ3E+ArW4VdE9t2SBjulsYFY5ZiXqQ+s
1chJr1LDDVgFhwgaMt5ZACoDy2n+CyjLqQaIZ+iaDoxqj5yA1a98IQw6PDe2iRIWt/40rQmOUnc0
nadgptXprLtk8LKXsiwsA8yWjleefOuj7EqxKmj7JAFmVSzQLAZirLOIqaESU7qxCn+U8afN0dOX
NO415X+ZZCxMm/hVaBekOLL0PY51n63xGCG/Cnl61VUGHdmndGzW/D0IUOHcrJTJwosEBtc5kkTm
mBhI6h3FSatS2wIrOum6gghcol6+s4q/BOXfRGGmYFY5wkxB5EkrixsRdKVNq0rXsMZ5LTIDStro
raza3cPoOnpPnhJ4exbbNeJVQc85BeG5Ec61y/NMZnmC2jxiECOtyosKaseSPMai8ButixPhrP4p
9xCf82CKCqkZJ8u3BMZPI6NCWDMiMTEkBDtW9I6wGm1GSnYmnlxY/TmbrovyRzHIazt6gZndQRKf
eE7N9OcpQpMRQs5EzLp2ovdKIUxT0GLYqNKE52QCC93/9YFSa+OhwXXem2hAYzu+qRFqSn28t6nq
cwgSYCC7N5Ww7I3Xs0Ms/KlWb0tC3QmALQDQtWcykTfOjt3uKAqx0VG6E1D1hI4+KkkWHhhPbzdm
0P+ncIAw0dGrHFx3H5s7pfO5b3HN5qdILUQSFkPXcusGxlemKr3iSxjdNBkvIQFh6C9rqIrBxPyq
jhGho687RrfWq0rL36gwXDhJlaAVbQHI9Dwy1lgKm9c/jk2zzuZr2cusPqBbLSzZcx3DSBlOKu6Q
0z1s4u76MzN6y+/O5FPReKT6pYGBLhcODnDpGDr0RJQemnBl99F8eOhW0fMfnxXudhtCB8Zs7q+5
dJFELzF1h76lB92eWGv7wHpvbm4sQXEoXWqc+FaF3Fw/HeQbV23J6hkxMr+nXkCcIG4vYhqtPpJx
t15R/mdMD/N53PsjNC2qfHuFp1P52V9EE1iNi31y43vI7U/LngmOLlSAccGWj77O8ibe4e9UcUuB
hvg2Kfcx7P5yBDo2LefiPF0zEsU32goHWPzZ+FULs496ArBKyjo26ARQH1fFaajaRtHpPjuAHAoj
iidRyQ8p32ZKx1zzzkrq81PeMXgMNk4v8lXf7048bxvvABGJKFX7xajzTnLSHMNvDEli0SegcD0T
ymM5tLfxkZD8iY5xc1K9JhhTHdWPKQWbkBzNZZ/ELv75+43qZPBBIoPUsFU0XDlP2wdhaQ4izp9P
TWnJ7JRT55PkULfJUJOe7vphnzZ4jCw9o9xH7XIb44bEDy+wUSTXYd8ucokM+DQCYmrIWWlg1OLg
QWLRN69N9dvAnzIgHiZdyak+taEVs2CIHQIBG+6QSRHHh6eEEolqdENv3S5UKuk1SA61ZwSS6txs
ZZBH0korUsrBXo0jQ9+07Snk8e7EreFDd50FjEQGCwm5k21TApsm/aTj2qCGB4MKxU9v5dxZJ28E
D+GuA0HphDQPeCtBzOznUHbp6YJYqMCulAsIB8jL7cShTX2ykDwsraKp9hE1dsRSOmgeVRFNkVe3
r8k/XA6iS/AsmEQyTakVU7goTy9OU45q2GH4sJrcFef722AT39Y5pF6whaNLM8txSPNIzlGmdzEb
55tyEnFI6wdxSvvCTr6h0G0DWrFOw+qc/MS260kwpYrvf149Vr1WeUoavvsnlIU/2Em7g+MT7Wwh
2q/tbMbzvPQaxyVJilBxOyrmAs0WMZFwbhaQM36HRN6c3HgH1pZDaRES4PqUT2BJkpzwrwaQJZZB
2xx4G1rbE97T40YKgykCV3ruRCv3mZjxG8eh3FracWjT3CyfprJijvDO6cK4ugtitAjXUa+gMmFz
ybagrNDYUBucNbnssO10XCoj6eEOcx8UqIpNoGnolzXtwzAbVuam9NhKK1zsrMpS43LHnWU7HwN4
+yMp+7kUcMRXNp/KrCjdomsSsvgd7aPVSACBuZiF88/Nzlha4bQMNc5JRgWXoNtPEJG0ZEqxgplI
xOy6ZwsACuuShwWLTo3bbg05nKDLUzCmj8hrfYwHTVL6hAI/vHapuMo+gRZYxHnt5S+VmiRl5qO8
22z7NgPJrZXH5ODzoTPr0FRLktmz2G/grPrwD8ExUD7Z/O+qMvFeNqgNd9KlkNOKDMnRDZgyxFnL
9j+cLAOh/VuqULv4g+TxqRrypDMMLh71RPYPlcAhi/MGPxdCOhlrSrMfHwa6B2PCP5UNbtwYsXUb
3IiCraTdMGlj4+hV47dmvcR4j5eDTY/JsS9ZlIAAMUWwkTw83f1H+tj2sRlHdXygN85KfQ9cawL9
npZPm7aZ33hRjQDyVsSc+CRJ1mZJhF0Ul6auATH1MIiS3oXRD9+9Ue8p+O/Ebms4EiJmP0VMZWmS
TGAdONDDKIrNQYBhi3xVTeS7paaohzmo7IG03pjMu80ZdlffnahJ3TmLtfVzX37udG+md1sIrkht
ylT0+M87m8BWbf0yAcbYUxVB1N3Vkf75HeA7Zwqd7VrlplWCvfCkPUsTys2dUFQREThXt9sGA4I3
Uwbdth/zfDirwLT2OstGHy6wqYgF5987mxHTQRLUxHOCeiYtcQKRHsAKnKt0x/tRbbpEOmMEMs9P
VH4IPhX0wRvH+AiZ7XSPzN81vQFJuUnopZiX3TpYvOuA+3EsdRk7D46/tm9yURMm6YZfaDVDgSSZ
ZBmLB11nsP0QZyStWWJTyJbuzw69xsBQ20VcChVal2GHUwRaT7227a77uBUtTj17qhzPMsO1MzTV
Wfsh+m3VnH5hlNR83qCRlWE/JE1miaBAUw+ydvYFkxwQUDsj32uE76xjC4oCQbJCEXh3mmUpvXYn
Ic+q7sJMAjwpPVYKt/apA3Ouh+dO8U3ZyIirmTzDAbwPsiGxr4Oam8cFEQzIglFKUPtvzcJZUEHP
X4KvrQKErgGvcUa0QO02HQ4ABHFBQWvcWw1JqbroXcK3JoEljhcK+SVdbGFQGeQiRNipd1E98G7/
6lVgrhKfJrJvUIfY+0wzbwXsXqSRibQE/fTd+zWit8XztI/qMm7K3D3dQ0BlZgVTIO0T+TFCuxkW
XljFJCvQtxJ2xAEBA2tC2+vXNgy4mkksuNJ7uXD536LFG7dqfW24JKXOqIjVcDYc5vZWYmNDeU5Z
xB8Ze8wouuludg+TFYnR55EN/jngDGrVR3NRp828xz96ntvF2yq7it5DmSsc9xI06NEs1AKOIfH6
0+nu/f7C2oQq7uLWsr6e9vdAkFUEn9gMWv/pyYsbs8P/aLIYX1bMSYc/66Db27lgU9msceMavguo
nA5H8tXEKqZJHBgZkd0yqj4Ry+wHEepG/xdktAg63l/JQQU7czBZ4L/9tJ3jJuwXwBSLaPoMIQ8Y
dpClqb+S8/3iI5SV/O5pS9luP1kG8f08ndQlNTJJ5a+1p5MG/X+76lAWsVyM7S83dFICkYg9QZkk
AmpVo+zsQdb2PeZsJK70evMyRqgzu0Qxp4Lo2HcO/FnwUDhcykBscvtN0UnBGoK4fq0ChPxHfjsT
5YHWnfUMXgXThLlYNXQIGbyhk3uDivHtWoNuQiIGbwC4DlLOMmR1Wq3zvzZHYLpMQpNBdSrevYOc
4nepRM3FMQZZnAxBR3+wJwZDrb2XYmMwpXU+BGm5OmlFHZ6kW+YFN7Ca7TIz/tcJuLLHodmvCHS9
39wNCaladUHanyu6sqLKiyR1tCZWvA2ScdHUbSwwwIIhUCL2joVCY3QBO0JKw4LyZ4TpnOh99Eqs
l0zoqDnBlEyIGE27h5a8AZeMWxn1SpJjV9XofVbKV9BsjXG9FISZ8h/Qxa4Gd9Q0O0VLJskH7ZNZ
Zi3vzPxTFryKcYbQe9fRKzy3vygvS+z3CgXt7MEBs4JNq5mW+OuYmdDsvI+ggq2l8+tB7+6jTPLl
w7is9mB29I2uSaoEDcE3nPx2PxpCt5+9QHQZZE3nTgY9T1vfnNUAGTUjekglZ4//9D3Ks/RY0FvS
9ng8iXQhNRlCPEbcG2b86EzB95SZ9cg4mlwJ+EPJSmkad9hJx/tDFXW3x5ykTdIOmfQj113ymctz
2RvKUwhKRD8EsFiEjM8Tnr4LwHHj8r0JwT6+SzHfHr42iUz0XZ3N7OTtYCSnLTempINaLkT5/aGY
WU8oq0wdrPuyF3j9ZekEuSAagOAhTFWeGZoAPUOJNC7SeiZsSGw7AT4HimdPwzj7fK+5LYYuAV9S
K+nJ5xXigUqfg1/PMnSAGwVPS76Ve+QdrD2whmCfo3oLW40A9LDI9DzoygIoMBqSg5BZrU6wBQoJ
qswJKMcqT4KdnkwJVD8LcUq6AzsYNAY0BIDnI3zMgOwp0fMvNuNDcMLYG8Hg1Wc8eNGFKkoj+vu6
1R0tXlDJr5OzFAiRYsSM5ImkLaXU7IDSYsBsE1fi6fiStcGqjkUuI9zjU+MZB9hNTlMWq0Vba7US
JfknW6f7AjRwRI+gfe5xnbvHj79Fo+F2ttHEi6ZjddIjOfwZN5b+j0MK/F3Uk0UQTl7vO2vMpBm/
XW8KnK3RbmqLyEWFuiun21OYUKnVmhvfwW9pgd3eUOYlXobMCRn28YnlpCe+WfPWqGkcZt/h9Qcw
5pSC+DToppNPI8axe4V8pDL+iTWJZfzqpXET2UGusZSI7DPgjvSbqGJNBVOzuaWJ2L439eZg+PN3
FJUnjGj6HuqyYO6ppYhBBHBQYtSwPDrRi2Vd5plpgUsPjjQWjRmygJBAWCZsQ0O2LqCuALBF/HIk
lFSrGLkg2+ddCUZB+dFdU2eNWVA8Fhr360Qsr0zyOv99oRhVTkr9uxD/9OBxWtQdpMHu+ibr6qu2
jlwghn6p+14XRkNnEtWnsca+YSlYrhOe0HuOCZeIBb8RjIxtDeLv5Ri+VNJkdCtmtY3TYlZPreYx
ykpbtuZECt8Nhw1reBDhT2tRrjUxMBY691Q66jXeC7gAyz/u79r2mcosKgRjNE3UKyhMzIQkJ6PY
LTkhj6la+pkm6Hoe5MK3+EOd9Y59hUtnZufPyW1PQ7cnTUWEqKkpmujkZvzkizJAxFBHCM3udq3C
l/2UQV7X05CLBBG+2SuEre2b8ByyoJXZVBvMRHSn3PMfwBViSiTBtnTmHruF2t2X8/bI9sCdYhw3
ei9FgVSWfdBUDVTwacHl3rtkGYdxF7e3MEmNxo7ncUNT5+FqfXepPaIsUKUZvFrM9ZpHeC0HxOcE
45FYG6Qdu/jFO+tpsexruq2cTxjOV9wGyY/up6IYs9+PGYkxO1lz0znbqoJs4U+/K6UjiaH5Hoqs
ugBI/na81PZTLWZWYCwSHteVthbM7GF7Z/SStr+B6NNWXhnB/5ieTeanVrqoGyhvVi97o3Y1iKc5
PHd2RUMLyaaKweKpoBVq9r7mK2KbgjO9uzSAgy/hrUZahmOKzIhy7cWA/0TyJBQGMv4pQdMjD97g
+kzYo0fJ65lNe2m/SNR4hyFQD/fHe2qJHvU3PnwTxTI19e1NVhX0K0k3AEiQK+DodTLmKga4qDne
r70MOMLoQrG8/GEy7Vyr43woGFIOjwQuAgo7UQVnxKfyXz4SgrJCebkJ6t8TwYVY0X/brTzKV0XQ
GyP+3Kb9zP1E5R73wg25zGsS+IQNGfIMc1h8R76GWdxPPbJjLgMAUdbgXcKIHXHEDInb3SAI9CxC
kobClnSXqVkf439VP38RgbvGSrAkV5HoGRoIJILQhZBLLX7ARugFF/gUnBpenNXHA9h1CYp4IZNa
oK4GcM0O7BhLOPyUViC7imMLqQDmnBO/ySmmnqgjW9B+X54hKEYweT6mzBOykcwwOnCXLLhKWYKW
Sdtp0xWIML516Vetsbzz0JXRREbCS7Gi/yhmTSNXFv8yFJlrdbRisi048vzjKmLg1xW4fOyPMcCO
eWQg8KxS0iZcYk5FL+yv0GVtuWpzzCfeSdYOI+VdsSPf1blB/01cvNLBTGEKOyxGm5RoybWAhbNR
/43+/VC1E7IiMhDyRFgChGjuptXmJxXw6a7wtfpMX/L38OtVDEdKJmYmrhru2EauPPiyLDlMavz4
SOm+la60qcjXnGzEaG/F8Iwnrg4Ju+qBBIrdMBKN697d49N3oJAWZAAbr1ok0wHpI/N/lYgUfQlq
n1/NgrOcNUPT6x0ZZH6ZHVwTn0rtsiy0rhgktc5ijxOK5HKJ0m7XoldNaeSHrHXZsbLJWyssbtxh
HBx4vj0g+M9KXAlCwbIMQ5I4eiqHyo/SCPDqo91a4vb+Lgh0FJLPW3dmQcI/GbUKWN0J90FExYLe
0ThoZTbWBXBZqM70o2Or4JsCGrnuW3FkBkCrxENg6jDIl1M/lnvItabfu05wbddDS8dztFz6DpRf
rXz0YXQf276/S78ac2flOUDjwzgeLGCFd6C1Tze2tERlv2j6RSUMjWmpdLFiDikcOp5vFSpqsW3a
bGvfpKHf5BwKYtVHS80u1OBdDdAxD0w6TG6ZKk/BmgGWreJNA4+noI3qa4pXq1+k55PUSUBFGCI4
+oFQ03PbsFldyeHbrWaMbEAfAy9/Cyu+6yBsp0kmfOvsEQYDMr9IIffd62VWZgkDdsA5O4MJjUfu
Z/n80gapl0lvcOQwBnddy8kGZUrcGYWNmxVV3JgN3P0zzfR6OnQoat8o7294FCEatpXKr7CJx4zV
MLLmOjJXZ+3GG3J677LwF3AYMGJx+7eldbkUIjoSPi2pwpYfimDYzDGfAcrcuLjHwVJnRUpLdT9B
XqAJQGIZsoPsnErpsmhu8I6jgJ6xNh8jgwWI2GtuOCFFVmJJxIximAHvltu5F8zBoYOZ7+8h9aEr
pikAnR0I21Wo/UOl6IddZFESq4sU6hcgQEXjcXnYQpsIkqEhDcP7U1Bv0z67A1COJIEUOdLzPFTf
PsXkFfzMHkhmx8cVndwhndQKbLqB61SFXUMPDQJoa+LVEnVDwldnWMTBoGrFreukCpIKrDeZb5Ny
Vz0Ik9QHERQ+h4Xur6m6HRFR413awghvduck1CDPjO61wy/IQwERPi0lFxNmvXmH4sDcyjIQMuyM
UlgvCGzQ7BoGovsZoong9q7UjcuQP/YkTCsj46LTdb4T9r0jY1YF06az6ZM3XIJg9J8dwNVBa9zH
CTgJYEZF/Ayo3K7Cp/7QDAymRCNBQU9UkdcvsIbjtAyUG1BfH6yQ9zHdYVx3CS2/MaOaQaipN6fs
tlzvNF8WRQ7mcdZ0u35KyEv1jAMQuJcQeXRxKCygOgcDYK7zDRo+Ogs/IxXmcAx7yb5IioFB3Diw
l5dIhME/SdjncK0heI624yMQmVMmFJApC3r3i0R8EpRRatISMKM3ZuzzKn9e5tIQI7D/uxVTLz23
QdtSU9cFlyucxshv9xSuqh1xwDa3VCkxfxx+791hpWA+ZBWKmYXgc9FSUqaEg9/D+KfCT8dwNEwn
brSKsbQC+meDN6gya2k+4fCZKegBfisKPdBZhcTZQcLClchfQrbS8lLG71cY8nq4BtP6Hm9Kvvkq
bSWAarnnd8KpJgJflxqTj55ZejjLmnqmlQYS8rKAkIJ/U+d41HugmJAjWxgaGV0yeP/UJmgXbSf/
rfi+9y9wUSkCw6FRrJJknXkYrdynVjrphlCd8TXs7lROn71joW5/x3N4MzhiNtpG9HMtE9GrMGDj
Ly0IO/KyZRybUVQ++duD4VEn8MRBZ+omXJPO6poAcZDDEsyfhbM1znCeXmpgXtF0cFtW1Hi92zPa
Xbek6FryYMjP2WZZge2szj3tGSWmPpVyQtk2u8q1boNkzRLwyYKz51cywqqhnSf/aCblt9KjTVV8
croRfr9IHFGe5kpUvRPQofBMm7/cC6vNZbUMov5kBIsDm8Wcc7oRtjBNymypJhv7e72F/cEkY/co
5JC8090XcStNcN7yaz9+aYD1iMxJ6DGNAds/bMrC08gXFpZaqoSv4v6PQoo/oBXcoYesVpQ1GFyg
JhlL26CSbI2WgnhTh1uZ6FA5RrFWre7F2hZTmoNymZk6dw1KwxYPD78j6ip1HTzGbhCwtmIjTzXv
7d0gmpkqelYnc/sb1uAWpQ1fGegcu7SP4ygUK6gArTN5YZoyeFLBl40vy86suUkb+SC/KSXBOMeL
WHrQnq2S5Z7pM35DVbI91lVI2okXSoUBV7C7XCyEJIaWj0nkuyHb4mIipkHUtjB3IPpsiLdOBADp
Q4/XJ8BO69MwoNfdDksSsAJHIzLfP3BJvmDstFw6aEp4lqBp5VcuthUu/1XhMoek5qEihX34FO/H
moOrqoulyhJbNoz4VqjWDeiBa07H9Bnz/k0+VXsjnef5et26jyh9SVkqgd39PbLwOsDEx4M3ZrBp
y8hBp74bMzILKNbJ38onXGLVX1yKgXCoInfov3UmRI4cCv5tKVzOaYgmEMDXw5+egUeCx8ZBwxMZ
4rYQoCgpKH11HnIYR7w1lDHxBVucXWVSKzut1HK+q9BWgKb7OM6PDB3OWDS3BxX3jw+crTGf82uY
knwBA+iAZbviwRrTidyK2PwBWf0gw5NKGfOA8HbOR9I0fNQ/9w40GPfnay3eHMu9tTZkyZbZGOx5
KWytMT9w5u3GSFyZv/nSO8JNJoBoUoHLs7MqrD/vJOxrrwdYD9gl8RRGUDn9xTT9to1wBt3riTzM
5dbuAbPoag6NICnceztV2fxW9IHTtG7qGMIGLguDwwEAdWmw68pbEIBX5b4t0jPn5OtXxw/RrU5I
ZAS81b8ybf2rKmI7cJY46wHVJdAXWkT2w3hZxsYMKE/hTQJahMxdD8nolKtsSUDUhLYD62m+uTab
4/ld3js7CfWL5/B39C1ohHjH1C5i+2iq6Kk9jdfyVKvCtHN7kUbgmQx8Nzkxz7bhAzhSCI5J//Sl
QDL3mF3Y91wzMK4ukvROhdlVBla+7cDL+5hQ1SQWebkn5BddNmrFrBzUPmk7P4YmcVezvKN1iY0O
xvVbAMAu2tlngGho90FGuMugCHfV4nMcOxcbmRtbgx4PEUoObo7hqOAx7HS2t+WQ3D1HWa10nzZb
I+vdMu1hqPjocL12B/BL6J+/FmvSpz5K9GOuX6Iq3NBda633Qzmw33S10nUKJ/7PdEPWon41vAwV
v3H0qglImDg9CY2KmiYpzrmSanNo7SDp+vb8BJWqNgIBzxWSedZPJBjtgtyTj6nIor8KeAnJwfPX
us+TOTHni2RINvIzLWB0Hx1TQmjWWw7+Iyx9ihMaodjSy8YGk2y7KgM94/iz8tHnVPn+hUjgAYHt
An73L08MIo9qeNUfURVpVGcpvclzwsAeZQ6gM8L9IIbzqTTGedA7pUauGvZ9dch7IVYBKOW1/oB/
kRUS1/kOrkt68dbpD8Xmi0qdsldnGbNEj00vYmFXBEllUsqXBfvu1LpsDNZl/OE5qDx1Sc3D9v5V
m+Z5mo/XjQ7QSBvJF9ECrbC2UM9t6o2/gH3/+wLOHUrQ5fWpERY/lony2WrGuYDxPz41Weze2mho
yeFmUN3TkHWrg0Ybjvh4bMakVMdIyKaXT3YjZUxDtTI79ewxXYQlsvakEqjQ/n3CVDX6D8AExnxl
7yFChPb23v0oHIHQu+r/Ek1sKa7yTnUobE0HQXP916Chh+cYdQMeaB3cems6CmSyeyrQ5PL0Rv2y
dMarcO+ZHS5++cNNNokP8uIushi10/tniSKu4rMvApdJE3LWNuaDFF1OpLvFeiBGA5/VixN/tj8e
UQNPlPDFnCB2CE+rcHwJ9HEuJbbzS/YXSheOLeRlUMPCexyFj6pMJJU3KUvZjofk8pqh7nGJntCg
SfHw1NyfoKG1fW883LACvncGIgnatXr+3dMso7go4/tcl2ATKVXCGxHHVbtNDEbb8SHITiLatDjR
UyknCkkjCM3U8fLwZS0bhx69inR7WdrE3P/QPx8vHFXv9NZhQaiWdFvs4KHncE8+2NJcsc4HFiD1
W/8NoxUEtDAhkAxSfbvv/gzUFo8dQmfkLkxgs9q7hQKUUUKONyv9v+M5nsmsTdWStVs5mY4XAVOs
3ZQMBCCyO0+2lgUjzASo/cu68vyLPceLOqLrrIYMTHstrucaBd6gywQcdK6anzJmlMCrMe766D0W
EdDrh+U647jCSmoGi7wyK8er8YFHxCOfbxSjXwMrZa4f1/XlclMeBGXDnzA6XSaZKwzk7UXotOC/
ma3HVE3Y/UY5mTSQ5QVc0nKVp94LvE4qRnCERgNWEm8EcqGCGeHIQtdgovzK5yjoEV2vzMnEjSra
FVXi7+WFTc9iOsOkvIQiBHOr1NUT6ccaPFleGUDG5FAhbEGZ4lBWGdB0N6LlnrT3qqzLmHzNBGl4
+t0uL4VOZ+DSG4NRtuMvTirA757t1diFic7hVI2tQ6a3mZ61lPuTa3GRaPHEWNozVOaV5o1wjDgH
qARg6BPzJ66FKg2hlz/MUzULaUP9LFKrs6OT0Yf/vOm00hoG2/R3PyDfRCCbmRPuIHSW5pFR9FCs
Ew+sym/mDGR+m4Tw6d6SFWittIr8E4yde3BVpxAXZ9JAfO68l34I+CSCh9DXcRJmPWxMZdnRX+9P
1eVfwKYJYLXZpGMHEcRdBOYYHYtYKxA3TcIuzvrDKBW5d0CD0hGDRX7anMTpmQng6bdk8O+IMu9N
C9FbFOqX8KwOFO1hELz15vB1EN0E5SByOwruIg6156FlY1/a7UqJM01qlBQCsYVehPowosj8jxJ/
08Rye9465j/la+tZE0A+Ug+QfOkqWofUukp60hPT7zbwcpij1rnsXcWGJ6dRIlPZQ7Wumptpc+vx
0mln2DgKm8/NI3j6ykXVrMV5OSg5UDIMZiBeWHn786kg1Dz55NmdgCtDkIUkApsgCHkjtMLWpP1T
Q3mAFBUDqUftBEnL4BHD8mFxtnsvbOZeHfoUJk+oD+wjykT6r1O6v6HGc6wBnJjyK0/5+hHi1Kdn
Z6qLnCqusAH0GESvcS8DSXt7JTumRbu0UGaEIFi9kZYMG+5x7MGnpxCoJbTyL8wHi4IOk7nOUOcE
FjOiYn/7y8pEMdwBvjABt0a/fnVpyqzMyHjt9LNviwcqX3iR5XRyw/qS+lnQTx/zXRQ79qtfb66t
I7oASCec47JSVV4L9jcem+2B0vf6nD4Wkq2sNdGY3lB+DTztI0kKSokEZbeRh5dHeKv0A1oNQBE/
dkworvVbgPxvqgZr4sm/y3GdqFYkjOxDssY2LSNr3DqW5SVTPjS+XgjLBlSxGKhDiZW+nUqEo3pJ
zxSE9bIgMKVG/cmPhb5xN2uD5UKI1DDnSa4N+LdxOxNWS3UdRCuoh/2zyi4pHnu9OzJcsvXgG4tp
4Y7k1DvQOMqUj/1Y57kgxWhbTignBgTROuotxHAVyzeDc7QDaCEcuPPhfZ0yP8d+uWe70K9+TdpI
uiCjUm7zDnPuf/q9YS3+BRljHlhl/wCM7TQJ8Xcn4eSbiX/Z66/+dUonQD+IQbpIBYytb77ZCO+r
f78A2qzx3wfDGARJWeJqGq4z9IIH9XnFjsRX8EKU42N+GC7KI3Wss5crsARNk3ZlFJFV5740fyTC
XoIs3sa2ej0TU9drOtHA/oAXhHCDTORkRsrCZMBZebY8ssCa92y3ZtpOsVCSeKX9iTb+UloBIH7L
0yHj4aKK13bFca5CFfoBrAQRQQbPtEuS1LLsgnUs33X+RP/NAQx9UD2JRBV60pHTLZQyODwGD3zp
CzZPBiDVPLazmgO/aM8otosCM50VnA25Zqt+6e+hJFiz+qy0l9aDKgfcUSN++CRVYhrcvGlY2RGc
eEr88l+kjJqfouwZwfkovwPMrszSV3uBRsLA7vdHRcxNpXLUkQNTbyfFMt3hKFoRFAbFLukgZuD6
uKJdCf19ZzaJUuGiEENHp3rjNupXtI2H1MA/KfY4CeaR65irdaXZoDrnZR1cq256Z1o/WGiV5t99
Ma128YssoVzs800xgN6KozQ+KrsxcwS5GWfTdO1T79tjQrffGdKFP8Vf/f8bDXFXHFZTk8QrzqYM
9nAcdWpq+LOtqKvPXnz81fat+MJ34g8vQF7tGn1uLaW082Kl4ZziaDo4XrqEBjSkKyoMWkjKYDKg
ros3aV+enQbvfE46LEDgMaBkGm9MDsh5U3Git06oVXIb/K87iDHE6a8s9AO4eV0L57P66NTi2XRu
ZbPynTvnqv1OGL4MJ06Fukqbww/espgz71W7d0JWoSXrkDedi1hF0MFHK15ccJv2SjP58ds+tEXt
bMCVFpLcInjD1kRutg6N9L9EpQon1ghwCpbjKcSlxrdxDCkA+eObdQUjVDWH5fzaCoyQZutWmckH
gnPmmJWau54EWgkOig4NOz+He8moP6nsz9fgWwoJYJyAEPnU3I3ID3u03gCRdQzDjTS0yGgzAKBz
m6qf2v/f7Yh8vakSdmiayHgNBHiw3j1cqdcbkgC6uCFzKuKf4EtOqhbIngtmfauhkudEvo4AxG6f
OovpNYUquDG8/iGo6FiyL89l1zOFaaZePpXwVSy1IF3OMiHqMqO57rBs5PNSsx8DKyhWGi3/yXeb
QV5wsojXY5drADLx/WzWN8dExBh4AGuLEuq9AOBu5juBzwd/np2wmRFhIV2BPXv5dImPDvFKzvw9
yYsMZp7CB5IuT3rOHs3KGV8EDirRz46UFnFaxEdKrmoUjxl4MEfXcK3xPb7vJi/ODC5OKi7ZEZ3T
Kj8jLpCva2PSVla73iSVN0+KiKmVdeMC8oju2zS+qBgUMsroEMsM/Xvcrg/+HVOFTgASH6x+kdis
iFMO/OcLrEG65IM21mSIBzrqVuEjphD3RiNLxAJ2k8N6o5t5zk2iku/mF6gOOo+pivS3gxqgSn0U
XsonaOEOJ4Abt3ksxmyZYvEHTnD+C/Nl6cuatoFjwkhxLYsu7GajSCp2d/8MTWiQc+qDHG4wBhW0
b0960TB9sILRkdCGUpMLfv0UsLLQcJzXl4e2h+Q0nDDVzrqxEHEt6mURXQBAv5ivLCcMEA/WJ4lx
BWTjNWEnuf3g0RzrWtDHytt9saljas7A47UD5o1oi57a+Eb59DQwbbO56gLRAe5Ik0lkhW/1PQjx
+xI9WtcihLX8zzXsuikgQ6f993DexllKytZnpVV2O+CBXr2pNpub6kb9FW+SzHjLfKOX06HH6RLf
bZFoAWobOCo2Pe2F0IefEKyF27h/sM5BRbvTd3hbnS89Czhv5EgkvE4r0OVAo9Yl3WZlBg7aWumn
UgogWLcSkjXUbB58qdv/jrpLEV2OWPfYGguMEg/iPnWLHr6OncsrSI4O6bUNAdG8WZ53CL6sC+P1
UTtNlLMf+TExjBIrgffLzsER03yWoxG+4h2Xhayhz37m1BQeTCwRAS6doaI2zFNarUf3p9ywjOp7
hOsJZ816Rwz5s62hkWpyzFwhmof10ELzQ1WubPlzsIBKCEFBZ+ZzOCHzRl0RBNS9XzaDI/Kfd9oL
G5fXISMxPGd3nrIzTEuLxEsDxKOOcsIWMdimX54rIMbHY+AjuyCV+HcHcbAAk7mVW1ruQORRFVQU
Prrslw/thry8elyxVLQNBHb00IEaWODtPLwlV8ErY9XZ8R9MPvkcMLTR9GKqrww9THcWkgmlF4PL
SgA5ggAJ2PLezYFEhoTJapOZQxu0P4N03XTb5JFr3sURv9BlWogo2T0fTIfuioJ136i/x8a4nYqG
Kk92LCldM/m/w+aWgh+W/s1nc48uxmR0WDeuCmYpt4rcwGuGhKQdkORMRNm8lljTK6W3ogGGP8Zn
AdXAFcWIDLQGrhHsst83HB7MPQsQhYxPlrdX6LiCpNSCtSYRMk36JnC2imL8m8dh7Lu5aOsg6E88
LpR4/JYWLWYuqigqECjf8njO6rlCcsYo6wzegkc0KThq1ot4OtuTYYm+VEtYWWoVNj7ZLuDHbL6k
e6fsZ4ohQlEwFEAHMqQCVC3669lHMGwIO4ceepuxJcCxu80UYkoyTDCrBNm4VikvhnKKZOZkq3tN
chiRzUKT4kr43zUAIYvlXEsSg9L5a5ZtxtTP5C2r10HDBxBN/Snd2v6GNXxNHQqkRcHxDeZI1+KK
vaNLb2g6vtK76185t5IomV1UUX69Il5a0/5jj7fel+sBdx8ERghiLa+bl/PwTh9p9pntLSdlbVUl
1jbJVuxGqixuwmMJz1+5+3Bwj952aeqSbqevKl/W7amy9hn0U/3ViyV4PtXPJTNTQvvQr4tJo1o3
3q44ZodyEZwwCLuHa4JltEimBvsMp0pS0nbiirYtXHt9CmeHZWaGFWwQY+h/r9vvwCCmtUwKqnu2
3WJrX/1ttgEw8DFcLA0kKpEPsMUbz2E2ZsxvP724W6Lhv+VwLX0Xkb+W1ZWLyM3CHGB1caIEQGVc
kX87fH6kN6oQQQjzkjCeIhSYAvpLTalAb4MQR38/iOJkfXsi/CLvy62NFQtV5PstmW9mlrgnHZev
2QoVEIH8rRENUBJNYy6z4EAzA2An7M+/tFAq6WXYH+XhieLF9oFeRRGsnZsfpsmcJLdgXx57YwT2
XAVFw9lp7/IRDJaw06eFju2Xpa9HB/L0rtqvH9huIN1N2CUdCJryHsDpvAiUJCedBNVcmGD71ObP
JkSPPDgf6REJDBTA9X/c8QbBGpZnIWY56DxFDRgukoz0kYFd7MTOJBQNMCS1L/ryxNPVszJy7gAW
GJVHMFx8krNdFy1/QhCbzGvYqIcQItDNRGJzin8a7ZjcntFownOK8W2U7T9Y/ahjcDOLEHIAQFvz
XwXVIDcsTSQV96o0NaKDOy9jkVvoDwJMgv3fYPbQFLagW/qGApCueHcwWd6bEmoJ4JiSJqP0p2Lz
UbbM5INLddBOzDqgdA5ecLIXxl/Xk1If7LoTvUFn34/2Lrf7GOChUoe0GZmE87wu05+veOyGUJfS
L9CAe+KLz1nDhCba9diX6bcYHaaC4LPeBkvAXYEGPsF9bE5y9RKpVOCiX+U/oVrpT2Y0edDrggSQ
lRLza1CTicXNry03mhuY+yqfpcpW7+B33STEYkxFm+dURlxvHg5660s6m2lhHZhJu3nAI/8FyBUT
kOWFrn63cZKkZgSgncSSFlF2H9JAoPwAbr6LCoib7rGqICEsuUtIuWbHUvHCGhUaBVAsJALYGHq0
rJu4+SMRl2QBPfiedLr0QMyk+/SEJJeLOeqOMcG8WsMf824WSrvzMel34tBxaVHq9rPFDBpdLfkp
+Q+8v4zdHkAZG0EPoGmvlSnyUR8F1lsrx2IWNZVRyd6emPWgFr4tCxmBPRFAC9AMmW8DMK5cDfuS
Qgc/b0gCGs9zS9Eqkq4eB6jOna5BvE3NBDBCrkQhzy8bNrV1RcheuRx+kWFk4Sj9smnauy9LzIaa
ImaLW+ZdKXldVw4IA/7k/JGXHdj3fh8yLaRB0RzWLAmt86VkbX9mrC1sbmYForKWH0UFkAGQ1l7A
rCO1dqWC0k/bc29TOUJ51R1rDdNMLu6lKYCVGziyu/NKdqlLMu1xLxiNQqHlOXEBeanGWG/z6TYf
XehObhxeAiFSlj4+BHzN6kmth7ByAeHOn1v+rZwQ+hWG6ewvH2at7yDed3m9htCozxycZ7zoLrS1
RzaKUMfs/tHC8LkdSVN/8YdYGHrYfk+UlicMT87ducjNDaClIym/lcBWHaE+XDht0Us8uQLaR6cw
XCZWiVwqSY+1LoBr+CKcSCKBpdTrx+68rYKOqSESQdCob2qkRQddbihpvmRO38RPk8enwhzOwvXT
kxFkS0B+0fTckC6LEKQoJddNCmLAsdH7fdbpIE7ydqKnZpwe83kW/VMJj9B5dFwLm/kDNnu+SccN
TVt3kLWA0kA6r4IVHmeHbyxgKszeKzzFAV0eX4MHX3i/KLJNuQUuiUAhVs3Hkdb8fjG2YNMy2gqG
ix9qkM4SBiNvUGIYT6A8bMwS21AnDx+ciEi3sgbFYbHf6Z30J/ab/DGooMnKwtEUK98CGlbroY+3
m13u2tovZFwss1pLQgloV9dEG8+mZWAsCaUOHULpjsZm1KlZmL73PVnjznEoE/LwY+MPLwz7brfq
MTNrwVquNQQDUVoDAJCUhQZIZybYcZzh0Hl9BsmLq5jTAhc1qEEwfOWf55lHQb+CVb7xvmHtn+mh
wZCm1xqRqq3gcyhVLegMN3VJw3UbngvYfnVpKy82tkR6nurA7WAc/3OD77adtpNz4VH12jbPZmc0
/EPl/StXwTyNSAX9TDsvU7HFcvT4R4SH5Au9x5yomJMcQW8JxeEGl4wkkvFC62aJSXUlx02nC5pM
9uaTsdvLfHQfoo56CtqTr/37rnv3GFsimkIvj9Myd04nV23U6sQfSnp1R3iTPcoZlXl66HPXX1sr
3pae5eRhDgrSJOYJ/GVW64DRGdkeFQY5re6AUchA7D5LT9RAkxnGNOQpOCGF9pHkdd0unbgw2+fb
Z/rRw5LSDtLNLCL2AsnQvFQ8u9wurzOITod/xNWclKVy+pFQduO3JuumXwt3jNYQzWe23Wj6fgBv
bLVLbxo/toNkXbYLTqr8jIr9fVs1X6KtCSRe2EcGX0vqO3Wc53MLPlOx5mBRR74iK3ZvN/3tXyr+
XyHxsN7RcpDIFtLsJcQuhnlCWS680cs5qq04qVCdt1Um0YMcsJIgrA7N2JDgt6n8YH3ToAQd1baV
n4psu4gR5wlnX+HsaFukrFQEQv5iMuno/1BFOhNPzq7WpECZX3KwZkWQfdPt7QXkrY/wsZCl7ljo
ReViP2pMIz++q9tUUEdt03n9u1MPZiW6aopKNGLrLJpbJI/JbDxqVDns1RNMsFQCeM9Ic7Ao8P3Y
/ssq/XkU0+YAoI4ZqX/gY1hbDsWRuQ3ArWrQuW5u2CaZqavFzpq/jXe8CvjkoLvhGTSfFdlevvv6
1tGM97K3nd+XRhYKppWdA+hinHNbPI8F2Gs0k0ATxPI8oS7s9i0g/h6M5b2VDIdWNDVGM/tz+J4f
28z2Ht64JbhCbZcSSKfUgKxMjoThg6ZLb1zyQfekDvS1pTo7ANOEXvk1Py8qaMcv/Y0zzxEe+Lb1
AEWs+lI6T3CYPZooMHiEKkJHn7q9tQYvZcj5RUTBexGxesn0f91Plk2X3AowNSmnbuB5PjwRkZHV
l0wfgExxP6HOB1ummqxXRu5tYS9qrCZHOTS0VtznmjsAhmdiHmYMp+NOg4yRCS+D3o5mx2JSDXgo
5h4+IqeR2R8AZZ2i4o9uDbTxdugsBU+CwnK01QWBLM4dIXmpsvIexKYyXrhrWv2A+XJ4hFlYLPh3
cJQgqz0aPLVEIE+Cm86JmU6H7JX/I/628j+4msuZL8P1HnarbwTbvEhY1PhGWSgZwnQ0ifuYW848
gH3mEyBe8rwFDqtqCUp5oL5M5WTyf6tdew4B0nOCHT5hTT7vZi456l8T//vOzmvS4xpHdaT0v5cS
2E5wMXGyyOQHRNLxsOjwtpODry9gSKoPNiH4qjmMYmNQu8v2camQi2l/jUh316jCgI2ux7hppYAs
vOEpwVBmJShfQ/RBQQqCLCXiZoWtploO+jT+OplYlNOUO5kfMyqtS033yns5SY+Sve/IZYTOpFqw
YLm9M0rTPuLXIGFH/vyLT/eKG3iZ+Prqwq3ZSKOKFuNyGikobC1UWyWWyQVcjxUHHmJbujsbH5Qh
zyZKEShdjTiXApY6N8lx6r1W0whqSqrPZvEbM2Sr2R0vdsj2ZgRM9PrQAZ/vOX3XrUGJOre3LREK
2UCIZdgHLX11zIANm0eo9YSiZPs3DIBOqo7naZa2RIEacdz3qzvQNTgWo06Z63wY56bNTMjqLoUT
nGyGUkj1E5IR2TWzZvy3TlDel1BtJDG3aeAbQ9RVf5aZ1IbWpJovxEkSTL//ut7EwQQoCPasBD7P
TZhAhtg/3Dld61Ozn7N/4VJqebrpnW9RnUbmfi7xWGkOHHqcFTSgRltahVu2EB5zS8R4WCtab56r
FpWyUoETO3dcLKFsSzMJqwKzTTMdM6LOEMPkOeyJZR/e5eImoUkzqDaOppVgsJhWtK878PvlEBJW
EJ/q1k8O2FlfD0g46PCBs4Jkkn610G2ouGT+D5rUQwcjli4BmrhaGf/mheT7KqbqIU00rHhTMoH1
M32NBckbwO3V8tQ92jO670KvR527TAJ0cDfgnMtqug5zTIZ1wOV0svNd5LJExoU9Mk6cZBPl4Jz7
AVOBDshhtCA9ZH0Oe4M1zurt2Qjck/JfqxZ9ZEWP51eBgNs1E+SC1HY5QDo8fr6w8dqYzoSuoMxa
EF5+rI5dBlOGwEJ+cIG/ULMI0ENbm0wJLxBIXB84+7iSsUwvg4cDvLndCEAinHsb4rD/n9GrAaVh
fUvIVJa0np5mSKOY0Jel/CfMgAuL9T0x6gIyWI4buZhZdz3Agar65n4VvrBBKzxJbvmOcA8JyTPG
Id7d71JrhZCxPnalpglv1ZUlqyK+P831pjJ25a7fL4Kx9lj6ORKhZqvP2yB3iBwr5W2tsB9bMMzY
oIgkByjG53iyzU+wB8ad+uRbTg33ao2zWktTD/5HCmEy/fuG3bKnK1VIVLe99UgTz46wX6mTL51b
vgC5ZXF1MyGyQtKMAcwJ5wiGym79WuyA4cTWpDjaH64EWxtnfPMpCxI+vM4u8E5aaXLs3AHeCxI3
ESS0Fd0PU+lAQ3EYMoC5rzpPDDBsByMxfquWkdClnoQBovQocGIm8mYtGePoLK8VpQM4B8+p3Y/H
ubYWgv6/uoBUxk2Ht2TCUKiBS7Ir4G0f5UXiunvJOwGLHqh0uJ93oO0dLVtw1PUZADU5xXmV5QO/
HiY2zfdiFoy+QX0gNv8Td9EoHkesl3aiFVAeXEibmwSWxTtjP1CoiZzSsFT+TFrZ41o92i2bH6DS
JsAZD/oiwvzG/GGASqOuoKStysQ4MiuiacOiJ1JioK0eC6LLVC3pfAcq0Q70uffPjLGLKQMMAOUB
c36wctn5g1VsMd+is7cuvrm3bpKR0/PYvuxk1gruXUZ4Ufr5NtNrJxm3ZcHjiPF0fE6WKI31kywI
2kVh2jSc0kMJaXVOHI7NC/53BjCiGPAHqZvxg+ljXw7h3Ozwya5hrSLnERxL4+o3E3Puf+P24v8G
/wgtHiLiwjbQQs43q1JTYsDlGoApE40UiUfboFNO5cq7FNK/lx/6Ega53pgEntfC4r+2GOLbpaqC
DkOuxsQ31UH30Jdj8dQrvH3ZecJZRVjIwL8NtgPRsQxLBFDpc4UsgtKQlvLtT/IMx+anaAj2VG0b
jCiWDmLxMvxz+1dx/pkPMI1N/mi41elLEe+48KVl1NepLWz5KlGW9m5qzfA2Irl5/On0XeRi3iqk
Z3+HMcRzcNPfA6pZpFJTcXZT/+alzzmzP9CPJCOSYJUl5g0QkVOJqrMraav/3JArehyOMZ92ddp6
1K3INkuxCIQdGXSUDY8qXJe2ZBSbezEqxoG6sIB3mzs2gPkKKriStki5gBJPGor1lOXitbrSQuRk
q36gfa7ubRKenB1WfsalhzBgjrEbQ6gfMez/MuortpOt6md4TGoJKlugXQU0DtoQz8XhxHeToAjd
k8jX787Pyh/xp4Yd0ky3ctGADSCqkOHCznYlgdg2U+ezgJIiW/UqUJGGLew6J1pPxXi0HBuKID5J
6qOhYnnrr+zqt3m+HC7eeFBTAR0EQhxmnbl3c4UJf5DlYFE0ldATnDHV6krec5rU3W1iSd2MAXrc
/CinHhewq+4Hnyg6G3m3GterVXr+Ow7gQtyweaVtIC1W6jusRP/PhV+MYyDb97HJY4AsuntCYaqg
2fpCOFpDII18K5WoUuWHwqikHh+GexBMmOA+UB0kQ3LLZjapKj9DcJe7reXA28Oc0/JD7QDJ0K6g
ljahF7uYkYeGcjJcGjqSpmo7AMko6GJP+hB1E2l2tT/B0QHP051KEJfCkG20awl3sYiAg6aoiTu3
yE7jScuYJ5or4Jk8+anm56GFjPqP4wQT7NHcPjaYw7JtmJmkLBRP6Zpdcr/YtMty1QLI2bgO7G2U
Sl4yw/BX3NxH7EyC/myoANDSgpXTvuZ1Ss/tHwC7Rqi40MKRyHlcvq/sjMVqobNtQSZ2BHoz1sGc
6CjtoQIyVj/1MBiSL5XPSvC2yZ+K/e7diNu2N3KieKDx5ouuDHLW9ayskhDP97mb+OA/UjbLtpcC
ZK941lcLg6ieWQ1/1RumbrJJwL56mFoP2jlMC/QoCz9khYLzW04HUGU4CEOrf8q5hEiTOHh+mjZn
Uflkk9HuzzmZR/giG7wXqjwXp91Dsn1ts7nqwpGR2YcNSsfQBtt6EedJ1/iQBWKUyjQJMXgVN4SL
VL9TFsahKqiERXi8mEaqbHhlbxbzoTQlUhP7IVXti7ly5oxz+m3qrkO9CZt3DHRk0ykfaa5zH/n8
T345vYCjI8jeIy3wzKMYUNFOUSHkQkkwiFbld27a8qhbsDgjLKiZs9pJd0s9SrVtch5M4bZ10RDn
6ITUShxrxwdx2zugoaX0GNDDX26UsBKUPWg6fwvUEFflJbolRdcyvFXPv+tu7ZUfe5WKavG4VFi9
2K9WGo9StXap84MqfDj4bLkQOuahWbKx1ximslLGQCbZ3k0Xt4cJY1oke8UAcn/TyhwiQGxKeyuB
bGbQlkAcfsy4XunD5xnOzzD89VNUFS9j+K7mdPI/PyMR5AIOy2zCkMvY4TJtz2/D1BGaUPXd9aMn
TQZws+jGFf76aw1uHbkjD2PhnWTZAGYsQADr4UQ7bVOiA9cNI5Yd3VZh1O02Kn76BdmATr8A8vnd
9bia5zF6OQbsxPPOfGFUIaAZ/3U1PJtcMKyPt4A6oqqEoPRCzV8f6Ow44TnkAjfwXv4kml+kpbJY
5ZE6DRYsKgNOcbeY8EFepZjK+rbNaolsM87aaiY57C1mzgk1cP92emwzaHHZRUA5/OLcqV4t4cLZ
1GqBviq/JpL2U3MdwFX7ZTHmsi9qb7oAqXd6N/0hQUYuEzF4Z75Uuv5Zm4cMk7X9uMN8Ot87irzy
pLHpF0XWtRI2rGD4ECeNQVWrmWLdjaWAjOHsfgIe69cJB1L+VD74jUXSBFdxiJpsPERYpnGNKyaq
qhdT0r5L4II2SZDrAPDKCjDJiFSd6BjXHxtzKP5vmEsJBnTJhzYeO0F67RF7GGL1gWdb2ZLI+JLE
3r8+Xqo+fa7qItaLJCwBG8QJKHW+N5Z9dErDukAWKdY1nodN2DeFJldFmCe+0hdE+Qh0u6Y+6zUv
xllxprbrN6CM/A/zdU1imSGEEqrVfLj0KT2NEUy7wVAYqW4z5qTZyUd5j1PC6g7ml+R1lBeTPi+g
Io4Y/9OgwzAtU77POqtlebKM5Z6haGL4hrYzLwoV0XOZVKOHWertGfpXK+Wei//qGnO5NjNoMe/I
PsyPEPuoH4bQSU1GLlXMHgEoST24udPtEgDmcIqYF8eBMuFdIF7SA1QhYpeXuPktb34qYJ+gcMmn
i1W52AssRCxmVuaSQkO7Cx0e2jAjqUJPan/eE+hyeLsOeR8pBxOApYJwEfptX4dwx4TEbXXJACW6
gYDQGBg6Mic5pHI2s10rl/apfWPpna3INN2AU6ofc/Igcu+5T75HLcqk5upxmj2XBxWaS2wUbzk8
J68+g04bks4Q7QALfr423QHiBwHirYE1yC6svrQhZTVohUN7V9C0XNANsYH9C9Ce04giTNFrxTli
82zfF2acNDZxeZBySZ3fEyyeL4EmqUTH8aTP3C/+RwJIT9SqqQ3UVaqOH4wU31Y820mGJOM/qbLx
OigCX9bOnL02stIU0HAualXCNQ25XIyWruF+P+7MZZ3ZBmhheMhdS4n57u5C69484jKLmfa0fFPm
ZCtV8CIXOS7L98YeVC4qwCxrxRFi1WL/6S4aOrT7nqiXAOJL2gs0xs0yY2IJPLhIE6TAVOz4c2SX
xLQTcc5L5JpfnosXVgivsS6NQxGSQfPobyC1yW3BAL1dsnEl+1bv347sqpG5/VoScItZt0ttNmyX
2YrQk36BA3BKr0sQtj9vzGbS9/aLKLhtXcVXikZ6z/0/dYyx6HpdTszhZAFsfrphW+StV3dG4+1N
PT4zAHzX6RGrWDYMX249e2UYIgmh0KSf2ay8Y7dCULD2yrwZvy4qwqHIsKwnRxTZ3UEQeKIsqwd4
75NrSq31Exmi3zq7l2lrvmnYKznt6GCO9LaLDLiTVgV8+utGaXCd3M1dIYYSbdp/A40kX2DOS4lc
lzGJKgTPB7eZtCF+qqxA9ozw2kUchXUBzcw4llR6oxOuFK+vFxIXaHjX+Ghu9v1GDTauNfp40iCg
8W37Rv6VeoyJylNZmyKFpWq6uk0mupMz1CZhgLTkz1mL/RgPGcCPV9Zu3qeQPbqTka8yDUuyiI9Q
6N2QwKliHxZB4tb1HN5UCGAv7KoDYJhsICWuGuJj4IleHfQS+cyplmgHUwj3M7PJbD2OhJ/891DZ
zs5Crb78p4Rp51RlLR6G/hanAH2/RbGUe5q/Y1wY4os3/j4Yx3bL/Ps++hZRXxv28ZFL3k3cDu/w
7Xw1lfuLDuVPzQU8zTWuAzvtxQsxUR4e6QdFZKsHSiD2JOyoWD/eX/883xVfLuBTy+Y2DWer7Iq7
Oh1PzfMlCCZAj7jiOEfu8iekvp4r64+WxRzbArvEkjtowg6TSW1SfwDdabXiAgVrwRXe8HOtZosm
HFrgJDq1+2r/QlXTsI9RPA/6vGK/nAe86tIVhR/hjyDEvKXD5X9wVae+rBfi1FT+oWjHW8qvPcNQ
6y0aELExrRWZ9hbzmEeMq/v199l31KZ2tmVDKTYm5n2/zTVGeV56OECxNwzapFHQhYtyXLOSjkdR
sFUmp0nULSoBcFMeKYie3Q547AWYHSmeZme6j+15cSkIxwoSPta5/qkxJXoI7FfWKLh0buo1nI6b
PtHwixL+a6JABT1QKwj82nnKhgRZQ6Cd6/UkQpLRSWN00aijt6qwZhXnBqe8kB2byrO9MJe69aDI
Ji+EgRnzGFQraKbv4zBNGto+32QOp8tmlTuh4RTN1JMWgJUuagghmYjpHux/TdhbtI6PVaFXZGqd
tQzZGx/3SA/AVzkBb30liQGT5xVPluXs53tq4IOm4jyo3IvO1RHvMYKm2TdDSwAMYeQ02IlGT7Hn
tozhU7hnf9iaBHXszP612mO5ByWvqo1eI2UUnP+4pgwjL5GIho2706twPagUrawvGwrvQV8o+rTE
KKSpvdsxf3MGy3Dm1g0TBqCEQHT4NFnXvMF6PmnZw5sM89qPWzEApEl3kCpd/nFcGx3RaHTXaDCK
qTQPy0Crkmy/iSdFMv1U2ouldOZWiaSyixr91PWSoHQc9porNLawCIAbU/gKZMaFhSd3kv4wptFe
/iPiE54g5zpBipXKJXCAO2IcDBjCe9yZbY9M4lJNdOIIWyPiOcSqPU+f6w91+qgL0puIfnouatm5
jsUGiGtbC8hu0ijNnNEz0EoyYCFxtGwovh0do0hGSeu9/7e3ytz8xxX0wCDZu9y/wNyMVMFEk8YH
zLWr3Nw4vIskc82e1eI3t4NamQcBgmrDTc9oMsUAjbgBXeD3KnYd/pv8FiaEDbfsZujFm/vlV+4y
FPNi73zID5hV5XhMeZXZ3Hf4Jl+6M8vlgjzABxVr0OB/aAyJ9wboYQLUy/44xinYnAyz0tIH0f8R
ctzxHLA0gnWkP9GrM112seIJY6QvLIxpdRGtAeCIIHTji8xLa21H9qZ8nNKufmxuA5feCJ0jQYNi
LGwW+a6kkoY/JQrKwfPXbYT7zjUwjvEr9i719T2jk3eEeaXcFMeJ5+XsYIqXcN0pVfElOlMYBSFO
rcqYNTbS9W3McXIH1/GvXIVMYtOdshHkqsWjSrKmpMyUglldmCLpejhIEv8H4g6w3EHgtK6r3oqo
60zUKM5IahIZKU8sAnzpQuvO9tCwQhnMvfTx6A3cEtn2COWhnJtPr2I/Kh4N6242aNnPiiS9f35H
BTvGNg552clmgXWKpLylNgGThrX9ebzTdO0Cg388/NaEKpgl/UIkID+jPdHnyz91QNlnL7w1Zcdo
o2++eQm6IOfEcOFq9XNOzKsmN1e6NnuVQAJg0HZ6OePZPTcU1gUK8ZqKXlci3PkVVeaE+6EGv34x
Lzaey9/wWfiW3YK7AGenQcuPpWmNQaQ1/aiIheNuoTG0UYJMkRZ6xvfCNJBtctaRzxtGsPZbQ3tF
N1Zr91OqXRoTvWGbT6VFOx+6tRoKE7hXa3ZZ5Kl3Nh4+TCt5yu+7pGqc8HiGsA1cW0ssIjZexTcQ
e07HgSfrJTMkZP2ROXnz59o6F5RTYfuPgwOSeoQAOaTT2Y878b5e82EdPYQPpd7JnG5dfBQhAeiE
Lj9nvB3JWWvGlAiODJy0la8wMJWPBeD2/2bxpnB3yaNFUMbLjVjvy05M1nbdy8z6qr02jupAZqyl
fOUJoWJKKX2V2xaswM0fJqv0svU8JjfldkNncfGpFqOC1Owr8IaqTPUrR39KhU6X4Z/8Qadh0aCf
2UrZsgqeX8XmOB2FF/DaflZMH/ELmS1uAVgst9b6nusJjhUkpgN0jGymuKp3b6+LhzVib2bDnKx9
7AQFZUTT1tcKYY9TUT5xV9UeOOMm02fhHMlin9qT6RwxXKsvBqyBGJu2M2da/4BiygWAKbNVzMdg
RQJzAPYO0+gwb2++DyBHXoZZto5bQejAlU8NQ7f+bnjEB5zkFNcRv74hBWvA/hYpr6VEyacXijZL
Sd07nOh+lcnI3zJ985vLeNXDYPy6bcKYvLztTBESF51fM3ooffWmasj1aUATU50OR30lSLTpDOJX
NcccVf33M/CzZzq7u2tGfR0yotfxC2ZrLsF5MKI92CQnsts5N2DsJoWrmFtmJVGZtTXqdeetDyae
Zvv8R+Pg1g/R5TAPk8IW8FdbLOlr+20rUgOjfOzU9TH7c7BcYBo8n9Q8mEdScc9emAYP7Q4JYqZm
n70mzOsTsImktNbR47DbfJhlG2By/GYhcYF2Pnrl+BHUB6D8g6qxn7bqFjG+e35bM3B2yYc7NJdv
lfSpdHd6+YKP+KhlWqBsogu8PJFYJH0J9ig9qMNAqCPiR9Aj2IFuI2lSWfOlXnS0S4OoAFxnOW9J
vWW6PC4rMffi1W8TS/bT3e43pouqZvdUdYr9PFuNWuJurZVX4we6aq1H2inwHko/eEH84DUJu9Q2
m63pzHNZaEbxSDGbtNwgw37hoRnCgo7Dv2HcITBo+xNl7vFZdDeSuPQ6Zk22GWclevkpHT068gxO
621L0g8UdG7DTOJrdmM77zQTXBMn4PLFx8uLewpuQQhhDvt23WwI6fyxpcG+WbsJ/OSNuF4sl+I4
w6pe6UjwXBNSE5SPHaXZgVKpiGhUVL/FttKp2DIG0mwcwoi+MYWK0T58WQhFrEIiWg0rR9wW8CfB
IYAPSGfcupeGsv7I4/kCOhx+6z6qaR87mlVoUsAdIdYQpdl+douq0yzhUtuXjYMVOQ6tYeYrJR4M
5NoB58e1UW6pC3t7p3ozjzA/KNvB7CCe+gNSKQLntihV1DWwmina6uMm5iZ8FRs2Qac9kYr9nwaR
vaQ4d++T04nWIQvaZ1szhKsRGZpBOSi6hQBvRNoDNilo/seEJJoTlydzpmpDodwfJqhSa/FtZL2y
AaxdvKtKt+PheeL+DQj1aK5J3ewGkL6zDmGChoT6mRjm14AVzEBLu0UN46KDXWVwtnLn93bL28rN
RbnB/+bOrhHQQn6y8MgVo5Ch+iMQUpdDAhMJtQsOcdT0HKFny9XvU2nB/h6NxQNXMB1v+NXUkio2
qF13iwewYOC9zld6viB9EHYRsjc0iaxIUZrqrMNHrO+F8fdsj0hKY5FHKbBuft8HmUiCfn1/UlTW
Sm1i/D6UjdVzg6+/D02r85g96VeVwNY6EHuxhe5LLKff8w/Nb61dOKaIypFrEJC/w782+1lwVszn
EW+ds2EHBTYyOnWlfsDK5ltylKmq7mEhg1ET9Xg0wnV21TZD0tEse6injLKSxPx/0/AYYwRTL2OC
ZPeOz+UvtpdohGqeuwJDWRkIRNXNVzEoBw7HDVm3/HGeoHJMJM0CiuIPK1fx/2h4zJlEQCDCQ0zX
S9uIQ70mwWbDTdM2UjZ1mDyc0JSCqhH4qVrrGI0of+WrrH1jzC0ZIQOz9ZxCTKXySQcJN8uYGtkP
ZfpzTt5j6f9n0t9foIz72tFsyq+oIt0ZhIh2GdoE1tY6jWDsv54UtJPqiSYEPqpUhEGHQF0sqOWc
0UaEnzOU+hiViSznrNRass1b4/hyEtxTyurhOzXhUU4uJgNx/MHnSaGna1BEg2xrMwYWZ0T3PpXO
918QB8KWkcS6vrChUoTZUZximZgaY8bQODOB8yHGEx+cfQ7lz3NsifRrLvsNabFppIpktK2sHh9B
KDdDfZSW+Y0u6DWNjWXZSi6xGfxNgzyTxSe50OM4hcZNCZKmm4CN70mT67maD0iD/YLc9MTbFusR
vIXe78+cCLcQLhoHu7/F1KzUIAeV5IbOLGhsX9lHMXxOEm8ebhsrEE3muiHC4sKKR/9N2Ytsxq9R
cI3W1oU86zbOfDVaUC28gpeUhtaTIFP2S0FZJ6itpVPNDFR/UChItAGhlivrJ/P7qyGQisrbQ5Xy
vmAnJUtYUULG6Tl25bEtZOXl2lqDUaooxHurq8Lwiw7i6lUSCale5Sok8K2cn2Z+UnV8og0mhj8K
0F5paTHaJsvad3GxswgaXKrpOEc9chm1LxnC7UbThIk8AO+XURWJicQmyVt3RrZPH5/99ZIkg+/n
PxHNa1dzBC3k/9QupxQhNLtugLFownzeawAG3S1bnTtKLBSf7AoDxu8/NC5xBCdUI+QvsXmLoOkg
WjwxxLeXMwWHew7UrQvFt91aVv+lR0phyZ6KM+TaVVKXjI8M496Gr7ZMF/Ti8Cr6zvdh0IK27XN6
B2E+9P8tQRAbnYd/6AdVj9zPpA8N2t6SL//W4gHawfCcbKojlmEUPTWKwaxutWjCNGlDzssjv90M
ZQgeotAJdcNvvtoZymLysiWYmscdaUua1RrnHbLAF/PkyA5UU2dTQ/Stmycgkuwl20RDy/jKXEp4
eVz2xJ1ctJF9p3X/ywQ8qbfZXYwTart6XdtCtFRutFpMAb5Jcmsz5meEVbNXeb1LAavjYIYbXHOH
2dihRd87xAlS9n4Cn4XQMM2HSGNlUfJ6I6RdySFJ0nxh3/5o5e8MxcvnsqwNQFDo5sp97D+rn0zJ
5DZH406MekyDcbThvB10wT7kTvVUfC9c+PoFm+vIVllY1yv4kvsybWj+ptoOqGUCY4ID8zQQcsrI
+plcHVyDRhD1u636vLzbUee3Bf0p4Slmt2zbSCxmHo6EuB84DJ6mfWDXeI9BFhiAwU8rUeQVu3iQ
RsZfd7YEjS2aOpvsF23CgE5JKpzQMk/b0hdiKwsS47yKtKnjPI2VwauTv1cvCVNSoDoG8n24dLZQ
FMCiKLft06QDiRTSL8snw1RwjJk/BzndDvfH3q4Ty4OM5iQAflsd/lLIUHjr9daZelc0rIjvP/yU
2jWyQSD+BW24oUmzeZn/HkrObPc9e0MY/928i/BgxTpDhikcm+r3gyCnTcvOZhiiZIwrF+uv/hrS
4nhhhUF8lfYjb7p9R0k0Lw2W9Ll6NZvBmYfwjVOwlxf/wqjTj9pSUPE7684wvVETfcqmawOpBux4
y7rQkqkkIB7irMFBEO98h2EPG8/3l16zstZcvkk6/LuNBgtjWCSF/Br2yLUqrYEEL+OatxrrKMh6
jlE1TsYXpzmODkgixj19kqUT4g7oTkoAwgjLOXHRDhXGLRD0dk04msnkAGJBP1uAcKF5g8tjsUmX
suYu529iE9NE55aYPPm/hIQ+yaxRRFbgDnhKJLzV5qket7aW4jyYzlOf0Jxere/JTMUlgN7INvh/
TlQvP4Bh3H1qBomnc5as8g4ACuhYUbOo5rbb96EMaW1V8oRJinmVzbbfrVQsQ/w81pusrYoVqGgP
hIJXYcM+DtyCUqRaADNcTwR9B9OSCYkzG8g8aKN6iFP/hdU6ootGAB7U01B+R+6foAB+N2fMtVd+
CtguMHiV8ZO1iEkYEcQiVjfgcswrwgxQUN7zerqXsJgopheCdoEgnmjCmwjzvQmQKKq68jqPi0fq
/dNRxs0NoRkZ97Yd8yZyh1FHIv75IrVf3LCXYMUeiY+FSG+VGc8rJTGUiB1UNWSmS/narNnJ80CG
WGZwJudMzHxY7d3+XnkJ87yWSz+roxunwL3ePbH7F74fSz3r8HbitBKEvRQARbpUSjJeZL3Mfh6Y
UfJTYfh5xWJ8B1gTNGjfG1arbyv07GLzWkqdHicIcQRRipp37tTKrU9Zugihc0oSnSwi0CuUgZSk
uyjEyhaPmctBlvUpBmcNIHnHSA4MXjoNh0WUdpNOGm4WDiDZ/GliDSmwI7e1qmFYNvNDAv9LJ3Gd
lxX73yeuNxyqhE9ZQwBlbtYUK7oL3XSPaoekqFyYj7B/fRj+nAXj7u+R24fCjhRdeVF5+TWcjrAv
Ud8ZxLiNeKx/qW86oNKAFT3ZkZGYWyXh4nMpmAlVyTKlfctokKNZ29d+rY1dA0QPhSsXyvO7meTj
x/PfyeVQUWf84p+R3G0u9gL/B+Jj8lbb5pGQ3YvcVJrjIWEVUWiDGcB/kyD93flmHpMTBKOfEvZb
/363irAIcAnWPhemICtceuL4U/6Q+9QAxP8ZApK3SUbPWwbVwW4NUzX8MbtNz3h2M6tY/q/HxBvC
m3Zhesp+Auds0xNPTpBFQ0iq8NK8PpdTzwEMRT9i+UKftGlxqpiXwS91bSd0BER85rbvM5ONVztF
k4AoJ6YJe+m9aViPQjbbAdD5OqnWygp+6121dEplKVu0gTwJvRqTQSEdZ9da/VcrwYhO2krvGkwc
jTj4ZnnJTcGMPnzB3TyVyFytwt4YLH7k1SYjaYPA/T9gINBTjlDUdFVA9yN8nRS1+XICiWixkuRM
1DKJ/VXqctim9uLT9ntdB3zCmZ3gYbttm4PC9aQbKbv+CNCWghSTo6shviezUQYZg0eFDYvDgkeX
Y/5wFz6q9sWCV70fzQf19L4+2K2GV7xlEbPsKXyy4WuvWYKhq+UbIqMDZaSeeSogYqfnRhYyD03P
Fw/KcTtW90mk+Tx9abvdxZiX4khog06UJLoBekifgbaEe9YYZJ+4BgREsRRrUqzjLhaTvFlYdP/t
06TCeLxnvIIANoOmijaINKJWkaVsktqYkjXL9XTja4BQsX6R5Eyq+trtIRklT1UWGrPHfH2Uk5uR
84D84UYurYn3kZuPmDQiU/MSL8kdteThW9at1IvxuwGU5xnJ20zhecLetiH33ZfjL712M57FBOYM
3NmvtQracdSPQGu3xtZulIeSXFd6dRZ9pw0neeW+IlfNRLxucp4FR7NbraIg+Pf3GIafyXNczU74
mqnZTsD0mmamhmT1QHQNk+W1e0tNdqF6UMMEiHmjoGdom8lA7UJMSLhlYbwCnqiy6rqPwcsvMuIh
3fQMBnqxBCWzaG1RR21BKM4UnF5nD5upROwsAJE1KPaR82e4IvUqeiZpJWy2oPnwtCFLDngSFj4V
Ln2lvoqYzQh/gZGPnc2dCa0GkOOVH5H570TqHfifZRmSDU1dShcCcdbxEW9S0kWaDuKknTqx8fYI
ksJm1Kt2P4auh4GzTdaFssy96KImazVKquOOWoeuuvrHAEVrGkDe+luluhO+0PVsUsLKTM9gPoBK
HJrWEDVi7dr3xKbvbefVbZEepg4SYCCQBePsrp2WRK/0q/8yg9uZFsRIJ1IXU50AChSbNy2r0RoK
A4oloDVAQa26U8cZjd3YseVdDAuM35fGOBMEE7utvx1NFG+RyDS8mrzUB8n9Tv1789+Wepro8dY9
HVmfEdgvgPH8SdnkK+vbaPTLhv9RLLAYewmXG4xXB47CuvQC1ym/mgOMXe3X8CSfr/wJT1M6LWwS
C8qIYzC4dXsG4DPEFpVXzTj9WySQDTpSELqbQrLc8yFCs6tUw0ezR4crTx8RZzQGKsg4QGC+Xn5D
o+8p1PwziRdFo/SHCR3b9H8GHxH340+OCky+1+kkHgt3w5JeG7IKrHzbvPaVwFdgj2KndGT/8G1G
QSXr3gE3zeS27k0izYr5O3CXKyDk59eB+Gh+8DFtYma2s49rFnA6FLPsLgtebITPrdZAdUukkMkg
+BB5SxWBzB2FRBsT72NeArw++c04GF8DMFeUS6mba2kkq3V3BagBee6vg6qRZwAZIrs33/Fm7OfK
sazpILOoRlGLTncF4SYXnw5zeRhVFkXqLhzW/4CINrsx1Am4Ps2V5vGJ+9qclXmHfYdi0bqNJffm
zEJ+zb2m3gZmiWv40FsF9Tz+1aRRaXG8hWVyGuLCgn52UTNLDQsrc2qNl6daJGkXiymK8xlO3NB9
cIOcgxRMaimAa9Ybb0XYIOPMqfr7Lf9Ga4/5fyFRdQHYKzbZv4fVqQCZVRsZhbl7O9WNWnZTNur1
5Ayvo6d4mx91kUSX2DvdqcPVvLi4JEQ5csFyVLGwUqetHsAl4j5YViuYb9Ma3cQl5BqusvqXAk86
MHq+0aZ0LSezV05gwt5nB8RBP76N3bXqPLUb2xB858tJuK6vDf+t3NCHYcOUQFS/VqvwaNNfN1WB
vlqxi6ZL/TJhmGuLdCmP/PzziE7OjlSdfwQHZjtVS9RjqR4zGmxUTT61RCz5KhSXngOzgzqjskJT
nKM/NC530qYVOFLwzKeb3fVyU6pO9IKcPDB8UlLgSJZ69c8Je6X7DKblM8ORN4fAh1Q1k3Up4nvv
R5I34ovBRJh+XsnRivLc0hR8E5wDgnRb5Pf41nz0hTb8GeKLfrS6VFDJq6tJlkzEaEM8TztcQAZP
xMjoic4xzKQuGewI3MPDyN0Pax7ZjVElut06A+enySZJSgKAigui5q6DbZiHKdUEbnodvDqAwnTi
dX27/Z6U4M2dHtMigYjqKrQgCrBCkF9/wGgcJbHuXr+0wS+aFNXiwFwIuJYIaEeH9ngzeJX1UcBR
zJfioKbzRtUf2OLLyOUQS3EO1NeBAVIkdrlPm7HWt53q66RsDh1jrGGOpXKS8lxToyCZ8UDVXL0z
SWQBv6lKd9TOP3i5PiBFq/yEGL/Nxl0IC17Gn9sxtdM5+XqOEtlRNdjvIHiX71Y0Kp43oJFp8Td+
SIAzKW1m5jBhU4QhKbkTjX9K+Q5Qrun+MMXphYRJ14ud616f13CQuytN5BYRwwfvmijVYX+EiTd3
8rRM/KX6mBthPATapOuq7Ar31KvkooGS6WGBGS2qqNacT348Ola4ccwpiDTp8+qz6peJF1AOJKXX
VEYG+CYUBhOgmu6Eh2VPut8NT5N51AKcbptEirI7HetJkh5+5f/KzTTaFZyUxxhGXhHVdf+yGC4c
ZOvTG+e3qkLM7LQhTeXO6aitmUJClCMMPoRcCCgZBkSbdBHXnDByqVDmTLD1VEsVbWXbJrzQkx7S
47rjpGQFdbqM5juURiDMzZRqREvZ04Aju2nFVvgm3WgehT/PMWEA9ErorBLNBdmsq8rY3qwz6kt0
4ndOX3B8/v/8q4CC9LciLtcQfZcYLMyQEydUM86cd+tSHhylfjF3ELeLA//x/LovLT8tOs6wcqDx
5f1PW+1ICssu6PRlbeW5ZubqGG9bl0bX0/HWHx9tQ5ro1hP4T3/7vOd5PVWaPCVlUySGvpymQQ1M
Tj2BWns2a+Eqx5jkH2wjCqGfuBOTJbUOFgV/Rsy1C8kDu2p3XRyx/cYvQePXZ/EVYcyIiQ1h7J76
txsh9D7TB2+GviwtBuR56o5EugDuvCIis8xuKPlkPvZZWPOUi/e5uEefqox5qocs72PvRjLhutfk
JnPjguVJkA52QjkL06zksUDeTG0Ver64zxF6SoEgzTnknihJfe45GYil/3kxDcC72uciPBOWnBZv
TS6naZSZx59XJ4eAQMkFDKu6FzcPZ8N4wf8lfFqCqXxsy+W4RPHsQDYcH2qHSHGxZddnTqbRil9e
tIQ2AqJQShkZbF7Lbu++H3qHcREqn2WcnpOGaF/4A7+sB7B7LDwuPlw3wVImn7dIES+sn/56dwdb
N37wGIKx2gQxuTqvvh3t87y2h3pTqMPluzedZQkAZHZRbw2XVS5fQwcYU+14ywUd34ZWuirpqa0y
xJgEbsXodJ5qShyN7k4os/3Iv4dfPhaZoB4VTGjWZmmqNsaM+79A0oaboFXJKAH2yCnQtmEzMR92
Q4IW3L1S9Ry2bBgDNphkKaLZq3KwRUlo1Vw6GaoPolnZUa+YAVol7vOQQXkOboyv7049Mf0dRLnn
zl3UnGd50AJ+bEYbbRgbHf0+2cJvAu1pKDemLDUPupiHuLmu6EzMaYMlijGbD15Z/Su3Qz5Fx19/
k5VN4Fb+BLii+fO6aA749peVgZvPfGR+H10OSjhLWwAZjVIULXNaXAEDzndDVGgd5IFkFdtnAlSj
CqpypgWoSBpCaUIwXjCiTrkg4OA87vamwpphf/PaZkzZo+P+FcbNYCwi1zsIftOnBL5gvLz2C5GQ
gC2b9IjB5BkIc86SyQd4GXnDPiXYEjAwSlQcWwyew8m83eGwfn+w+RR30VRIWfSoRb6EtD+CxGqa
7LgHbv+kPS+kXzTWqOY3/ysNTOusgS7y0VPgdpHFchgto6IqfoOba0O7t41T43GGjlnKiGTKZwOV
eiH7PaKhCQNAELEmgx7L6SQLrib3jv9sAH1BMd8YlPH5wUDqq43ykvSwdWq1zQ5yGr14TkVrrkqY
N3AQUt144bbuuq+wkywUoIDA03/iChFkNqO3pDXvp4igVnubyyalw04kXGLGagb+tJBNouG3oJS+
ZJBNIDD0qF1EjA9qpMO8vbrpqK1b5STXP+qNK27FN0BOCVqhrL2xJ023sbMp9rf2bF7nRJ7eHZjU
qgKKWkJcpK9mZxocpdB3N6jFDbvCMWtAfWE6JF7Z/h1Kq8vfCZ/zZK6/IovKmeMx8Z6OOkxTotEQ
gGrWIEhp7lvDmOe/rVt861h+7Jw5biAj5UVPNfaO9H3A2T0pNw6erCK2d/oeC/hke4th+Y9ogFPb
y7QYeFy26LEbTU48IwyRVQvPu7VV/110tZRjDmEl2n9M67lY3zBwsuks4GiGnp6rllc5k4Wrbxkg
L+o+vEa2IrgsUqQi/K83Lu+0EyltIYXb5sHeBgLQePLZjpLEQQc9NXE/vRsXAYj7hn8IrPnEZx7/
x4RwcMgfsZEb39QFntUXel9P0YoAPBvMMsjV2Qr1CtsJpkSgeUGeXFbE8H0P8TZJS728hL4PRcmJ
vUzpoitDPmvesZPO8R4I14GGmTCprKDNeV4VFkvLRLNsJhTslbeXEP42ZerdWkB+oB0WFLLICg4m
qbDd7ZseIHX9BBkLIvlqPEm/hj8KkwJeMNq+zvh5A1GyNR++TzagtwH3h6+ntIiLjWxc9Nir71Yl
1wa5qq6pfuUOjpZonpx9/YgLTYiG+PF1M1sqvcZPM5VaytDf4LrH1l98FbzIpVJJCgnT5/eE3xkv
3ADMsoEUb9EFSfbmtsxOvmtaAr5apQcdruVyZ2S/MIQNaFfaMZS/FwR0HkTWJhebs+kJ+0SyYYcg
gZLiF6tT20MKKqdkWARfLZDd3iPOHClRd6b2G7jU8S6GxjdIh0oJ+gUeEHYuj8U4EPm83WoxGiXr
hUeNqo+ZyodVdIP9JWg4w8oVzLxajPOD+NaqF205LHeMkeopB0MB8EVeCgjjgSVVp2blVFbhDuE/
2XONu4V1602PYFRON3p/Y2FvYG+hINoHwKz6NPQXIHvlG9hu6R+zD7tENInHi2KC6mqhsISPTL4Z
9EexU9ANn7gFvZkmLzkhf8qx8GhltNiMIBwtpnDRNHu+83jqUpYCygs6lbreUhZ/BQo9PCmxhs5j
PI7ZzEfiz5YyJ+aMu51OVUk44GVhSJQW9H7C542y3H2N7lrIhKYLGfpFo4ba8fx40+GCiIfyQkVO
HamfmpBhTfkv41ILUxy0J7hN19VYfS4WeRJi/TBarIlxBXDjuCLkpv69ZmBn4GiKSRGf61/LB2+E
Mqb2sCm+XmFyWQ9Lt/pttBhppedGBPwqn178wE3kMeYRn+mn3isUUlrmtlwyo0k+MWQvxlmFd9pF
fGQvS5EZzXh2AQmFXN/WF1+v/uVPg6PAl2cjRfpXulxXeUr/xZLaWhsQBiJUFCLTzuRvajUdDzYM
bPSJD4Lxw5PPR6WhmvsxvJ5dKOv9U7EcWwjryPc8DfgQ9dyo/vjbSfpFQru//n2ztgDconmGRd/V
7MCiLyyYR8ZnRVnmFkJjep+q4XJ7B0JpZjaNbqm5pdpv/SYbZoOY1eDslNhd1leyiTQvY2pzd7S5
J9jZIdCSvk4Ea6WTkmVISbRCygvispwwYwe6Anq4FDmVJnJqK9nH1kBLC0lcNHnqWf6K8Q5v3M4Y
IxrAsIVs5fu9vmYU/+FBgMnm+68vmabv4sZlAz+wjuO2GtFWAJg6GnlPUNqTYSDS0uNOLN/a70BW
7jIIr4UTvKvMCkHQYGkm5BOrAwPV84HRPkWLBNLinUJEKUeUy//o/1LqjI8Qb9Xh8vxIEL8YDott
0lUwoY6AgBRdDh4zSqzsaqgXIA3k3KCQjP9dfyOCFe6dHxeRc5YmMaWpdXrXcxYFp3m3foV4wCSb
eWBKNd4ip3r9ntP9RCVuMf8s+/5NmcJZFhBtQHWF8gOkw+Kjh8ut40w9BRrA23fDhZKAB2PXjxxr
IVQTPLOGcDegL4NrqcwRz3QBCylxDp8CMlOJQkxx02ewJnQ6UyViSE7Hk+IIg7DVpjFU7aaLOtLt
75159drjNTA9XSNmdh0GqdsgWY+RuxCcP0/GbRFuuPc3KPxQxN/GJbwuWV7tw2RvhGOpkV4Hdmy9
SsEbK98Cqk+130mCdizAY3P3jDIBxCVJ4lqWYRBNljVW4+1uCsBze1aPxquEMIMLabxpX/Inkf75
E8oDLoSxFEshQ6hfiuOiCSzERBHC9iFIrvsKuSGS8ja1OnAdaK5CHFJoyvHhbcBOuHzFQzAKUflh
0SpMFcW3e5SEadjj7GAbqANgKIn88wk1xBdweEHTgPmL0qP5Hx0h6YtYJlflM1sCL4yE3kIKw94v
8pDcBmJoUA49bgWNBkQKRvf4HdVEUJtD4sct1DwjmD5CaId084wDzPPCLw4eSeW+KYcnPDvBu04V
0Sr4EL11Zf9Ck5sYAEh7iYH8QWN6urX7HaWfJYLyE8sDgVQ9P+mO9rqWnYcQkjzhIKqJq4Xor5fn
CkxoricKgym0LRML7/trsledPhwF81PMdcjEHWn7wQ4nxlEfHW8K1lntdoPIW46QOSC777PPq0eb
kuKzD7JcZTkIm/HXIaQrgLlvADEAbinXUp2Ar8hFHbQVhnaEe3B+m3rA4WB9JEAjj+SfKkgvZCR6
aEcOulklRcoOvnWSwPaK7MyAz2UKmWYkiL6DQJD27IHuSZ3fkIXkDXK8mdZCNMVdzeW6m5GsNA8Y
EP0+uP7A+YqkfoOum3YRFysVXKj3kc4jcWXeX6MqVjLfDaF0qRY1s4r7joDViGBb6Cbce4DCs2r6
XM4VWzP0t9ldaS4i3c86x/fg0dbODcqOfSQPDlmXP0iAakYQw4P6qOwGkuZXPO8+52KO7XQQN9nG
oOcfgGsw3HKhxUxTWGuJSOw5vnRL0lAaJAEiCVM6/5UjRVYfe4QS0h0UesGSB8ixoToPT9/o9Xkn
c2ET5CWYq1yOgQQOsj3bRdXW7pAbbJS67pl82Uhb+58Hh32clghNaJv8FjiUmRQLgcJz3NMpwgiZ
d6BwFZIi1fSFNelyscpeAzfKWF2dTGJMPVUDl/wtNV5t/T+tGV9AujvZJGcPO+hCqhD7Quf+aKmN
LJFTflvILeplXDaV3Wb0bcXp/wP5LCuf6YjKemWT8OJpAOWBzFyhTjjP6naHzDpTNIX5yCqKXo99
q3o2+aLDJ4hJPvj+KPAGLzUcXA0m2plTZ3PvW28QSPPPGoGgMt6gKeKAz/GlCuP46NtYuAlJV6Iy
4M01zRQJrHIkwlxArUoX0AQkntmDy8oVX/VpHnz2eU0fWuOjvFOYW8hXSAB6kS+Cc8DGDmBUX0xP
FoS7G8dkOG4U4REePG4OCn4rwgOjI9b+r+gwd5AHmkWv7OSI6nqnCyjoc+fVJoptEFfNNRu6KbsG
icN4OP2rmaDVqL1OjJtcVohsg/z8mRu8IsD8xj1govBdlozwNnodLCqzUONe7wqrnN58lbh07w49
DXERUDNgy8Uif10fKSR+gIm3+HNXnaRvUZmOYkeN9xjT/K9FIvrRf4FynxX8Ik9ve/O2wB96RgS4
VcMNSRVYTsek+JpEISvG9Rv+Ddt5/tmSRL+IHIfOoU5ENr/8Dk6eGE0V6wVME1yoU6MgtjB0rJf8
m5qINuYmH1aXG4yMs/MA/uiYCSSy52gLl5K3X1G6C6V1W2K3hrtjkFI2Z+pD+DneYun5iEqLNkdT
GzUTygG1JY7u77JyVPjik5hmqA3EWld3B/CRioqkFynGB5YRErmx8t+GDlPU5se7XDE1P0a+t5XH
f4KA7hGaquhMh7PjdhoLqQBxB6PxQNhxFSrbrFWmphj+5hm6yoTQ6fbsXipEtPI6kHMk6oUBk3kt
4VJ6ammu0isw2EFxhQ+PjQK8Q/C2QlwOPamulUB2rHA7yoYO6TZw8g1mh0m1CclSoieM9pekunja
asA3+ok5JLVssl81/U5PuSK00Qy0QJVP7+XDR4O8FzQ6JHx55DU9N+domgW3gBANYRiGcEMjoKka
Yk2Q2wQVlXPMASHgZOq54CnOc9JJ90XJRrB1ZwzYvK4Qz7d8NpGe1m2qJabSRWJha5ldLKgbigAS
1knI8o3gbCDVd/ns7FMHGRDCde3+vUyQMhUPlxgPb7EXXY/XgDumx/oTOzYAKOQxdHwYP4WmueAY
7sw8S6qNTcIKQ0HtY0zzcS+ImB0lsD+4b315xi5d0rugAqT+BlAx7Hnh4mVLI086ll4gvXkKbvt4
8v9GLqBWj8NwDCVQMW0vGMW7MW0rN3trPnw903QNxvRrly/6x0tFXkTCohi0s0dGvV4Dzadc8B2P
R9NL4zT3FiFY6/mGU6T0sr5eQWJZYcEEu+hRkUoO7ad2DlK3HWr2dtsPG88Vwr3/UGtwxuwExgDo
ooFkV590gYWpzZoHVuNbbtJce4/5N+XbHii/MfUTtWR8E9arym/J0MUukNi2gCW67/ta4aLsUdZN
i6zVe5Ch3IRgPSljNHJscMcNKb7TXEUJZfBwQ6zARI9W8A7B8Gr64tbM5MNbFkuEseVN6OKIMJJr
H5/Go17WOUlAvppRNfzGSVJclKO4+tijJpBvFmE6CvG81b5rrRS8EDhqgyikzX6tpN/LqAOo3r2h
5D28bqJeUqtEJ7TMhTOzR6P5t/DRX2WYFqmt7VSI9c/bHJ10monv1rHeoNcdhnoYQmjVLjWdeWyL
q+ZS5DUQKT8ab8Be1aBbsuy0GcjhpHQw0XUae9yArW+QAK3GKJOxN8RgniTXXCqhH5hWtuHDiLk3
wA4AHQj7bq1A83q3b0NpZj5mFOmA44kD+O5ebt+aJdFoCg9oYhgCDNaeRpLGiWiuBRNDoXrHQeLn
BDO6d37B09i4wkSvHbCp33mRPLCKCXaHebtvpgWLuLTDfVrkt713W9ZML6ykFaKhMXaqJ7/OyCQp
3fw6s6DX2HuATj4eowrjThCrzB+6rdx+LFl3y3c1bqrYCOGzzRUmByc00lg8FG2Spg6z4C2Am+k5
iTtveHKrmVUS7T1ggLqbb8mgVxc72o4leds3PV6ff/sXO6FmM8J54xhuu4DMGCOj5zdDoo2j4Lws
hpbacT9lttASmXaiJsZZDv12XnQSvHPQAw+FXAwOxw3IHGs25Q/S7aDQtb9H7sT12E0x2Nd3H82W
PwwIBaOElQ797JH31JSJKA4+VCKYbu8Hb+aDW9h8gAOHgCiJfO2/Jr8TwHMt2Ix4Ary0qnnh3W7Q
P8J3qEHCHJ6FNV3+I977Milv4XYaK5HJ4P+aFFIUWZoy9B6BN7XVfZf/gW6b99T8u35RmbrydItg
hPTblSo7mU2kjIhM8KaEXv0DW4MssiEVXAYmHDrMmT5KofDRQwKKIR0qqeoVB2FEDLEudwSNgFZr
8Sd7UMW+ThHEGCK8kHn/HypzZQh0I4pwSbGWeG3N9Hpme8/oS9Hq+neGNq1hsyM8eiMNiNwRGrVU
XDNXkZMxGYQBz37l4HRKvoXKBwYTMS+GlT67igMYcJRUO843hRYHKANEQwbOck6Au5GO8MDwI2WM
1w7ooWcx+jexfrFYSn4fId0swEBNYvsi2oy0uJgoXfdRb7cvaX4t7Cq0xdgZ3G1lonqPzVhTDBjS
tb0G6Pau3wpV9nt+adZHrB04JqzMyyWiRlFIGVAsomGCd84EFaHHoaQJI5tU10vn6PQ6BzQShbBM
QMA6zqSQxveuBQP/QTZwhszgMi+WXOz7u7HPT/VS03T/aEHFgoi3MxsVqsqm4UlsmxlmQ4DBzO3u
iSEVuyLXg8Czb0sSD+fx77TbTsz/aiTOiI/8hEIgtnDuxX0N30v0xEywYn4lSen8+hHPGNKXEotn
AgIh5awYWstjUlXHHAFrud87lFldYI77r/mmEnrEzrR2qd79aCKRZqZHCSUZlDJBF/WPX8tY7brC
2uCeu1zZcZbHN3zvlLGRyl555VQLwXY92vNyKLNQFSNRQ8fxxQu+CIE4K2d9BWqmQqgx/BPu9CBt
CnQaTvogcDfFgzwd+4+rt+RILGTJzdxm3O72m+OwGyYVr0BQn65fAZUWrHXeMOAVNj95567sPAP0
POyQMVqcyEB/DYq5SF8+4e45ER52xIs0kMlsqSAMVDEoK5AbqIjQoUyz29GpSwSP+rAIl29ESFoo
W+xbLocrfhkDce7uXTnArMT/1TmBlWpsYRVEPIV92d/E5z7RbGk14rzWjg42wyKJyvrZe0RkyxLp
WS+hTDOTifVOdvr0DhuEqLncV5txzr7J0OSlW1y4tbpxHyu9bIyC8LxZ5WeF9SjNlcJnG5lf/DO9
Tt3B4nGW11Mzh4v9qv7lpb2LKkVcKq+87sTQ2tcxpqXtfVub/YHVNv1wHt3CXiBO05xXKCC3i2HP
h5HIqesTUzvGXRi5+v2CrRAwn4U5xMu+kJaD9WpgIFfP0bn1khlLGFuSihKmtguhsc8CKUoNGG1G
g5432CxU/L11srKsaF13TgpTFME8tRdRzENMze5lUtGH+RolrsiZCjV524Hqs2hCILq2xUwkAN56
O0RgIw2Bw8awka1GZB3BE3t8SqlFlhusFtJpYJ6lDrUisITJnktj3WejEYAEj6e2k4Sq/x/JrSTW
vj92Mvrgdl0Uvmge0LeZsIufOSiV2ok80BBZeE+nRxDfNsTKso8pwsqKKwBKrbUvMW/HYGOriAPE
xV5xbfIaJ3AULXqu8gX+lSqjimYBmDjjDQJlH4d0RnCF51cJoU7nOc6F8ONbvCtilW4APH/IPS7I
TEgKbZPYmZ/Vi2uG8wqWnjrKgtEFE/uI1uI47yBIKirtNv0b8E3WZpF5i2cuVLd5PvjSg9YsN3x3
YdJ8R4yAxiOgKa7BuNexh2j/hJR4ebYt4OD5x058ne/ESikkxRrTnVye3DWUipVWYw5njTk5TvyP
HIB+8A7LvaSZr0SVcjQYJyKohbWhW81hlctcSfhOuss+UPmeyIAPs/BikKv9OJz8GMsTpV1O1iLK
Bb9Ik7nq5K/MC5cOwcmQcmG6lOclWw3XMcMlLGbQTMGS/gM1XkP02enUnaa+qghoVuAzlv+9TYma
eNOA+K99Gq/OhApYivMBZ4vJgMZKkOr08XtcxZZNxj7zWPiyrnIt9cNnMqrYIAtNsgiyeOt6gUV1
wBMZTESWtR06LN8DIYVzSsF5hI9UUhxXkNo+fArGknqsgBrVKtDzmW1U4kXXsWm74XtlM9DbAtnu
sIwExHJnNLImXPwRlrebSABwb8iItmYEorntwu9ayn3rM03fcjczZ/djjprQNn3uOjYw7xGQZ+Eo
Iah4kppihswdradIuUqoQrQZlJyygFnEQO5dJEkd9zuu6t5miW/VgRMUGhwndeBWaLlMBpg0X6sJ
ioPw3LUtZtUKX4m9gy30RuGjb5/XamVyaAgLpsIZ/KvezO/pzirBjFirf+cg2Xe0uz6FJ6tiqk4S
3sset3c4qb9th9HDyc8pzIFRSO6AJi1XJzAXK+HjPCRiWlklGH5Ldwcx6O4crdO5Oc1J9WtKLsaH
KmmargNIad3oVRUwRTyjbGxpWIHIy+xbcOXga7YR2hj4OU4ic7LtUFOEhZUGrMg3lwULI0Mya598
W5eKnCO7J4JEEwBiEeCby42EnUGRgcMCmhDwebFAxQGckxYmMy6SiPpjxYDCM7CYVIuMhvTfa+l2
02yN3AKaoA4Xv0W/CceA1ipf6n5o2tsnHxRdofNoflh6YB81HFk/5TUy9n7m4zb6S2GkrrIyEU09
rF9CxtauSBwsSXNI4VzCNiMOcTXY8cnoTpvPcuF4Wgubeb9wYWIMfELBLrOn0kKWJELKe7/iPTKp
N1RBlglTKldi22OUs+OoSQaRWgCHp/xvaEKvrkOZ0LXSMeUDoPmY0r0ia70tu5/DoJVdkJlDbbTC
Cm8SUM5UYwJ/1KtSrSB8hYTpYKdoOaxBJo6V2XbW6gPYcAF+vSEk2GRwNY6b7I21jArxk85X0Ykv
iOYPIJm8qZFyEf+3aOrJilDgqFhGrYRExxyIBZGFSPsSpZJW8URJf4UYhXed4Af0ZA6pI+UaaD5r
4m0yclGRe0fxwoRhhEHRnwWiaKBFk42Zqs2XDIhVJmrSY2PcE8DjmukPcqF8iAGEYt1XbLXSEFKa
d2+ajDw/v/lPfcS6EIRAeYuPEp1gmNaji9NQHiqLF/+tF9qJnkUlF0A3dLMbUmEVLcouWpke/MDv
dt+1jVc+KJ5tOKZGNXWDXeUlrjAreveiuRbEb0bBOlRoSjn5jTnJShW2U+FzU+84tLOcy/bRAL3x
v8T3CvFG//+gWDcmEYXCVlXQJqG82tX7t7dARtE8rF1XRkS5i/i8UPICHyrrbtofYAGNaocowpdM
jpGZ54uXfK04yxgbYnDn7TRXB8L2etnbbZ6cm4xAUtcxXfShWClG7BlaksL8B+IssO+oovUTLg23
ynkQPUfTHjJs7uBndE0W2ugw+NcJH/B/6mnTnF5zSe9wFy4WNv6tNo4HTq7Snuq7MqKAuAQFIO8J
/F8y95314gRnFWqFhmL30I8j7ms3CXdmXqBqVsDtltUaOmiTUDGh2gS6ZLLgk/3/b6mQlCCRx80M
/7hZwB5ASlKLtDRh1n+M3y7GofwoITq8vw1Qv8VfmmmVrWVFEjdFfn012xeXysd79CLf6q0swm6N
qdLqiRZ9MA0MigDrDwzdlTR0hPzVndH1EOhj1qPQljJVbBzOe4v7jyEsOMEZFgaFMMeAMl0cepRX
pxO7TAVCAiJLI8y/YYxN0fpd6tNPK9SmaAys5GrrpbRqWgamfwSNEEvkxvadeh78C+cojZ9+vSjA
W0k5p0IAtm+JCivdRjACFyEhseJhdcDhJ/OByO3/KRCBPVOcD7kJX5iXDiLUSyAaGJMMIrk8pAiJ
02Q/CBkemVkI7PzZ48wb5xkkVQ7Mq1Pm/MIncAshKMwvuEnaUQZU5Xb/IQx/E64PZU1zVqdFvkPM
JymHyPdmi2W94tD9wF+hWLHeiu9Y5oxpt9/z9BFpnMneTW9jrJ6E+iYPpSMyfHHhifXYwMLnrQII
aZp1x6fxdxBTvoXRASTAyX2m///RfTfSJ1+bCABQg9pZgdGi5p6RduMu68K9jmu0iN25gcBR8ExB
1ppzSlo743Pig1tQX9mUPLzj1+zDz2cnSHJLkGB5QpYIlxkjiDzMKTp2hEG/GYQqT4taeTTGvTJD
/ZdkMYyHtGnyyFm1VrM0+o+NiFaALTz8IrEWdTXSkLKoNsVDQ4jWTo5kUEI5FsRAX1x70rtLlxuG
lzvexoX4xjyc6mljtFmbve2PtKSIZTzbKHDCD1zWN7mMLSvo9etAks/0zsbqt8H02v+jfO02rZub
qtZ+97R5r37yN2NpZerwpwFP743A3KkQ95z19cljzWohAUc0ei01qG+n6Ay/fGaS9AXTdJxcnNBV
p93BdrIV6iNIZxFKzCEbKccDef+YYJo7bJTr7brGEzUGXpX0BByMcXIlaO40BZsQ2NAmLlmdEl7Z
TNU0+TLAb2/naZ5TYFOgswIEYnrYBkQnf1RjQWAIriO3TWkheigXM9D7ChsewpozbFEP7784v0bF
HBWSaWgAoi67mqFp/huVOP1vbXE9WBk0qPMlqzvRNhN1fx9jN4of4mDpP/smGf07nB3fMl/95jZT
9lh2i1apq1hMTUJ4mnR0cQHG+SunW3lMIeVoSm55xPHiE4aolWCDUaWtlbK4E/Fqczojub81VK3T
zQMvHyFVkxNnKHnpPRmtWe+OLdBdfQk4VhpNzoxBGQ0FZkp3SiNjU/GZ0tqtqrVw3R59bGe+A5Ap
L3D76yzUMIO1zyIGmuhQg6bM/7ukCLkFbMH7oDn6OujDXLL7Vv5Wranyc5JHxIXGUpo4drtJuB/f
UJovyIy0hGTAyCaJINerS8mt9etNA+Xn9vpmsbz7TjUhU/Vkos2cidVwWSDW8Mp7Wx1em/xM6vA9
XX8TOpucII3UWy9Qd1Qw/EF9Yryhjh0huudj3iWBeXsJcrFkeuC5TE1bWjhbkjuaADdGWSPlsh9d
ZAOE7Sqze8+6w+BCQzKouJk4K3qp2Up0b37IVoKvTqgp8ZW9Mh4UNtA31mufOjOuTXUDrPodzDwm
x0DKnnHr1xMJcnj17srXSYi3XUjI+n3Oj52LLYHYzGV/FLo0tGE8r+TP3pJqDAqL5WT50O5qHdOk
k7J6inNwbvlTW5rQ8NuzxlwGzSJirLwIP7ClKESCKU++JYCN5lJF1MXanovWcfK9kQ7gRnVEM8Xh
1iHzAqEnJCRj/EqvXnYOdwoiYa6xXKwS4kW0S0v8THb38s/Z6RJbeOSkzqVBLLYdZ8KIyHJcX89R
nyKvQQgZ9N5E6RLYrmFDXVcp2lvnAoInloBpzmcHffgZZSzn6bAc+OXJ4nGLVnO5p1X6Jx3rWX2J
Fmcs6TNXaVf4XNgfDfmgxRIVLFyirj0t2/FNK2XrPSQr+qNTtx1dIzYS2aYdK1kZWX3VS0P5SVkG
onhGgpwdRDWrgQNOLH1Zkpfy2MK3/2eSkURB3TPr+wv8oXnlHlyobMRUmRBEXibCLrgPeBaxXooe
Mu2d2ZTlqA6hLVOMgc6dt9zBh8YLl6sDeJbT7rBK/YrhG0ZQqddj42F39B22wcX2APY9bm5yXTkz
Wz46SMjTt7YezkSOUowClx4i/gBwnF+Fm2KFEhHWCSwKEjPvxMxPf+xiWTcpepySgMcZjmPgLUHl
iZsXEa8bdnqnZcEtT05ViA38ERvaSWUkFFZw0QyrVsflfVEAbk0Im1QZTnJF1qWrXYGsO+OZISya
A7v3Xomrg1UCYGQV67F24lYCCOM+5liuJ18Bx1vzjWEctvrnjX1TALS0hwKEZR7S9Svj0fiyR2I8
0etVi/DztdovTYcERalU0VxV+drxQhIuvLKPUDjFbnEHnbVvtdHKDUpYOuzHqDCUMQpxEvweRGQ7
sdZ26OO5YV+vk3ewczG4vqBa2qvDFoaqNa85bCLTTfY9C3rnOgkYF8BlXoo/qbHGyvF4WT9lwKwa
o5F8Io7SKjfevu3UZSXny0toMPm/2ajFq5Cn1JLmFcSGXsQIxnVMroDc/JW6c5vXDiC5ZtqMufo1
Py4TxvxIGggurftCa3x72wb33TlxI6VLtkp5bSoE4OQn8l44FN3fRTA1UgyxcejDlieMVqyyXLBI
YSlLe5L3um3L0vxl54z+yjtRmpehcP7VW0TCC4MmTB3PhFQVrEanFXrex06fuXjmi0arPQBQUOQw
XpbV3N+lJSrYUUYXSjA3/k+9Xg+Fcq7I5UfMsqNc8la5Z/cid+kZXBYXv9HYdm1S2POAnPPYwBHh
lfvYmq4eG3j9Ybiag7eanncFXVYlZ8y/l+HIQ6KBZoXyG+uTouNyfMthEFbgn9wSds9mDp3Sp2Gr
d/s/sT3JL9e1V7cOsB/GejvQs7KB9avgNOMq2j4C7TwOIGB2xOtv37vxhfZwgWxGQE7ZRLZZods2
NsiCgBG5LiQxDv8CTxhC0pegBKoHNaZ6vcy58xLVDeE7JOOUgO//TGThkQg3go8SYjXsuoqN8+Qb
ZyFNDSxfbcWI+sRyrYeM8jHuN+0ESvcB+6I3bMnET5vWBYRjiEKMO7B1d0RANQ73UDTEoqlcpfSx
sJhdaXfNAnoKbdL4cZpbcb1iHxrFKkcL9EN3wiPvTxOmz9tyHtoxB0AVacKw6hngxDPPvJJmH5RJ
QO3gvcWtoXmikHlb59yEKF5sDe3Ag1aZE2zX3yvuLcZsxOHFfYOjOoJ72PCYtjU9VNysEfnuLhlk
dksIUk8AfnCV2h069orRLnxFtk1LGIVWRbIydtN9MMpGWWw9zuk/tQ5CS+O2vzz1osatmXjFPx6V
h1nidoiOrdgkW/TWc/sNYT7Dsl0PnrmBlmGRIvpsykZp0VNp1f4N+akHSENibEQYoUgagDkCkrhO
xTwCQwaLok3rI63ZP5RBCh9W2coRxJ03esX0mPImm+nPKA5QAFuZpxf5uEHQatGfe2QXCXSvABs8
cgfM8bzquhi99uW8LWMKonBNAZDYqgSPtusJ84NKhav/e942hKegPPPzYaIOHsd1NumUnc0dgzWK
RFQlaLlnTLemmK5MNwNu5PtaKlWFjxmz4GV0PD4PdviSIXUSbiz0snvtxnvT+1RGm0drzbpoi99h
zP4JmhAfHGiLxfF8GbZjfrb8GqomJWmtzToqosb6GQudVmhJcyKleMHSdglnFtFTqhVcbGb2DCCF
83Y3v3KXdjDf1eJA9zupSyHlXkJT/KFktl2oNMYL/ILsMYOlDEeVqYf2Ehz7a3pQSRO05pK0Um+m
4W79zf3S6YT4f/AJBPUgfWT+Tu2Ibv1z2iUrxm9SbA82u41uwFAs78DrM0x6EvLANxRd+J6FLCgg
Zhxt0a568veGXCkORhSfi301IQjC4et+7LWOeU4+hp6xGXQZkweGapk5uppn1w2A+8weQ1D01JXf
qC3N0SoW7gZYnjVAe/kLzW/cAlpuRUDap7pPnlqhSeHaevL2w7PvWw4StYiTZaCxfVnPTOzeJkim
OCxd34Ymb1xZdnNMQp+iZPI0rhFOi45Smv8/U1jnOFB5gYbeSgSvCQMN5fbCDKE2fQGlqnEys3dO
YEHwVGkzRl7uDDGYLn0fHXreaugssJTZUQZoyoB+TVySYWy6G3lgMr8OqeoAUsUhjJ1EsbKbwNus
gAVmVSeLdALecxHu0DtT5Gr6UTpIef0KoT0kJhAksZE6Qhm9cIda50gSXPjgZiwCmZrLNG43nz9n
uBZ1uLU44n2IukKemHwvOSFNtfUPfjNx48F02tajt3HFp/icA1MXSLaN+HLkr5dK6KKnpNjst8Ei
RAO+Fvlvli5R+vH4w9JxyYkXpoRaYxizuVykkyUBlPibQ8lDcAXOH1QM6QQC7oNNgpVDMvvReHq4
YM3hWEfIfgj72E9mL4wY+oX/pukBqSkhyQG4YHaGdeRsRrQzFuKfY9gSBALwjff8IhtnTLaUYhmH
2iW7CgSfqIPS914vA/Q9fVce9B+am9lA05fXl5FPDbtdY054l7waf3y4FwFMA9cqd5Cc9VKL9c37
SBf7wZBlMXJgwLfUZbpQQS+tqm+nl4DJB6Qp67TwRULV7evb/0dsR0+OLh6LbexuyfrbrUxzxcuh
a/9HPZJ9CbXskxi1DA76qYi8ZQKUPqtHl5CF3NjxFmYqLzeRJEK7wwvFCDbCMyLeKRCgqqWQfDbc
aHzCcQzU7bgtwRe3sr0/179qraqxbFL6LebE3ynRt0i4fOv9ciiH2ufxCRDqBGJJZOKw3+EjMghT
XoXjklywZZwPD0ArISx9VMXnf6z6soLhpMGxTB1BtttovxMwvIQhsTWpLg1lfJFjiIULhkodJdnw
RMVUKY6Rq+EN9RXGgXu2AX2CSXY8VtGXxdeFvGcoK26iMOeh/44h8wW169jtiy6ZdcIJIDV+ZQhe
8lk3x6UB0QcqbOrxxgK4jZfvpXQUGE/heEa3j2Keg336cxbgM03kg3hIjnS7Fi6zSkR2ul4uXLm8
rVJ6ts2lipXHA2sq/Aso/gVWJUwcEE8rxocHwn1gsJVIhPgHf1N8TL191+q6EVINgnZuoQXHG5m1
pIePBUF6ihE+FiLIHgnln/nSWWgaOzUupUBOwvbUUwFVwlHynXSfHfUupuwJPYhfCPbwGTbou7+C
hzu1C03KYNRU8X66/KIDTROlZKpSZ77OsydwaWIoWOd076QwzbsPcDM6qfiMcNduGkGQv30jtTfE
21Rgqe73w4r8QJFpesimSNnxhuEQYpsTr1lXP7MprRuSKMG8YBVIHxHooPhK/Jbv9FsOF5ffLesg
RY8hvAkD4f2Ei9P3zbkkbfR0+cs2NF/hsNg6Z6A4MJ66LfRyDPDgH5pZpI6h3JXmzzWkrmhnwIx0
iKE2fwNSAHfaDSEaNcwJW8Lqbgfo1arLdvHubanA0iWtr/N9bB6h6K4I9vnWexJyPD5EIu1D8bC+
7C/h80aszTCAnWpnK4X/TdoYOpjD7ZQzpCx3Ng5w39ZYER7NrBsV92FZmYJOmAHIUQxcAa7+YXGi
eDg1TrFQ98Myy3Bn8g04za3RNE9aAErMgfVCBheaxVY6B5KIvp670uz2K8vCc569uxHciYFseA76
qVS4Vi5x3TOlNxCmihbMvaMm6WlgD90M1R9/qA1FkImobLSfC7azIXVk7HEwSHitt4EdD1Afkcv9
IGlKYik/vneQSaXkn25pCX1CCxPtMb4Mh+oru8daeLwk3sVwjvyqin1yNzwDThoqgan5BH2LsdIe
48gJWvgBmGJQ+ThF4IkWk1k9P9PSlOZ+8oy4HJstblIw4fHxamBwiUlSJcHtWJNZDO93RUaXdsKd
35GBZAE0FOTKBMwaHUMC+3ur0ux+SNG146T53/btayxONLD06WSDL4gDmSvA6wUEl59kmVtyZPEw
YTVl2Ji9aPbQrvfqoid4rcuC48ryG5niFBFDdbxdPALTr4Ck7WhsvlfpzmVq/lr+o8drvAIj3Ikq
4BucXq934pjQ/hDzf4WFWwuQBvI2zrOUWgWuvp2FVqfoyYVnJ45yIBbg5thVvKQRnKP2s3zckjaU
WwaijTIRINzHePfPBhERRRdAy9DA7BZv8E+AUzrpukY8H7AIx5DoWTmYUvJrvNSbX/Gc1UGUR1WU
3Xz/GOmupdWWcNgh3p2Rh6gu+iJASSkXdRq6hDLgN5Fy/fSXNNI6x4YQRlCIvX9AikUv31DQMfXW
umhuL9AQfFVOJByRoVJ02TT+pSLFAQuylHZU9c9ND+Vz3wrWEcVIv/uO8PJpfJ1qTmIMK2pRsVeo
/489ZBLgVjIwbzVIo2Vd7fs/3Jx+5FD5NFxrhcDSfaoZWwDZBG0r2ZaZ6MpMf8+bU4Iz3oRwaV4T
35CVY5u61HbRRwO6+DtgaYnKDz5Ux4SxI1mPot+3JdAEND1zWfr/GMf9TQWUQvuxuzoNIBpbCIzJ
6+Jgij/kb5JAUWRQRgSiDL6KaanKHn6wqeMuF1nR8tr8VDFOdyHVrtt0NTtfqB9hTRufHXer6/j+
SpQ+EoIo65n5IXjPphOsWd4ldqRfvGVqeeNUigS0Jg6GKKuOodoYC03ON9YijPyC3tDMlAdlFf1O
ggugSaACLBsrQy2LKrpUwMtcr58IncB8dJXv7a3HaFWJeDB+g7RSfWoNyo5J6srzjNPK0Z6UMlcI
IItZGi6+hxxM5OjtEJsZ32zFUYzzq7XBvyflJqXtuu4r3F6MRDOSCQCSROb4aC4pmikvUmC3raYb
wezDF9YRdXKA5wMx88OdK4Bi6lVHXtpwM9wMifOJ1awCvEp8PKqdrlv4dnoSGm2i8hhOnfN2kJ6B
ZUirLBcsLKORUSbErRwOuoPCHhxp3XDqqI941mZ3V0ByLThghxrk182mawnlk7b6+hiFj+FiKYB3
dhkfYL4+bFcKBdN0bHkZrxHQh+4RlI6gngB3OZVkiZR5wb/DsW5+eV19CGc2BPWrrylXHzqEMTdN
d9l1xF/dGtZVXgSrJuxiuTG2Wx9SC/qn6XUlWiVYJyAW6EfhKpQNUH0f8ZJLqCyiPcGzcsBLxq4w
qtNRckFyejPJHtjzeg98WGZeZDDnHmzqCNEJtAM+CWNFNS3dLi6I3GnmXWorrH1pS3bY0z6Pj14M
AHraRvNrFvZv+FWKSXR70uJoaJ6ZNc+XkC8g/3m66F/9mFBHzbMi9aa6NOLlxmdfkH6QtjeaXWwq
IfXbnDYJI5Z1dUekxU3OaJ4rDpNd354IFW75v98TirZA29Pc5vlP0yoVlu1/6wwbwjT9RqIO/yaM
P03YUlAXg5y3rQKIGKth6V9ILGaJ/iZ/7VmzhfiMraD10QtKqEGQyHNDD4MqvHTKxAdnTC1eiXpc
dXxFlcyQhQeJUcFPTAo8gaKksAE5GjV+5c9NfZd1sp/Medg1mQxhEgz0KVkSaAPSDfTudhrv+3a0
asYmJjU2L01VJ1/pRHmUvzmjxxSyAd7JpLhSy/gJFQQI3kOB42Asq9rH7hhO2FHuH6RR08/L+FCH
1CKlxUxsgyhm5ITZxU/d+w/5otD31bYmwTTZxLL5GWGue5QPglZh4Vr5lhZJWAvViRK/8wWr4k6P
xn4pJfuhjOrjod3DZj/joOtIC64MR8uKneb+jXRyRk1vWOpMqj7cjBcUhsnHrsjSbTg0xg2Cuw9H
IEvq/xPDuvJqk45Ucfzr/bhEHjCkfy9rWqdYY0tV527ZuLbM6/e/lUyVg4FsrhgSKlEwHfiFKWgq
MbahfesJjGP6Ei14vbTAcECt0bIDzBNzYajCmjzV9M32q1seNlZ1a0y8vWHtpoMYesetLlqfI6Gw
oenfgPEpyxRFP20VHUyUQ5m/AvcaAxlR1EJurIHacmYtfgWImV2ETayJSzuHBJbrf52vAlokPYW8
VLJInKm2wM87gODd4th+6/9cXf3PAzgQegmZYncu4KpNk1ov3Ey2MJQMANLsZl7ZaU8SHhAwDLaM
Wo8kYEi5UwbNLZ0KKF+berY3YWu2iG926Xfp4RvL0jeOdU+IVaSzTWAujF3uMxWCvip/E5ro7ohP
9pap4peA5Wnau2Nfb98sKDEQYDNBrIcJ6mxQvd679ujR2ZfmXaQei81aszxUaLZAAEVIvqeJIDBm
JNBGsnd0jZRDZ+FLde8tsWdFIZ0cdlCEdKufav27g24ILaQgTlbfEBbTEccK0aY38RT+PgY61eMw
QjLK+whd+hdYkteRL1gWjXjEx+rTis3wddHdE1RvB4r2nIQVrfgeTXTwmxFd9Ydpa33Ma2X3a+F1
02vZl8SWCOdXxKG2AMliKg2Qq+u3wqNQHcSRRiNSBUq4+hVq7J9wivWM26J1wYt/Nb+d+PblK8Na
Ib5Sg+qt/ulWj9vD7D8d+oaF7k0r6NnhDRL4LemsFeptM6y8OMzSzIPqFH/YRrvbvh8iKI6BN2Vq
g0xMA62mqYcvPQgzb+U5tJDjgk8mgt12APVpujj6LQzB8skkOg5qx2nGLZfy2JsFr+5MNLRVdY/k
9phMUjAISU2KEu3n5Lm63LKufk9bIjULvv1JoZ/npd4hZeVyWde61DqUgnicrDIRGueQYyjdNnVx
RfM5/FDkIxaHQP9jOGCiHWe08rgos19Kz+twnqDV0Q6zEYDthK7aTrIac4lQva4KtdPnz+eyfaAG
QIrrfDmj/XHCmxCBXMBklG6n4k9TEDSOVcBePSMkjVsOES3OTW+oMnXkJ620Pfhu2jwfOFnKMm5H
02O8dJbmD2Wqe2r98abCBn1knqkvosdwNEn8F2mCWQoxIAC2wIWgne/q+l+YlCDa3FdouC6iJgI5
N8INhF8VeMlOz11cT+eTRzQbQkGY9KYnWNYZipXzVub6+XSro8bLjcBU4EmEtWsTA3GmPBK8m5kc
FZwsBKfe64ln0x+87XsKhee+CNd9uj1nU1G2x5DRYhnWxo2BMd8lH45o+6r7zEDnbSaQIXQE1xbm
4StV4mFFVh7C2a33uZdoV8mo3jYo+dsqcFzFyOMHecMq6uIX4SKZGYbUr5sNXZwcRr2iaPk4in1i
5oC9NHWf1kUOD+B5nnrvfRgQ55B4hP4CZHtzVPvyEPVDiirkJrNyqUzWdJ+dnkvSSVRzXwIwKJkz
wRXHyDnpuaQJVJRHeXjoa8m55mRKhuZIXBONrA2iJzKK6MTbVJxZh1SSgxTBEAoODStpX2R7TmcE
bgM+rdmnQEwngum/YWKOmWTxixkJXLHNwMNjbNWb3ukkjEyCv/obL8Us6TddLYG/jRu6OjnG44KN
933f+tn7QZ0z4Uqx0jZW3ESDmVJxQgULr5Pe0tabgIUSvxVJGVh+8+uIIX5jG8wLb5yu9EWBx+4I
BwZFKVn1DDdcmrtux0TAbdIbyos0ETiMOQLuSql5eIDHKkIoTgfqmhc1LUjMddxAljuS/m9DEliD
FEwpWdmhzX/KTZhbT1qlsoeh1g8uqpR8AB+LPKqO+Vgzc21X/dJzZBKQ/VIb9XTH3Qt/BCIzXFfB
1LZKcZG2jwGmtfKpffdfWMcYBjly7dNeHPBg2y8SbgBQuiTuKjlXDywK88o0gwS8pJj0YEHCE5S4
APn1lxYjsTzspjdb+Rbgbil4A10nC6HDPWidg05g6gKVYbI89yt/S9vLBfyfO6/9z4pQqyqIUZuL
xK1ZVGGmqY5rXwwILnlYFS0tjuegZiYZbzTjYonULAAMK/IAUtoAlXieUvVLjz8yM1p18Pj93mvt
FiLQFBabrMU+7XLw9EXN200vnh2eTUyVU21NtHLrhhf7ww3T5mlDSJkPT5vunRuVsZ2hEspYHIFs
/qtF/pf/H+rT44qEmtHFXsV1VBhAiL/ANLZF1pilvDRamL/VsLav3P5DbwA+e23LGer7rRWjx+DV
J2YbqeLTZIBrGGflGvORI5+F0yoyHLqkcmoiejmncZbZSBk/KkEJQXaQLN3Ru5E3rcu0NIwjBDxW
aOKFfwFQWwVzePRnsmnAFs/IF9RBNsSk2/fc4Crq7Vib//IyP3JtqUEWs6bAdw/ifuHD3SWbM5sX
WaiVknkytZ5r/uYRwIzScwnWtk+RFXfS1oXAekiuKqx6VRnD+7nekBqajEnwxQ6MD/oUBlaPJrtp
63PId48WJU0IrVxLNRVOpCAOcP9UNtVoKi7tjOb881oTBhrfbE8N18gNbPrtYacJ2AnBeTtMyrx9
b9L8NX9SQFm+HF6BnUTXpz0wsYhSjpUzDB493+YEqwmCrlh9MFkkPecQDNFeNaEEhJH7uqfVzX0u
3Dhr4NS+iRY0Vob5zBMKgEWZ3ELmb9V/G1l/cirUNdTAr45vF8ACa1wLL+/2BaFwJTBzd7PK7jBu
oJy6B559xuVA9Tev4CskCmYsLSrZOoFe/Gs6zXu8lCFplSQlATGFPrJvkfjd7Ooo7s8TEVMLVUEy
0U9vqd8pditl0U+pEFXKtzWbHnujQHbtujK9rBsp+KNneuWuUzDY3BCS15BDjLVMiHjGRC8eA6+1
l224rJB87i5Wu6z90PZiaF9/w00nwHaYs2SPpO4ocJg1w9efFIU05Key0FMtP+ye0f98PP6gCh8P
1g2eujYjn5xr6bhTkJn/EBmJ2vW8HAsbOzMJnJnIETEqOJe/RhRlJ8zEztYp2Z+unyfe4Tq1HpSr
YRxjmJV0ps9NV8P6OPLGPtudeGnhobnWCncMgzLOBiMZ9eg7bPduWLg0JzPn+bWqFqK8CUgeu18q
dyS/qIpFvU1yLzO0h4qjtToVebmBQkk/I7MQcJnnOwEM63e4HGKvSq0qrlTsGicy2dT25x9Dku59
w8/he/sVA2jzPA8ZDCUnK3q+x+cyyzyOv6JBzGEd+j+y0esDjZ2fJ1XQfkXpXDPYyHfX7oMQyLkS
zWRLC7COt3sFCI1gTmTGij7j+Yb59gr/LMUx2WsxjBmx9uSfHxAwv1DWdfaR5AVVOAVQE0urkcyo
rPgcMx5mn0N4DRFydrH6TBc3lcUJAJxgX+Hi59RyeMsNbOIMmFGEt2RpAwiaHiq8yvb27xJL1+/s
Q/pOc2/GzpeK+IUdbUfA3n9q3v6jfvSB52aqb/grFYbWoLS3TPHK0PYtKdL3aWWeCEeWsI69U+K/
TogGCXnI7EFP8QHvK6k69wer7y3FE1HEFgA4qm8eMZvFpoeJEAMSKqWqrJPcsBWjP2t/WQfV80cw
seSJpdvAcKWnevLg+EhoXLoN4PjZVNKhfx0tJISy495DSYL3H+k+GgaZGhN+XDXUI0r2jxsyeOPH
+eEkqXcnjl2gR3mzxQFU6aaMYBJA1LtK4WQGCkbpPI9tkcRNkdeb/9aYJqOXYLOKJ9xQui13wBcx
xo7nsVOMl+6plVfga9h7wqJsrghbB4FM4fbCmSZmoj4LV8A2VvoSVtsPH+rVDurKtuu1xXoRX32c
SRs0DLdnQiWVOdxDeMqYNN3rDZY8h6/K+LHaLOoGpOgEjsnZLp/02U72CWDfnQib7BLr0dU3H6Jz
f7Z4CBCEEyDFlE93lT4JbuFKcZrYVOv3nZUqeEIOs+G9Qi2vwa6xSNGuCnjJL5WhOk56UzQPVTq1
6kXwfsZ3hZCpmT7MdrsqMGuNCPjStLSOI9x8SE5SKljhcFy8LvhUULaAKy76P7TfFaGj62hWTxuT
Rg4XM8V6jhS7/0XfgorhvxPKA1ctFRma+zIjvP4aah/wrU1QcjF8WV7r1YIT1FvemoPyF1DSoIGI
fUw8YLyCqvbGKdY5biTBoxbP4K1ANV30FqRlzU4IQpiGd3jo6/aoV6AwDnn7eyQ80L0BGCSGdTNg
fLi4H39EGV5waZPW6W5oK4QRhX4LhgmERJP2RYuc9ON9+7fqk9Z97eoLK8iB61nUZSslsQgiaIgD
bg/MYNq3pvZfjg6hMtlGb3+07sOs5FKAKRgB/E0w7T29Gswo4tcLuTeDpuTWY4aVYMqepim95Aqi
wP1NhhMz17Aq+sxwP1g6x3jcsZuZKMhjmfKPqCA4vGTdBmJr9AuMsXujeUu/bfmUIFw4vFj2tta3
NCJguwydcWMrGkgVm7MPeWIhqY1uaK4xKj2zasZ58RlJWiIn5mitrKnPnPVaHMBrEBTCh+z8d4eP
/Qrttnam1dC+yHfzvVuWxBIFmrNPY7DLFobP3HedBoTy225ycP2saq9nR/E14Xoz7VCGg+5DmyMb
My3wdjKoLOmCD2Mbhz+2KdkJCEDCIAzXAKSF7plqdOhlAc5G8LDJ+oMW/GnhQsY3tgFRGLuovcRo
wnu0d7kUZQhQ5vlZA3+evLuXzDtc0zXfsn6cojpq1uDgkSlRQ8YbY8xIHFp7dhB4+/m5FM7RY/pn
5y3253p6HMJoHWgBBFl5FoknNJKxC75yGd+6/ZyIXpVjR2RxDSrjZqcKg0eGd6w1h49b5Km4vF2X
yokmqAK1QfXu25Ys8hJZq/xRiPmr1W/ClJ/sOEGTReeWthGlU+6Hhc/cQn7ClYwEs1bTvo3a8YUI
kM+HK9VsiEBq4pCrsKa0CIA2/nqY6H2bhq5tBxvNV7US2AsbO0N7RRjQmXCXCXgr7kO+41THgwWU
nKK6IkqfVmpRhxw2rljsv6uQeEaggpxvJsoEqHmQyLgFuIp88oVR7nwWLJv9JsHKNIIMbxrhOIS/
NPx9QArnGX4yfo6zuHJ3otyyHtikO1jbqLc5nunX2LAmxqA2gTHuJOCBkDAHhE1i3v/XrVgY8e/+
X5PXPM6m1dLMro942dU8Dds3jPgTuFKiVudKIEbWwakymMzN9zlmBmzbZskfrIMpVjOeNJV+SUt8
itYCaWsEpT/OqD3NoUztdYqAxYp2DcQlUMuxhufkchK0MMUCpNKijy0Z9oTFLHe7wgU84lL8oaZz
0GqSdqw90rP/B2ynPXNfTiieDqImmEbG1oXmzG/O4hMef/QrrtggFIcm2wT1Kut3l0zHVY4I4k5D
gblDs9uJnGTYrCYlYWo6+6nCEzweR+wioSS50pk+Fu1OVFko8Qq9nYxNcKIurfEDWQxL5+cRhzCR
19UxY2fvnrUPpOJQBdsa5XfS2PNo+HGzxFojPQgIyg6wQQVsMmaXAD0K2DrdREzdI+RSKqCn2VG4
edwlWrb4qhpEhMDFr8/FecscxoE4YjgbJjSLP7PC9okjqcyRvcDJfXzjsXeANcJKoG+fDUcl6JxC
Ftvtygrt6gxAwetj9fsmzH6Vb5LpCx7sCkfZh5XZenaP/UDsEZZg+Ll0bj2QXPZCmJj2bzCqhX9t
9+jCMf6bbHo5jzva+N2Xrufq1o4GbHujOpb3O1olpaI7qq5PCuRJu6K7ZjrvGH3Mx1R2tS+DwxK6
zDLxLdedFMDHj96l3bASQyMJDl9MjVquA9qblLQXlUkzjv1gDGwWxNQKjXKrWGzJEJRSVWB3HkBU
gqs23dtyOMafYaXFnUo6UkCsb64Nw6v9pUt2sQEPWIYDnJMFAAp8Id+mo/sXUU1VLmpN50/i/bDu
c/ucJLMx4tVfYy4ZhNx+moi4B3uEqCCU7W9LKyQCBYvzLMVANZ1Cg+SEH5s+vcvKqREyvLWjqkK8
bi+WvN5o0LyLsLLExedspOLETLFXY4co/GZQPKjhXhIUdGITHZ+oW5dCH32YUliVrPIXTN/Y0iy7
K3Q/ScDsxde0q2lAyOE/C8ayQwSdIpyoc20lscdfxlS03Rx/LPRXgFa1gituG1f6mEGzdff28r4H
UuTSPo1W2VNVLwCNf5IqU76FOeoAr2jVrPj75nb5gXlk/LFwCo+FimXrIUHIMW0RQoqsilFPb5eV
arIF4gLMMCC/HN30QnxQ5ppu8sLdbpFYE7OCy6ftqsqDwrMuVPnZzL2sYOftFJhi+bmzHCbCbpWZ
unDISeH25g9Y/5q/oXYzaVVEXJWCA4coCUSWDZOXmQSMkZ4vKl5e6Ux0tYggpcUdHuSDBJZxTe5i
HX/MhfILrt9r2GrHPTKJ+zuO6NilATUe6YpctueD3AiENV8yC7fWq9YG4fc4jsZ7T3t8vWhn6tXi
wOZiKtz+cJ9a2ZmoSwrN7n6V/RN4IVJn5HG64koWCVlCmhlbZqPoIPM2rkS3O1R27bnrkNOJaLXT
0TQ3SIc7wUv2BBcHRcOsK5oYEbwMk8oG9SnaKn04hOKadUwLn2Tu0HzRc8Lr7Sbp4t97GfqRDoXa
iO0x/fslI7maMebZoKiQ25qxGFW+CElPI5FPz0xIoIiM2u+m6uJf3myu1Dhsnr3jXE1o1yL7jIz+
i5yiBqqPDD9UYmecdYqpFqczafSokpMbi9RHExYZGl8DraDw1m+r1fiDmue93PBUsd1vT6S36El+
EHbh/6HD3+ntvdvm4Gj1CqtyVoesY7HGE7fXdjQ5dw+aF3Lib+hNsr3uIh/32qdpntSx7w4TAm5J
NG2JpAgLU+1SgiJdaMdySDX/p0ohlP4iGETlscxsODZuzgHtGDw8HLe6ZEpfF/NHt5y1dE92j55l
1txfL98iQsKEd/AW0iXZ3daNMl2J312z4Wn8s+6pQiYN2eFQOSEYjujyvVHBkU6CK21wLSwj3xVU
uL+u7fzJ+vuo4Bf42sXu6vbXOM7+tEZ1Mv0hDiWdWU5JZAV3wE/aFcKkQb0Vv26Sueqhga5Bv1hn
LKLpfgTIPecmb0lFcMtBWG9P5M4d78pJvopQhqNKFEVjsddbSKubbwtUoTWympAY+8sQ6Y7xs30j
w4x1bqosQbZX7Gl2ug/b00evGLUGQbe4tGwS/Vj0zEDFXafuT7a5qKdvlnbYbDgCHlxxNC3DePO3
/0MHA/2CtITkdbaMiFemRVn/gRknrmwLbXLi03+B4QZZ9EcI7Cf4pPmmkZnRgNHxApjEDIG7ueHY
2HAOUSIswl0oS9ohJX0fIDujBVnP3Xdddvkh4chAIt7oxHxAsrGQuL++1GwZP7YGVkADdlq54+Ak
qn6J63Jlg0Ma71QeN61svSqA8F2dSeyjWNq+kN0DoObPD0rKqN+1NKzxjRL4k2WzUP80K0W0nKLg
+0F76uxgSJ4/vuePZKp4qucp1t3ANUmWnpnCqJ11wf/1v4XHX6JLjtdMf90/fIDQhyAGFlW0UNof
HCupjMG4BxkyUS7xibTXi+PptWn56YFGc5TEKWxiMfGodpd7y5h/qLwN6E7jTm9i/4YX0IX7B31H
wHV25CTOYllaE5TOpIgxFuNNDMnprVysuebJFamb7N8SLrpC/lEKggsbhTmV6e++1eSfmSfjjgor
nTtuqHbm+/gEglYFwj1hweRTXcJLIKtlo+8TNJoDVz4qY2HuXhnvW9xzUaD23I+yLVMd0x/PIHPx
z6uAEFuVDzOovbDT9Xs30qZvz5Oblg7o/7cKu6ZfYzoWk8QD2E4qJe7p/2zlFXalPPnVZS3xLLDH
YOanIpRJjqLPaLWdHwWk+tNgkEIpnFwrSLK3MfLjXVLKKdBadFKaidVOOBmhAzTdxzb+8uvIEfBr
BRUSw9Jb/68pIVnS1vHgRF0AeplDxS9L3hQhluLZ2kddPJkZnklJ/E+q3UytBBem9p1Yx46bHPFC
14o5wrlNFP+rDobIlIzaRFHo8l7BOZ2UVBbem3v4ZabrahOhNibTHoSiBX7jkwP7kkYOqiB8XGvB
EJlautNYoFioxuB1bRnUVjkarcqlb2n/9VcUwMiClc9+oj0iI7yDdQVkHZQ3W5PF+iOKWAB0xceW
TAOstoueQmVWcB4QME/PXWbj4AJsddR50Bvp/X925ZS6c80KwjpUcWPzu6QQ4hyr4nRASFhCo6r4
z+CVOaTnnnuAXmZkO+rSK7e1HlHfjnFiaDfeERhO/wSmiGa8+K3IBukwNMyyBBj97DMLFIgLuUgN
7j9DwGEfnzjoGpabXfAX/IQakWZNTYAPTDmiC4xWVXc1Mhqw7UPr6BBoSTGa6GABDkBUcRack0eS
C998H4ki27J7ZnPFnXJzHKojBwWipvucAh/G+4EZhVNi4QJFRy6pv3S1PVfh2htnjt8Xy13AkqPB
1W+Ez6uihvVPEZPs70zuWatF/k+2bRrql752P6PwvS7XEYkrs8tj1xhUgjzhQXNV8H/e8MMdz1zZ
JpdJXKxVoAOzlXC92Aq0ljKyAXxRaeLE/7v8xjC+fdGrRwqwJxOfc+D+32un9H5s61qkrmJkCPoR
vFD54KnTBZHoKMP+9Spqb39jebfrm5CE65BaR38cCrkTZw5+PjKgWaVOpTeJz/y9chACOT+0ef8G
tJBp6MJgFJ6N0/j8A9SvURTk67XfH2YPSNQ8T0ATJad5VVa4SEts3/ztQ2Os/jrX5Vw1Lt1vnxD+
Brj5uP8crdKv/zNgedt1IiIlu14jhSeslRvdublmqj+uRpbXKzlMHe96JpOuyN3RmUa2QQReXZP6
upqMfOIItEnqFeQCPu0CrFx9k3n6wD9acuC37JJXmtX9ZJrF3R0CQ4JnOh2YqZ7Fu3ZowR5TD52k
Ow4eoNaGJRplwgAhRFv43G5YrIzNedzJp92wyhT1reVXX9/wHh5eKqE+p6d55ieDXIkU1T4FHO6j
NpJtm0/S7z1TIo48Pfgw6W9WcStoZ1CsnYIZpQvhLTrR5fEYAr4ioxy8p8leoMXbKPQeIo3X/rUq
g3ERLTMY8gZBw6qh2q9a3PY1e7M7TxEc7YAVjrhHgQ9+LusVPWRrZX8SEehkoRSFpVrYU3o4WfXu
5NtprwFcWBDNnbTm9Q05Ms6EZtQuC7HuZ7sXw6HwWLIpCxlFpqznOrH46rnqsXbUcu0OlmjBJI+K
5tJneDJW0QAyWMcta2M+9y4puLEm2ygL36mmpmb/PiMN0LGbY6aNK4aNR815Mc3VkSKA9hLKVhHq
iPSuSuq7miPdf+2+ygV57elvoLLzuGUd+3kakiaS/dKKdyARKgtNsdS7fNRZxGZOoecA5Q1gmfb5
dizIvCxe1Ws3YPUQ3pAh0IXvt57Xl7JBq9mImpiTDxiO2jBMFOq2aemjbZ2w88jEudryqzz+U9BU
/1aARU3LCzyZDAsb1ZliITLpRRpP/73Yq/acwP+UeOZ3TZMUSGp795M740nORnG589TC0kYcAZqF
HnQMZcU7BM/B49I+6QxUEGrbafFXW5Xe3IvRmD0twRFlhFep/gvp5MwieGhctUNDBgqca6bYMb9e
2K2SebuWdFWyNBd5eBN8NK4pC4hVIcakLnPFEWbJgU6Ms24DFSgD9rEW6Gi1BqjxsewiG2ZYtnGj
Y8IAE/Tgb744ubS+kL4F5viaO0TJgoo6IrPEWORKntNOmq4BwQQ5CUiQ8yJ9fUKer60Q0dw1uYGh
Zn3EUXxQDtY7nSD/+yIfTGGOAo+kJYh1p1Y6CkI5MLPIBtILRe3LOZZvhJS8c0kMTNhUlDOPunv0
jAN5fs/SnMCfc6HysgyVIwC8kV5VpLyQZmtGFTyfSHYikl0lTqUhp+Oi6WkADhMmC7Wca41Fa2+q
TAnUSRg55zN+NQvc2b6f+5catHGmTarjKpxd+BlNHJ4CagMO5mxewmTSliI3hhQnfTU5XmOCdf3Y
ml1/5qy1O1Z3wMqAvRo2G/kzI/tMhQCO3+QAylcpOfGtTq6305ipg4SrPsMM26Rh7NVhVcewKL+x
hDRvY3y1FdLpKFFq7haGOM7mthmo1dahb7uq7athAk0Jxdb7YaXXDCMSdfmQ6F7tvJQa+qUPUw9S
tJa7qLzG9fwguxk9yvsIzNR0V143V73dL2IxyathdP5dpSRKMjoL+JBnokHUkxJmVrkzclDWDxxM
GajKtvf+71+orWxv3Ix1C2sZv/qOAIagctHLMrK8PFcFD23IPlxqexhx/tkdLFOCnRwcyjxzZSmw
NqRpvzn319PKtBma1RRqliYlk8BBX/lSqoB8oP8RLWrcM2tAFKHeuNOTHLSVvR6V6V1hXC1vW1Ro
zJX4l4yig9Z6OU/rRCxp8Ll2ga52zezXQyxqUlfYAz3xkNMd1RWebhC1sk1om8cMAWyiTQq5hOIw
lydUzyyGPMwC/MyQWbI4vG8XtJ+SpoyT+UiYRDV2usmF7oma8SOWDfD+b9dj7/o1+XejZH+b34X0
zIc67rW+qeStCXY8A0ON/sBl/tkCf05KOEqXh+LiaDTXwufgvKyHi6BQFSFoUsFVEGzg20p7T9TP
JsUhG5vsgS+pZrAJBSryP64OcPEb9f2o4Lv4xQfzhBieO9B2zmPEH42Cck7p8FoM1J8qWK0Kt66F
7UKuq7sJpUGVmi2t8rJTGjKFN1AWkS/Zabun0mP9Pko+lpXwYcxbTXQiv0p1EZLR3G/Mka5SVmI8
BWj8DuWanQET/T5apnTKuAFjOaI+AjHGO1wDzsZ3zIr+EHDKenAU5ahnvlCjDYUwonvDv5BUvSNE
+DH9FacDEAIj6aYkNwT5pVkMU/8/cN+V9ijSE2x+E+zoseDGmUoqUUINCsM+0vtHxOC643zx7nAC
zYHvcnMSJIq6R4CIZn20L8OY/fhSnB51bhddPa2pBFY480wje1lre410zl8fmTRT6s+xBikiBCDt
I9Ore1RlAzctNFXXLuRqTD3OaIh3Sj9Kd+MGuJEKkv/WZdlrat5xzwMqMuFtb6W0dVCn4lGaURO1
FiTuPk/4l7BLn44OUs82ycr4BzhQlowDs03JxR6UhZ3P/b8mZ+Po5J7N75ZUgLXJHHKPe7U2F8KS
eSv9sYSIB7+MRkWASA1z0vcgpNQHrTf5vuQmRkmW60UioEZBmvycgM35/tNLVF2fPMzHB+S6bv32
w+TP5uV9HzVCagw+UQTtuJIuUhhKutq3XxmYKpdb0xhWw267CccCT7/1bCEntZBosQhv/C6AyDpI
rIUbt9AI24qjUFdGrneNbIBHF5qoMkpzZ9t7qAnBBJbDE9nIx8mXXGP0WP4Y2nO+XitpgnOh0cDo
vyM6GOhtNjRS1e7hTLGdR7EtEUjisNzMJUadxY8cN1LiRg+7kFuRUnU+h91+A1vLmRhXucVYaNrO
iKcUEB7pZoeuLub2pBY4seE8B5Wv5RQmz3uMjlD9dVrNWwPlo0cHwAMiniEbflqrQSfZJLQYx+ah
SH4H7fw1Mx3FMqPTnsKTlFrcu9XH7N1yk+AcVCCnJU9LizbFuOsgX+F9IDBzorFIjmSy9vo+5Epw
ZNf2THbbXI7RHmCyVra8Z7+H3A3+63yu8RbiUH5ITc9RAva1NZL36bvJwwe+K0uMS4pCBaf8YpZ+
vC4IrexKk4sy3BAdVeXeDLg/Dzsk8mof+u0Us+t9HqliZ9/gcCFWZ/yUInispbl8bki5Etg6NQyU
0qXUk/hMQxYDgikjYLNobJeP1GtvGOrkMQ5bagGM7F9XKVMXW3O5flpcSGbzDSsXdZZLjMQ7efRP
/znSvp1HevcviJhPJYyXwAfTcMFnS179owGXfiyA8GTWBC3WhGC5Dr2N6ol1a7smNRSYSn2LuI1C
+pHnZoAuwf7eNbr8tK6Q0hlnNgQJKy+evi873Lc2hXEhxbD6nx68FzjfOtUAe8KT9XwDY2jjIX7Q
LjR4OfbidD4Wja5O80Oipe7LBHKa7xqeKQkwZxEWufP89KfR6Q4vnal79P/zjZ2FY44L91tmmC02
qdFiB9X7jxdCNtX/NtLrJFaVWKolB7bDWgjFcw866T7x9Wc4dqtKUQZrg8BC3Hw8mgCuhd86ZyxW
aAKdP9I9yD6RhZ13WblaEimqtuSb9MHcrBPuDpvPWg3tS/kAyg594m+Zmirpw9K2F9FpLXw7sGVa
MroArv8RIxNtgJkXq+iXLnBMj3yqk8xegcnipWEDWjS9t0giXNzp2p1o9vajOykcN4JmFjtJ281U
V/bPi7OXFeZa8Ywb56ZHJDgu6gFr1YFKNAbFwoqjK1A/wgtNi9mm2B9+OFWhGSsFaFhMmNDDoZbE
akm7aVgJSEMYU0dBTtQTO8pcjWHq2ylrAf6tViKxgUJPyBSHiK3JQxjz5fU2N9RrX8wEeSgfUiYX
+tB+57slN9RnPRY4C6KTfFF16x52GIKsqLNBQhMvfYFKOR2m5dspRsrl+gYGh9XlgGdqzUyQXKAS
S7NcGlyGDsS66Sf3xjt4/V37WPfe2vinwu+xjPjTneFNf9CnNVHVePSQ+zv08JnYnlvwHzw/ET/e
p2Pfxs3p/wylqXVftib77AO9ho31xNtYPOdfGZvJu9gwMuUK0XzlE0h2GdB6be15gpTSTvfcZkLK
b+KEX7WCFgNkJB4cWVlhNW103wf6r47deDy0ujvsPlSwSJFT5qcOQaQoy8xwCfkILXhDBIEBitT6
wyPkBxH7GnPcA+GS0nsKRDlEWJSHaMUgrLBATY/q8MY2LLWyNc24Fa03gQ4Dcn/9FCBJLbO3S8At
K5JrxA/91trgQq+lHCsQebT4X/0bbMv4V9/19zXr4k5fVAGI/OnCThWDpVGIvzJM6eW2mjih6Wi+
elaMC0dGlsadH9RYbD8xX1Ul0QrjanI9ZaysExQo7hVALbd2RVDm2PXQ5WjZczd/R5p7igRGc1YM
P4NRVn20gjy0w8TTK+bYy+FaMDpTqtoM8TFSqnfSQk47SUQPjAyHO98TMgSXY4NIrZn/7hZof5Aj
IfCG+UG+XqUkmwXYTfTdAUojUWNDIC4rGqceEsAzesldD7KI+ZP87EtIhSlUY6ck8NjmNRb5OC6g
ky+5LZPJ/ZNg3I15ulT6S0o6yK38mAuPfOEjZhSa6/Q+w0f3NWvCnH9veym7Y1/bTSC1HW+aa+g3
L0HrAEPQRcGCn1rT3Ds3NxfD9gmiL8nEviyv4eOnniPeNeu+5RAdPq0nJ3LPvgg3Sd4CZ1whiKGX
V79QrY6YP9IAnDE6feXJYJO++BXQa+WGM7cVJqbJU4ytNjQfD0C22cK1Fju2D4k7MmoT1Iu0kwc5
5Wv2EqOphyVAfxwx9nMuojwqA/dSEI1sZ+gQC/e4ta6PFJmF8RooWCXgQdMfDMAt40z+t6skTFMb
9TwkbFQXEwvaIGR0ZbGxX/yaeQ2P9kukKM9BEUAbFatTbK8ueGS5dIius9WSGiPkT+S+Dtg0qvaf
oXTWVx3A9HVoAfxZ4dryYnuLmiKDKn6TcswtJYoXKUkOpzHLE5vOPXeF/Nf1QYpmdCGvqsQOY222
iY4Op8e45OfBw8fsiWM7mgbqy9b4EHxhoFMn22PfBDjbiugdegC0MhVvcST03KnfNbQo0TN27FFW
GykQmEUnk0pNHEOGr5xD/3UdQ2dbAC7FF89IJ8O1H1ayuBQtegkoZIDUtsRijrynVga8x7+xKKpV
bfE9bwLpzRHgHwmIXNSJryOS5ektQjB0wSvQIusoBAfPVJPwLXAIN0A4WdJ0oAXXe+T7iCv5rWA4
kc4PzEMqsZdbEbfSwXKWs8cjGmlTU2eySF9AG1qH21JkoIpBmfG0Up8Qj9D9dIdzhqSXs3axYRpA
wMe7j9/TT+3lN6x6neknrTllM0DYhTqxdRPzMw8pxKlgKL2r4sxnaDYgOfLBNS4S6SDIitaTwo43
BwLdl96xEyBTLdqi7tae4UB2V8VBwycYyScNjeJxIIlmgSKrTyM9UkKNJYFgXsLQmQchQMqxjKIj
KwmObdVzPFUaeXaizw8jHzNjctpEBad7Xt9Pvod+H370+4s/pMOePeEVhD/c4zDD/7a1TfbcRcKb
6mrwPVc5IK9mbB1Kcr2Jmrq/5ShMl0Jhw+sCII1T4wCBYhELKsbEzJlxMoJAQzfwr2GtYg5TZRFX
DEy9iQWodReilo1TDMJFW2xAdYqn6SHLlWjZdh6hE74KEfGUjpt4198rhZ1u560lyiWUCLAekF+l
zFdHgPqCb+X0qFsw7k5VmTofFzKP28pVaeZukrnB0O4aFSl/5HKXLuBd+pmKaZZVgYKhog4M44vG
WJ0Y9gjmAjfYrUeqVgh3fNdjk+NhOOnKbbu+JJHr+30ohctnidDWa7ADikGqxL0Vwwc8+4Bb6+4C
AzW69k54wHMtpDNxTKLd98Or6ECHnjHomUfcJ1PIyxsmrJo3QwXQeou7Gw8aEsG4VYAsUbkP7GXx
0LNmMni0Iu4TrLW3A9SYBt+bwokyH1zl/j5afSRoQbl6lGT66QRtkRCWErawAm+v6wdGRsNomlib
zEmtqxmRf9nLe0jt2/Ds9RfNdvZQuScv02vnuiBOdw3/OupyustIJEKKBCPz3UGEVo8RqyTn9smd
XcQ7JrNGq1RTosekjaKpQIhRJpbdlgpb80DPkEguV2IVR3Zz92Zd5hhfoGUMKn+2tyDIs1V8WP2p
kwER7OW/hDR/74Y/TiqVi+eu2zEenfcOLKcvuGFZQaXpCcNjx0CxZT6Zc4xrbo7gBS63LSVFj64L
9v950MFdy2uDqmonr+j+k9yOj86PCvL1xBdLe7h+QOz/n+0VGiFlw4UC23ao1+8HmXjjTd1i8adk
BWayLDhLP/HgUDcdsJmItmUdEyUtIRZdtKLEkXwTIThISwLD4DkW26w+jaPxGsGJCd8my48llwF5
AhiXc0p+tHZqNiWt9mmli6HxsZKz7ICXrSTGeBQ53bXmFLmJhI4NXFvO1wp02lrDQGuKw1hneFlx
GKuUltG6WhHOOyicH1z5Qfu7Ro6dljyWl5Pyf8bKK+mFFkAwKDfDFaNTntZ2n63wpAsvcJElN8v3
KogcMg4d27TBvNnU/5qXdvOcEVQbS+FIiukQQlhJ05MyAzBaccAF1thwD+CcObY+22bX1jZaBO0/
vGP0Tylt1UQAZdEbEx+ir/VblKH8EfyYhhCpBv/oHNnHcL2E8pnu9rnKsaKf37ljRTjThATMJW/q
4MDUpsLPyvM/CT05uyymLWBhf5oGd6C2xEYvRkNK0z0xFNoX6Iip0q/6JdrNqbQZXBUOFbhitQ7v
D2dBB3MDW4/XYMF6ZcCSr02MvRvzEYAZPowH/n5QJCuw77U/RIRG8bOU/kUdMPjToh5KRN8nHSq3
CJvJKKGUwNVEYzAKQJQLQ808XHIHoSECd37cFjoGOGloENipeU7hS2lnwcFDYMdGXjiVstVv5RDW
EKDbg+zdPYio1alLkzIFTVCuUil4jjmdMoPX/1eLvHLlB7WGDzPn/U5AraQkOhXIQKH/CJ7JS5wJ
R2SodcGpipbY0HT5W/RvjKItbOVroyOyWQaqdd4e5Gwl5pBqtA0H2MNH0FlCBFGCbZNq0wE4zVww
mvxisSMzzn7EwoOYSLG/TCM4x1SPmLu4qCrWOXT9pxhrt9ejpZlK9eIpTiywfA/HwlFfdb+ogWUW
V7UH0r9OYW1Q2JqYQy+WsremO8kcv4RwX7yz/Fn7VpJw5j1pAWK+ulYOLULlewF97YFYsS7e/v9d
wT8RUsGrrsBkXQaOA2eXSae8+abvqrUWj8WXM2ZMQitMMMGg92wPPYliYvCvSucU9l22j2rryxUj
6D5RunC2wJj4f9cPyizXbgXus+q1iK9NfehZOWJW6OSgbiyzA8ovCEhZ726qa75Iy7cyK3rUTQsx
65ptCI1BeWpTObSv5gM2DhWA6gw74LQJ7G9U6v12TqpND8eht/5nHAShPLJFa/pBZfVjy9Rke8eO
TUVOT3EeQy5bk91Ye4XvohzMN/GIrhYoysxRZsJQ/wkT2dwlzx1cGT6jcotDOvowdD01z25llVhR
mZg99dupQ+E1lyLi9mrYyZNNpqjE6jwyCH0VzO/qm5mF8AzhJV/qoT7P8Zb3iTQ25udk+5Cbd9uB
+Z/393JTrsxxdPqX6/cF/gD7xCocJqmpR/rBeiR8+f3LUyaLzxWGncc6Ajjg0oUpbw7wsWsts1d4
9UREdGhlgpBIMg3ooZdSUy6eoQXGHJFfI49hgACyXeDDMFmTgs/twY2HmaS9T/kZN8tBqAcmaere
zBhU8oYYi8wupFheTtjbwbNrWdcGli6SEzzTOSFdiAybXu3v8/ISxlvNcjvQKJK0ZlmnRhe6gEBR
B9HUfbNeKufALgfXQOt1POA6yMu+WGhaWzH8uQY6WkwJkwQGIhqlF9264yWY64XKd7qpsHAMq8cX
uOYkGP/JyxiozEJIvtBhi3eaFFowFBTAio1LCePMUDnUTomc2k9PXbmz4KGM/1xIBtHzEVmskJ41
YRfWcWZuJdDtrokGhy6nPU756vVXhNxaS8jSQFAUIHDsqU5XtHysWkrfczmKZa+Ky82G21vV4WwU
3KZy+h0VvX7Ul+DawDHgA+QiUTVlOUX4JVetgu1o4OPG/1EHZLa0So2s/lVRzRP23vn2TsSlXETx
9Lv1gI6nlTh8Q3s3/vERyQXFdByO22RWfpHsco/VtU3n2/e21KvuPZOBPylut2e0mOBkK8XPkjrS
GS6plVRY1Ho6TbRsG4J8KR7UeLsna2Yjjbfx+E2rYTPySdvxh49tTWOEJUDRezStuPkqY4MdM1Bi
NbOUv0PkNiQEv66IASv3nukhw5X4257+DnF/jq8iSdHzGxNdve9onbhPpvR4GlDqeKhIcv/FBRPx
d0N5vS1n6/nibrCrRDokye/yK4KNXckBFnAA5ArSUgwJECQvUd9HlougqQQXMSBXVsBBjdA2O08o
Jg1XZkqPJfwjYw2tPLHZJ4cb7XL88nBweV+1Nn7Kx9HFpgLWjf61QAx+Ain08ePY/+JEyb4ujvZO
8q/pM2eWx+EiUIvoRJ/3MELvTdxhRR77KrAmoWfni6TR0bf0Om8TNmMUNA8+YJ9YAd0917XBiuaA
NbBtI4uQkxy8BUKTT+65TNqzagqE+ET07X2l5Pqjyj5uGnJE9fwllX7odNzLzumw7lQmR807Mx+b
AEzf4tq7jS6sXXEFv37o0JQclAUpnbATi1rghMS93YrYMokPoh3eTnilP9VA0UIjzji9zoYnylCr
ymgUitdQQs7cm4VOAF8AG0s3iibzyfVo9RpmDEF6OqdtsciksAbt3BWo9qPivka6dmntvQ6KhMmI
FSU53pkO29DEv4ez+sZBMbft2kA7RF1CHpvkQ/Yw41bVWUFfYXP36BKFpAy1kBP+fVWUJtWM0aFe
/NvWXR8WhCUVQ9N43HJmGdjIMzXwOoHzRtE9PGux/Ih6TZqedwii+zmLixiWzC9TeCVEocjpoIxM
jOKkyYzWHQVjFiX4V1xkrvYGVmVLY53BXqlp+KM0LNCyzFzlg0defM52Ha2EEOaOJB8mJ62v9iO8
izUAwUinGR+M0ijK8npuJS8tZURwLlufHaqSPFAxYAjMXCJu9HvMxX3Bfw+hExg5LiON37cnQwQK
mA/klAyTFKKVZMIz7apy8tiW6dUweqBjtvBBOSydbrkOhh4Vy642LeK3t5zmvKMo/nkDHh3yNBqb
f2ShvSF66o0ggOUN+zakC6aFpGndIaVGDOAclzrSGkNf4K00GDl4vn1YwA043wHNeqritw9B7eV2
hbVFeVtvan2DYEHGyVLWw8yQsc/UCOzC9GN6zUT0XAK5O8KRl2MMEP+pSoHTcBns/apfxrTfB8vY
3th9ZGh3NoEWfYlDgnjX2J3ssCJdbpUmkZ75zytGrz1lTxoKrd6ncbBvN9sk0n4qvWLk9ABrFmE0
LP67tDmBt2ylWkO+QgnxCzXPg+bkexKrNWQOJ/XOvg8yqz4+rCbXR6nGdqr4B/RU12Dtt2Aq+Mhn
06mbhrM4LDWFFT9LM06MW1H+rfKKcv2uLwqBoog41qQ7SYaloa081VwIJZKGnNTddiH691Gg3Png
PLe2DPu61eXm34rGQeFeaSjTUnB+otUZuZrwSTHSvrf/3HGCbMmXOw9G4n/IclJa2/rk3b2Nowfx
oEH5ro/4TbWmWDHpmw0A92jPB38Wn3E8y0xCs+vBX+L2R/ikhX+5MtZR+ppr7psw67d7TsQcSIPr
yS4VM6T193Gyx6821r2lO9tSvAZPJXiNOESIE2oSLzxCVYkg4cfV0zHSlrVtudoQGfWeaGhAclF0
SF6AUEtbef0JVp6S14yXNtjylTXM70ZCg5wpCQncs6kbSgIFLFMEvRtDW06H5hVEZyyys9jMcWgF
hci/lO8aeJqkG3ZC1H01grqJXcWg2JhfiJSHxSGgG76PiuoSn+MbAWek2OX++btPcXycwA8fyvWG
6TPH8FZa7htvDOapgpG05OK1BZS7EMkjWZU/wInS3wTpxUCmVcaw+lslfcsX/qdFA6aUS0Ds4gup
dhFp2vUvGQx1Z7trHyrRbdb5kpYq1wNiAQyD8rQrSHAAWMJ4Tc0kQAxleZiwS304bNAjYArh2dnC
4i6cbE69tXOgzObEEcc00GcUp3gKPKgjjj/EM4qZPCejB2uGN9kBtk+RifO0b6DmDatuJ7TuUXLJ
qK9vfYwH70p5lyOtYlxBIoN9a93EfXuU9Wpakdjlc8BvBzuc1WvopCKa56zkP25pFIOC3Z9BjfMg
zMiBUSK0It6bk/olbCOcw6Z44777jlqZP1AQu8HjyDalyc/1SFSV239F6Qw3cSFOR9eEoegs+LDS
swHltCrDK00mdo8Pl3kO/hel5rbPKrS3eGq0m+RhQR1TJ9Upt5hiA87bZv7vhmMSXJGSXaM2YY6H
YU9q3I5AB5cQ9trjby7pnl0jvysHQ7mOHKsLG0Eu/yzG6tc195XZxngbZwynAweQl9LroUoe8W8L
D1gwPGEUlYZ2ZzgMlSF+mSpgWMxGUPyAnOHi6T0YNZu/CQdfwywSHh+xFq05W7BJzoiAMwUecGLz
BnWzxNw/pfo/VDJmoEeGlz9lp0y7a2ef4lsZS+avmOktmhoLihv9vJNgVOyNLOgTkzhZxZ0XekMb
VTXQ724ApZaI3gg6lsN0Cv/7+Y7uu+RUAMSsKk4ItZyVPng/wsTDOS0/uy+3CIRVFhWP0XAQC2aq
I70mM/45npqEQDtDwzdHtmFkZj9KF3mGvgjb+697JwR8UKG7r0sBvUnXmcWy5Ph8NO28CuXUAFbv
ppEMz8foq9Q1pjWNm1IroBKwdvcokXMc/8denfFArdaT66RvbsGIG8blIOop4pPP4e+7eR3kLbbm
NcCMcM5b+PHaUnaOxKst2MehIPWWd9YFtA1uaj2bn22kLX/P7cdxIHWcxYVbReqd5ZaMfgshSmp3
l1JUqKDwBGzNsWIu7uDRwXJokJzrltIGaZE3itTN3LPyuOqkmYxBgoK7orP2oJT05UtpAEebyTlo
JKmXv03/JOIVdEBkIoOY/XUArbYXSl6kvgzzXu0DmtJr5laxTXlm8ewbHaKIFFcE+bQPopCd3v7s
g887xck31KtwWFEDhZtsOLbVQJeCf3QfWUyKx7snoPMWwp72VyN9vZrrul/yGsCFisrysJcKTpXf
v3is5i7Q9WY6AaClTLxEG6fFIe7wde/IPkeg7+aCFaoB22J+oOsuj/EMH5OU+qk1bNmMO65vx53r
EVCSOZmHkpg/Mv1xoOiBrgm0pKLoSlEChnjRbWQ4S6hpw6XvS+aWM3RR4zJ/ws0+fd6GvkdWbxIj
dX7p7BAqpu8+QJo4y8p02zfciJHkZDvEWdTgO9SH4+vSvwh5MNpf0h7+eSLopxeN38Di6fw+0rEk
6lCN1GZ5szdM5ONLtcoZ8/Jne6NM/bBzPgqvZZQrGceOFSem9fLEtEi7GoD5Xr1XWowYNGiWYTwt
k6YbJheZa1mYqKVWf5j0E4nwAPHhBuUXPd0ydQdM70o1xQY8suXoP6eMYHv2bB9OMs/IP8HLwxQE
KpioKxVn+Qv9INQSFjvss1t0LGvXCUhmYGyeX3fXuqSxkb1sRDqdPH7Wf8OYJc5R7byWKICl4ZXt
hqj7WCPM687hIejnCJz3RKtQwF89PPVbkiZ7W4Y2258JcwBOFg+sLcSm/fqLWgLL68vuWXdDlotM
pijFzlA+6ufhJivKHw1FEcCj03jWjpiPyA/HuADfntzK2lNd3PvbVposYg/EfxCxntdnS/GKjuZG
K47nxKVxE9AV4v46z/ySbfW/eX36ml3U0k4F5N93VohlO+/5ixBRD16z8fQs+C3Jczka/t3mC3rI
O3VeR4zU/xlHQuf+L8gkdUy0twu+jaWl8TicKI6v4fNs1HHJA3kv9/09MNE9mdUbDKVa8KJ0TFRR
QxFjEOQoBGhRjCwCE24JhGvJNHFdOHeI5p5jQtwyhpTko+oTPxNEVZa9HlNQLSnAgujJPPOMxqLf
9S5M+t90k1F13RcBzPw2Rvjdco+3JScuMbpzOkx/7KXWqpbaWtxZldLzC0HVd4kkgr1PY67O8V7n
6XYcyDZf6TP4ds+l1gmH9O7wP4SUNWxKHh9iYqscRrZDBPH3CbEY/B8ZCp75mmrAb+l3bYgWWFnr
vnW8zV1tmT2BmcVFU89PZMY/Gfc3+kLeVXp4g6nD5soFXDErqZlI6AA7uLTwVc/Fan7R0v7KrZtb
o3cGUxYjTrJI3eiIYF2HeJoo1JVB52y0KXdbeZwJ/y/p2ofEB9tf3QSOAsCFYbxjNW1w8VXRi3eI
12XaQo+j2EuqIioYUonTElFCM8mNb2eme9yPNoZ89Znb49QwHFxPwuOW+cncdwG1abyzFe7CKMty
ayrlOzpAhokXISbFSJjru0e9cjmRMlen02MdOFktsG81j0MkWZuHA6suVKNM93e+TQjCEcrU7gtA
4iGCax6v2dGbDGsUrTUl6aF5qm9jAQVCgAKbPz2VC892QQ+bNaxm3W61xFzbuIPjN2yRsNLQA5Xj
4NNh0CQQZ1FOTaeTv6/Jjynck9zhjEDTLhq6bzknMJ3T2h7xm309/QUWFAhpx75o+++q0soI95Ch
RTI0CT9KrmydiRX6pMTw4ndTxdZP6T9VNNpAsDfJzHQ2I0vBddZR8cvzFQWAbCrZ/9uLxEa0LdUi
sneNsiejLBi5891rVd1F3U5O58o/N1haBfjnSCZ0DGr59T3TcZwPkbTZ06/RzrrxaGMMKPOWpTbn
167zcoPlqtrkI1K39fFuSoscv5ZeecOdBLJ6jZVMqWDPMPmkO8l23XMkh+ABoVLCHEd+b0rSo47Y
glY33wFbwAWs8TVQa8IV1ESH5pCHwU3zd2w1CygEWYexB2VzAsp2u+cTP+3M9m26JvLrqlyGJsRQ
znoGpRNgm3GKyhIzDTeVyw9w8tc1aG2VswDZaO3960igv7Hj8iSVrbxA1KXa4GHHaXFNkTiQaRhv
unZhHrSYCqm2anCjtSKWOsYXQs6gbcsXKoiSyoH1HXgK4Q/bGriu2FR4JTAcW191Zxg7bYd0Wnch
SK4O7EN+6FyBVDMYTwWRtqODIpiPXlVTbA3bBO8tsSvYFJyRwHevbeTfkgF6Sa2X+DZkD096SPkd
VmJa3NV7Fvi+mpfi3WpL0wpy08q1PrLo8F/uws3QW3lsM+7r+GxwJCs0KK01beWOCbF9PTsuJyAb
3FWZliHGzX8KWt7+zF9FDJKaGkQt1eYV33S/h3mXvNAfByos2WCIXJoKwZyWWA3UkLdAh9YjYCz8
Sx/uaBZHmvU0n5l4G2O0eDrADb8pSpqQVlU3pYo60hdrDy/+6C+Sz5wH1HQc/sOqr6AxpViQ+HRm
MhHN9eI/cDXexsH/zK9/fzu/KmdcRERNlYE21iWoKOLs0bQY8AQF6gwCrXRMJxyhvTPZ31IFZzm+
DubJEx5JUEfTNzrGFBFjRx4DdWgHDfXIbNLqqtj+3yGv6JAaxT8yaowToOMNrh4FZCcU0MOS/UyN
cxG0rcv4QuSYrrFwkzJSif/xQFcO5N/CvrtE7sSheKVKc00COPr5FvTxf2QcYkHqA+3a+CfruxUB
hzPprlXAW8gYKVMOdGXydIvFgcvV9eqlDSyOrEl82gX/5U56JCOzQEAfFTDhxUIpgvNVjdkkBa04
vHPPpsoI0DPo4ku5OD0gtxSZ8/WoLJ7Vn0TAhSYZkgURuljQwqSLeOfwN492ExdGNoTS4bM+UqyU
hFpvPXsT5HLvLtc+5ZsqHEfDD3hBsI9tF7/mmZPjwbu4ZBYkJz2LrX/Dm/4uN1vWWE/3STm13fkZ
a98AQWd3vJKr9/NK4GyHtEuoF9KgFZVdycMEITWh92pJWJT+luSdQGwnlbOm0KuaAIH8Muti6OMD
+DT7CZnFrmb5RbHme7A+SfzxIu1l9os/p0CPjLrG6wWyPTbL0lIkMvOzy1RzNs5+nfi/JLALNCVO
dh3sfdL/BH+2Fgy27Mj9Wa4NhJwqS8EqbkJO9dcrENkC8x4010tW4faXiFLxGUM+XvL5xhhvL+1E
tADlJQcwS5kFk8fN5l9RVmm+x9hrTd78rFexuqltLPELuJOkmBphIx6kNed3wwsYtdI8Z4vF+rK/
eS8E9Q0o7ZIPQQneWt7GaRsAybTWu8mquGYwVhQp4DhPMSoUQrkaKG8/Wzli+KwNIg7/zOPA0eyx
mVeMu56YQgtLrw8XHHjao51VNiXESBkAPfK1OknzNmfKiCR8mqFRg5+vFHgBle8bGI2SjElMl8rY
4NPgLUDGZkO8z6BEGkSM3TLjxAIDiWTHQZpmstj+5AfpDMfnurMvcHRMlXyHxNUK7DD+B+vft+F2
VdHlgZ7Ii/iGfmr7cdsbKYMAVdaoMYXHWSTkzA0BT687NTq3RDkLAAJu0W4/smNfamEYFG6Z+X39
53OpEuHa15MwEH7p/chfs7ognoiv9VaE7PyI1mNgIQnA6pTXjQSl/lWsHjiAUjEFFSLVZ+UyuQ0k
T6knjzMzVbcJqAvPYxJoBmjPCmOCF1qFQATL73pYXpGkQ1U4wX+LA0Fnw28SZdGV+es8Vg28A16n
qeQ41ULc5Mcit9QZ+SnRvsYFf/ktO6oEHFeroKKarbB1zpDGupSr8WAL0mnj632yLxNhtYVHX3d5
cI7XZydy5RXGPGr6Fe0gCcIpn0Tsr7pYnwFqws5X+Vrj84X66UIPbztYJZC8kqS2CreTvb1iElZp
Pb7CLnhJAsBbVdUwpr+lZb7i84YamSFBDPP5SmeKBi3QD5UrQQEzdi7+gt6nVTcm1BtLkGaDgE8n
Gn7FkQ4/xq7tZNu3wj0jZ1rvPSOztzEPKS4kWtE/wl8kscIv4uJpGcea+Myj1ER9RES/qiZ/oWyM
Rg67tVsKXaAwAMhwjpgvsEnNnyGDEcUh05c2Lc58aLRAuHV1ZzZUw3tUE1oLXeTPjsjt04olC1Oo
WJLcN4qFi4hpUlIwBvZ4tU5z1spiHUhd98RMb+oTUCjtBZ4Oo+cb9gduqGUkoOlK8fqqy1qalBx+
lDX+ZyCo4j04ac69bUge2rVlqVdaLEsk6v6yoBBQyBX7AeGaIwZDZKavohjqlvjtcM+gGr9H+5T4
cNkRe3o0dMOkgwQge/M0py2hnYN+bVAulxIjDkUZ08uGUKEi2hsF5TMiDhQHF40klbesoLTTYZHL
4tXKUXO2fxoytP4movytkwnIkD2t9rcq3TbaqTSkDigEdG30m1PbPVYkqv8LFOgkY9SgrLpkFeGQ
y4g/MeJ740wReeSG1pSfEy3RpbM/DByFsDksRRbntGeZzhVsg6eM9hX3OWzMWI8lETaZnUiaqq3/
xDUrAZgWNGZUceEDcSsYGxLbxZ/hFPV9m2yhwCgXKuIZcQ8vsT1jcih3drfCMKhDmN0xZaaSJeUj
0fTWspukmcwSI8qA5r/T+Ui68GkJqJQAheXjJtdMlupOiVnYJFX8PQkf5H7oku2CNugNjYM/RxMB
W/ULHrZqPhkBH3NWPF18GH4Zck5TsvZtOtfQgozeOih4d6EnABQMOeQt6zZUvz8MEEPRHtebc/jT
eUvMerijeGtRmxJLBECbstk2UTauvvUDXZwLrJARafKUdqpQa/mrr3en14ov4CNHist6XvRlMTEV
mEInCc4lkAcdM1S/tzqqesIrdmcy4KwepBU2tZTTHxOHhPfrB/6ItNLYKFJFR3AiiesPoMxYn76o
vWi6dNzbS8nV6tmjFMQYtqJIUUnDErtyNOp6FDN5+6ZJiFotz3NNOesvHBvJ485O/5iJX5926f/d
g/2HUx5b5VSmeCWnl6X0a3ArC3WDhWwzKVTzNqxa+KXq3hObfm0QMWKTx/OxLTTLspXS73puLPHY
BJ+l2hpz6RkotBYg5rPeeKLb9v/cjfH0PfBwQMm75jl6DBfo0/icfhC8HiGNPltHjvwzh1vCQd+I
GqmIiprg0yto/6nk2ZqvPqvxldEtdhiAKQhhBH3WdalaRT+JswF6ybOQRANpnG3krr+fSxytcjkI
K/yMdtSFSjWI9AJygHThB5CkKnNITuY7C55cwgQSLiS8ZBTowm7UBPci7kOqJVlZcBs8qNG6ATD5
P2MTz5sPYtFGrRB0+Umxk/IrTrPzdNGXfa4P+V3oiWVJlbqfGlMm2Ho+qqCO8wrGPzmwV4ZLUyOn
X18mk7LR7virPTCBPMWMFH0EUwp5/xB74Tl/J07wqAHgvJEB/+YZvGN0HUIfA+//MeAnamoL/pvB
HzpIgTMse3xtBRLNew07G+piBfz1hk6SsL9laeVvdYs3/FC8WPsxMgkq9wrTiye+d4OZwYuErVxk
CV2+KwHInNJqsNynl2yOPexX+cDxxRgV2+Nf/WOQQR88INGIyWIQcovtlD9YnUF3J1onv4CuyHEA
x3xBT6b5vBOdBexKex1SFeNR3OVp9uw8IZOdBrS+cioTWgpOew7hwfc3dkGSqQ84/SRiQSJirrvv
xxww5bpO0y17Pgdhk/zAcj8ZtwtrJ0kBmjsSpbKaYvCnqVZIjrXekbV7BRFLXClSQP1WKzTHbTcV
7ByU0yPhR6MwOtC3tDaKGa8lOQoDafqK5UgbGk1lGZkaOJ4t7eBMdTP1Vvm/PzHqxRmOyoEL3tpJ
lFJ2AlzF0H+8KMouyeAjllWamefH4XAYRY8eC1LuoJ2nqXDpJbFsauqzTyJTaY+sT6d7wh1K4EY6
w5QImQrYRuSJrzUMYS7dYsXvlExBU8gEaLVO6+ZWXwk2mqhwPfFIXjVuHKBC9RozCGalMRXE5dtN
SsLsXs9EgIsSrTuTmT1gFsLETTBRB2S3XGpvZkTgReMlCXe+j+IBiF+FX+7kcroJekPt9nSt6Qmi
sI0MnONvAIFIPzUeTcpj6JIfFIFOmfNxsUe0cyaicGeRi+ASsrfi5AoKkVueh/ZAxdBDucTiWzqg
LuhCXggGTXps7EAck0mScHR7xxrCDiEwi8KqKUbioP+p6fwRFNgBtVEarccOcPXSp7nIqqeF3ybH
hTvMYtYBdPRGXVk1b4rQjABx3f/hLUJ4iAQlusHoblOXYffrHuECKxe9NtW14ig113IgFpN5tuU0
JB2RcPyzNutS2mQJLyRVzUNvi38VkJgkzJ8apfY2Dru7y7lKdGyRmYapDUmD26VJpg/LvqCxwfP7
yIINHJoS5Qsx61TRYtm4YDIEKry0gQWhVtnUDtpOpNJWlpcxJoZdhr3jAdbtoD66dhccthBQjLoZ
nOIxpbfGdXLntmN/ExpIfhUZ0FXiI7FuhW7XiXfV8CRGsSSEkE+3ZhYAGdxhKyt+e3xOcY4wWApo
8LdUjm+WaSu5OJRfJy+Ya3IDPvctcSpMFV773Trs4Bp2BW50Tn1obInFcAWZIjTeiCmiPh70LJpM
gKVViAuuoJRFoutlEJXGw90DFJFhzFmFPX3wYzRYb9bnnCTcXWzXyAcjR1uwbLDQb9eLEPZi2S/c
TPY3lLOEboapf3zMWml5u5Bv7fc3RzRe21vSZStWBsKG5+ehAt/qHVms3up7sl3h10ZDu6+uYKLK
j/WULuIz2y8iAZV1Ov/OIrKOlurK6bJKklIYZ1HAJ2kJuyuB5kSJuODwbz/l2WGMlRKY287SJJH8
8PmHjaf1IP56ohgrWGBz30wRnGOmewNDoqSfatbkvSDn/D9Gx+buP7fD2j5UwYhSh0dpa3n1YuL0
lwXlcOni7hx3y2GvUQyFn5UPvseV+EmfdaHmbJigNc2UQMbeFPO38DuTmu7zs7OoY8sDAUS9GePd
CxyJJ9+pG4rMhXE6EAkrBJ9VNDsTXHmetJBEk7nglBpRUOGco1FVkboarpviIwI3jkcfruJTk+Ho
nCWANDMSv0QClFGKsA4WnAWDTO9ZiSph9v5YfX0u1I+uikeMdXO5EGidrc4lDWOtqEkxAKaKtVbu
9kn8dBojU87koysj/8ijFy4UIIc4EhdM9cUPtN0bxDwhT3K3vB5v+7UsI37/9pXs2F+KwjFNgxUv
lHnavNTCAIsIXkhHHPgSKetzpfTQZF7NseH1VIgvvTftUp47JiiFxInod0KdNjWsSp9NzAd9Yhmt
Mqgi2nWP3KqWlhAQAhBY3BcnpDJBVm5bpvpkqm1LrVWnFHccdmXSm+lpY/uXG8u1GxXXxN+XtErb
vxnQ0OtGem9qpDhQCfGZAY8W87SUXuFaUDlSMvrDqPVgHoTnoXScQ0KYC0xa5+4cdEH9faftPp9E
+l6M4ZARexAP1l+RLwBmJ8bQlieLZEMjUkXBKpFzssGzvCsSPjeGHW3uXdt4BZF6TjS0+PAeTVEy
cQ/5OOcFswWvMNhWluViSyK6GU+o0lbS/TONWp98Feg1SnFjNvulZWnZzOcBEWWS4FZZ/pxv3Vmo
oz6Iv9Q20f6kAQ3+8nL20pBew9GJYUgqLozIz1+7OoC6tOeCud3UflbpEn4ht0hEek770ZW4/QUQ
JdXXkNOKkv/EyOOW+npuAcnrheKwDn+F4ba7+21fFFJ/9p2qM0AhZfBKQx4ygvlnzvBAEa37d5H/
LDifir3rmSv4L8OOWmcaxsP/kI8mL3sAGPieWwbPxsfLSiMsannhlJrNS2mk/Qu1t1U7IEsLD1EQ
PmHGJWByfCq/xH5fWpT14Pa5lmpN2zxqjGEF2Pdyk1n5TLn5lAAklmaB1CXdWaMz8rwSzI7gHUNN
GW2wuzj+LTh/51QTsp/bekA9eR3nkDBK8Pejfvxv4yDlauHtFuqfIQ0mC3x8NT1MFc4rGEU1RTvM
WhzxTx5DUxRi7xWRCSkuZYQbfvTXTMtfE+/kXDiUET56zeGe0dcbv7q5s1oFMKBcwvJFX/S1cqpO
x7KzcYnLlPjn80loSz3Cy+S8GE9q8MpGweBZZOWfK9eBaIDj5WftEt0kFYfd6W93du3UOMk307hE
bT/rItprWlbz2fBLPre3ZyNNmVQLtqelz1DNc1yTdN4pOrPD2Kko1PM14o1VAYvgJzOl+ScsHqb1
Ux+DERrC0s1Q34J1b0fXGAjrYPhiqwppsjzPhgmGODU+B5vn3yUrlMPikia4vd9tM4vYhjXN05Hr
jYiIx7mnUEF8fh6DxpHhr0UPxgeGqAgsFEpMI8dkRqvAmnfo3zn97SRa49X3toaoW0NlWnBD2kyG
jVsZQIeQDJqll1s+hR9XpSqXuXru2eEZ0vA+TUhZEUI/BQV79b+ZIlXotxpu5IzH1FmbnHRWzIHy
zYjF5wYDpKfQ6jxBs0Cahab8UYFdZWkCR3UIMKjeIuHtTT7FyvLEFLaIxoBjNAhO2066TZT6VAI+
pxKUmXv3+AvRucZJNvE+0Q7KeXLBRsUO/Ce37nZ4sKqx5+kq4j7ielLUGkben4Sh8dLyH8L5XTWY
yOSv8pxmT8svkUt99uJyrOMk/LGYBdMH4r1ODFwoN7TOhadtE5l/RPRMIndZMiDcEacZ2pEg259O
VDTxg5W2pJpBPUsaYK6fMS2Ji2QD1jTFk+toZJacCmMGQvlMi0ZmWZ07wYhdm1CpM4UyLVKqhGmB
Xc6aDUeChiafYh7yY++w7ZEh6t5wSFwmzwvC+ZzLWWcEd8tV1HqKh0Bp6cpbZDqbyhGaY/t3AlMt
1lXtCAq6MjzGY62q2V0WT/9BC2m1HHDzGN8LvNH9N+KG4ccvWlFDw0gAI9PS6MSLDWltXe41LltL
RPaAwiGK0QkQ00j/VY8rDq+BzUFN+fmmVFko7CzaPGKS2PzfTi3o7oClYb+sYSl+JPBudUcUhypT
EVGk0QXRL7gqI2WmwcR6zMHhrVZAYGipxe6pdHBbeOn+T+MdogaVALQg9EpL0ttotaiRZqOYLB3M
TcCMiqOPt+QpwWwkF993ZUpbPz4Q0kASwwVJCKh8Zr0lH/pkGq9644MuJrhG4txEokeRWoVW+3Qm
/icPSUqecf/66GGfYifHczcLvgUju1V4QV6ZLBw0HVKn7k/p9w6yOvW0Z+OWm0BXvxp7DoaXXvHv
7GmQsrmK5PTwDkVafO6ZR+jomI4xzTV3pH4YclMibQVw6Ldeph+p1I6pCicfIEw0Y3lvYWif5Xtc
mioaU8xrvEYa/Sy4nxDDBUx9hIaShtVlFAdeXOHYwANvm1HU3CJ3z2lsf75mqbyC4/btFjE/RQxN
UJYQ8CisEfI9gotDOs9cQHnl1v+ptnp+lglvoVVe7QEOvztux1sa13VQ4WGabCAH3XH9fdlE4mTT
Bt2oSxVH4OqOAO3OJ7zzIH6SylzTMDUB6ql9XRJZUbbda1hoSSLWl75Y4jV1Vb5VwFS7bY8oSA8I
4mpCdPd7dHDEKn8NsvzvZVS3VqMW8AZ2sZEuALP0BmzOnrvc9rywFpPo3g8w/Ap3L5YT2dc4BN1N
Wp1TJNOYpwpJKBxIIMtqE/m46Z2fRIF8EMh+7cQIGzpjudmgl8yDEfLQkQc1UYYemXMm9pVJGWv4
law+QKu+a0iXAcQuNhjReJWFW88GhUg9j3Ry7OPMTEKKbpjH9L7keaZYl48A2hNqUmZBXUSQ7dFV
YIoOSAlLGMiGjH+W+BJClMyTSDBdNkYYFGKRxksioan4xsA8tSiEW6PMpVNERcfATA1YEVP4ppJV
aDbOO4yjzo2OuyqaBKHzwkDvAP7wQQdf4K9AWKsk05qYXstIFFQfawx2bf1eNmR5IzsgzfLD/0uH
hOfvs9mPuVstRR/A3WOH3bPKbUoePmDLeCO8U4z8s8b7xcppcXRk4iagAc+7u/G53eRXH6RgsAYM
dKboX8rc76K1Cy2TDzMALG5C7ImB1u/wnb/bb/QWZbNtfX9eMa20QdZVkqIhsgWDDttFeep1DiXW
d4vgxROY49PLyqhXALtJb16VY4AXVomFRtAsllRgpLAbaocDj9AJIwvBwEx0JuRSF9uI6jyaO5Jj
2hiiWWTnx8wCsSvyCcf1MijZVWfpJtw0W0jjOYfqhRX4hvORKf0M4yH5y3tx/8P2ydpmjr2phc+P
O4Q0Dj7cc2bUsPal9aag1yXI2lHOpm0hlnrkwtJrvbZVVJ03nQM8MoE8s3x+JdGmKy7yvvMFh+QU
vNaTgWynwYj4O0a/IvMtjW+RX5H1JmB7bG7X0EiAuCVFFV95f+bB7ielQ0XLlI+W8urmw4m1FPzW
gmdsuEdLTAx4zwjlr7UBBHP25QBbyBs8hgDynxCsv5x/tAqBlhhfZ7UC2vRUANxweZlkMh5eCRFB
Bw+3jliAgppAKmG51lmUujdeo5gagTAvR4YQx4e+iAzUcX5i1tIbbITPbOfCi37YY5h3/6E2r60T
q8U4st4ofa2SrnB66oFCGVCqp0a06q/m3LNsJ/q93SdjVcgwRn4eRsqlCg38/tup/KVQSEfBpqgr
aILpymm8cHBb4gfv7WbbyYxbcRxhOqZVi7hN3qxP894TBq4x8hk1bLqy7Tuic77Ktz+467jGnk6F
lCssZAnQDXReaRabFrPAqoQOO3oiemTEaAxuht5gXoMEb0LkszCNjwbGExC0cfRmV7Xb4dsEXC97
IaLNzgYxaVZraw7Za9eJ93TLgImCTRrXl6RTPNoipAd7R7LHVqJPVm8A4H4YqRSYeqhg1pzwraen
ZK4p0qUrwp85ypMV2L/t8Y7gYpGMjWUOA2yr4c3Qa/oC/qiF/MQV5orcJZWpcPiD0JTDR5k7wXUE
kwUn4Cw9L7HeCTr/+6+1ClQm0nah0Wg1N+8UOxd6Fpn0qM+GRfeWAtduygtSOObdYlkYMNyfP7AU
04NsTUEiIjqCmKx0lAdSsny/rFoVkd5BBOk2rsojjHC9/6wyLjRfUmqPJgyeOOl0eUYWT4Gp3EmR
jCwBB5o1UtBRgwMMrB68fmuSXsUIudLL/93p9PXDIT0fz2QBSMmAM5Vo/zT6/ENoWwRzVdWLAnPA
7jYzpoIvh/2/rh/m+dwXfwIc/7UQgXpkh8LUEu+c6WaMSSLf+a8WpqN4wyqrgizMHNirJSyZ1D80
or3gzOhnazQbaVGsePkamT/tIKtoeDcha10bBwn0mb+psY/97UFvr5eCa2rDLu0oTAIOqXAj2kg2
1dlk8MkjbKgWYz4yG4h187hZlYw2d48gjNkgxcuxPTSaiq4XjksTICDQyWXU5HNpru1GgvYmPtKC
ECAy6iHoqZXaaPkf4JYJdBqTClZH/lgnNf4h44VE2bKvnokU2cXGYRSQRzye2XHR88466nNd//MK
yaenbiit4gLM3K6638feXqD/K7j3QeAZa30OS2IuS7Nmwhn47gNLPL4r4G5wumF92rgfv+MMgvZ5
jQXKpsCGSIgsotNBIynlSTL+hdktFN57xhE//EhhYkAF8P7xjTzoGesEWhplGaJQ0pBxalcqln+G
fIY//BsOGM8L857SDEQe0/eFXzO76QzAVmpmpQE9tgrTORjKQcnd4HNajjB+6VJbrQCfJjgu1Vme
68Q/aMlTMPmHCuWWEw/wZYqJDiFlsoeKz3+s/4RE8V6Hvh6hZW5cj0bjCDcyEibmLdzzMvvNR2lH
qZvsV3yOmf8Kg22/DYDimk1147L6YUkrP15WAvubVbezAfvjw7H1pfJQSuV0E5GGTH6s+gDOzeRf
HUF7bCClxvaNO1bMaOrIl8cci+ujx9WFMp/JUemafezYtCFt3fsMaLa5wZ4LDEQYsM51A74ptURY
UsQDbyVKsNeV2cFL2hgyUMwqCZ79J4U69sc4jVVnGgaIohc/S2ZJA0MeC4RAHp+tikzoR70UgTYS
ugIqYWiDMcw256o6ItBGa1NmROnBHdMz9Xqu6hxFv9QZw19Q3xaME6fFdSm5QydHLwHNTkdGcInG
jV2cctzivpIESRcF0rk8CFTptpKXIyWQhJLc2BOxvPd6bo5F8rCH3NmTHXPPKowfORgTi2kwiRux
xd+Rv8NlAaV+MTyaNOg9BuCh0BFWrL3HXzVWDHlTshfXNczAPz12t7YQQhLWvPnz8rZ1goH2DBfY
jwQ8dHgZlO6rB+qwWGVUm+ZmlXw4uT0wV3MzJBoneahUIN24CwhTGCrvrb9gCo7Am4IQB0wLfHAQ
UkWL5niscHQV99djOIZYr4K2Rzq/nSY2ENPaMsRRyPtsBTH0Fc9CwU3RO+OYKQ1WbRZX7FiIIN6i
s30w4rTiwnFtJTlHlahrPBnamhhuVYi4A2bTvXUKQVYFXSi0c3c5yvu/sGgbzleDLF9VgdvKwsdA
2i7bUB5bEjxyG6Dq66VI4OPL3USAdU5ybLFr9hO/FG4fEjOyRb08UBWc0SfoLhBdoFKZ8H7PXwSe
eFNuT0+OOp0fpXQdTZSGHyinbMt9Sn/KzCUqJgM/AXetOhfa7/SliLBf7CihyFHlejwOe/Twee5O
AzmfNCO4uNspaTTWemoG5tO9zv6iptN1++Dm8X5R22aciRzeDpY3kPrwbLILOqVRWXIItjttBzsI
9aMdRd7ZHP/BLuPLzKDupovNYzum0iA1gCldpGesOft9Rzed5df9CB5qMLGu8bIdItm7fMYOJqTa
KxXOj9kr5cT7usqsnWiDseBuMbOAvUOAqu1ug4eQ/XpE2DV0FIMwO3YHaW4rIBrMm3ODUHQ/elal
CK5hWtBFW/j28lq5DZOY8eJWvpEbtnA9bI3bnyVHgLU0IoxrxBDdI0VoUbZ3JDQr3pcnniT1aubE
f6THDWKegmRZJ5+eIhL1lgNkofGXI+U9rSuY8KdqhLI28IqESkK+DYUdigVFfVdL0rnlELB873/z
iN9DrjdC52IygoNWj8yfXJ0eZOjYbs4mqe1/jSqMzu8pdL5gTtEK46PhEVPyZ5l3VNSIG8Q4zO7E
8UJgvn6YH0lv7DmrTRt3v1yb5Ktfwg9DWx/AVeKNV2BznU/TKQr+poxrhd0loe09jVsE4xpvY2I5
idbn4vfelShlooVT6u0Ivly8gXteDgSpFquX79OWrJb2KoW+7ZWMm+xdpaIMa9KwistFbCxxlCO9
lbcWom5O/f7h+aucYQOEI9qQcXrWpD9FLc62k+RqyVP9W+1r0vNxf1dO4iin0wxk7YDZJ8nBfaE5
o4vg3JUsAnPlc1lWIWB9cmqA87qs34cWZjJvlVhcPWL+JABZcb9jPGkB0cWNkYq0K6NPY5TKTOPI
/jHp0vRE9SzN0CKko+n9J21k7HJg+DqfCAoW6qM7jLe+bJoWu2sK48Z1YGnmAivORsfyZYzNQ3tj
/0+NM8klGkNFOQU909+eHSOyRP9xWuEeEfzn1kYuleNHnaHcf9VGcItoZ4AnXB80ZJQrTBgxynbm
d7Jhwb0+IX+F9OW51dnkozGxdhUR6sIKCzh4Zr4CzGye4ijmhsdsp81sVCe5mgOLsSs0YkfEIbAj
WrDWAFJDd6IG+WxApxG/TrUZLgl/Vi2yFiN2DpuhAEqsTW8HJiQUxLCDD8ofmgqM+c4TNfqDt6H8
T7nkUFu9CLFGVT/duXs5dFObMGGiwJ5YxeR0JIWd5ewvdRHB5IL9S6bBECCacO2XdYHPJ0O8ARKA
GHSbpU1dVEw+wqBC/1hVeHTkjYYkkWhJEVCudYqFNV7Z0cDv9FGcYfBI9CkD1ZEqJi8ONgMvCaqN
6tblOHZzZovEhML80IrABZ/aPANifbq8Cn6+K6zIaanmYsHJEePH695GDd6z189SFUleHvNmvrnS
QVVC0iVAC+LfSjAjGm0mjtJDxzNtNvqoE4G2lHvgYruwDsH474r7qOiH5D9Ks48XNjMPH5cz21nY
WscSWYqXY7KI1OgXA93O1VXnO3gg2b9+mK6K22C212cVOQ5YZtY9E/Rvgpdd6BsZeFaf9ZNAKNGK
q4N4LFk9ZFi3QVkHr1o8qed6Sifg2L1N15zNwdRaHH8R3+LoYhh48YOE90snZVRF8K4j14qYxaDG
aEvWyMzaavOZfAzq6G/a+3wZlGrkkJwQGssSLw53Lb13MZ82x7B5v8AwvXJjxnNt3rxcOi1ZDPVh
TEDTzPIMVz1/teV4vMcoGuT10usguVPm9Ccuv8x5Nivx2BqVxjKcgecWFfatwjSWwhKcVzvIxhKE
pXG/eEeoBEsnXOD1VmBiBVplr+99VZBfAzWMmesdnH+JkB98lr/CmDcUspfUMgWrvlOz1mu06XLo
UIWSWmuPdnlasMQZvxejdGAJAUO02mrO6NFCg/0ckzw8TPOPyb2RtsZ+Irq0251pI3kjqMYylsiK
0hMFz32nDpII8JDNGPqOxY4Lj62denjnlMSz/rD6agWP0/6aQzr+wiNpJhwVVq2Hswa3+DwWmXmK
ML3VBmFSmi6vk4+S/YCRvHEFQIBlr4dmyJiA/HAgtH9okBaqPT6L67Kb1lCqryyNkcm86Lo5eyI+
iOq7QNM+HNpThrOkTMh0RhJFK/wWnK18TMgEeN/6shS7r+bbO/CBt4RLz58SPZG2MIxf6Am0LLzB
Ewty74pK0nMmyFk4UvWgX/WG6ZNtXWn94q5IVmK0VWFNlzIbJvj52DB01ZgkIo5GvFyeCvdtgt6T
SzMeSOymnLxDH13mkAS7rp/e+TuSTZQXRFz5KjUYCU9skswX4RB7/Mhi69q4Ex3dy1tPBJNwJmbn
rc88Fo4I/tsU9oqvSJL/2ff1OEgbTw76nTZr0mqSPLd6WCKTnN5caPSpuTTah5VZcYuZezRei1QR
YlvKU8gFKzKpituWz6ayeeSQ/oo7k0khpgmhTDPNng8OuPPKkqkGy+FQB8ZYs73USuGffq0VgZa3
ZmEuRGqp3UE2rd9OjgPsniNK+Taez4wgCvOeDuAtx+z1wLzX1aUiJ5ggebjv0UoGBScnmE0ZNZCu
p7iW4clkfNfu77Y+yBfgrWgUT35+ePQ20zBfB1BUm7cXEn+SJKUtJWtBmr2uOwRfznaZ28CdWqGa
fzLRdzhw59VqKfWxLv/oepGgGt86FafZgA9pJ2YK5nb092y9iNYYObY4fjNH0Iyj9TSjxkiQX2Zz
E7/xGe+9CpAb3Kch5qOTURIqya9rXN0ls1wCtEFDW1IaGLROFl8CHzLV0LTpfrV0ZlhabUdOhFji
9E+1HiIF/HBla9+HndXqcKooLR9aBQ0Py7GVrMU2SVuMf5/xGfd8/dLnLL5hhGNkiFjzCxDn7wBo
LTbU9UaS5ma+cZT+wA9Zs0rKjrvs5KwwJZJ1J6Z8UFK9XK+hps+6pNhv6VFf7PFN5pqqnVzapFzj
o3ULrkV6mbKoszJsflfhAK+8ieSuhby2dvPkpZzZyu2YTcuL+4Hh8ZP4PI1OSZRtDQ4JnuAAI+zA
x1dq6HJD8SR6SqCNPjL6Ufm0OT+jOnuuKpJnBl1DJNutYIA1YdZWYty9sefUxn3zvhecMbDlKsYB
ysZLecYGIHDC7VKgsrOwh0EHsiGy+EmqbzAqTGSnGIF7jSpgqhsUhoQxEp9tZAaeBUMHnoAT9H2r
KuizVIecqQMFEIBiOm5xhR8SWcTFNm0Ajppeuf+uykWmn14aloukEBPETGzvQ5+rXWk3VimFFWu0
2lZ94Zcm6ZDre7l338YjgI4DQXaJSbncStnFNXz3agGg88ijDc/nR8qvnJ6rQCGs86u4EJy51Z8V
ZiBxUE89SyhK9Y7nC6mxet1ME9dDw3UGm+BK80uQ67tLG4bcvnWV3On2UI6aWDoE55cHdUdPF8LY
NGqc9KKRKLYkdALtq4VbKMO29wNDmmo3q+zUJXf4Wq/lub/37aXlBpUfolrJPVov0Y+CAd6wa616
9SagdrBMsrt/2h6okeZOuThF0qNpOhDPHNHXPDd6bhXm/pvXJ2c19o+/TX2jbWViZdRPoFT0cKZL
7jAZEFenFKgA6jnBqGS54K+Oi9zWSXSY7tATWuOJ7uPOgkBJF88ovAJ1IqpbB23g3aowiGa7ncGQ
Slmhsm64ozxHYha3a8YOf8gmFa409v5P7XW3n1/TN5sH0THOsNTKtaKJvQQkPE4kJPzBNmmI2vtU
Ba7xWqC4GwdhRi1+BjjN0VQB+tzJ60RM1ElIllAjUUIRKFyykuf/WZlJtpCElo104DY0tIky5Qha
DpZ+8l5X+c4MunXFo3BWlDI+Y/SDhaslWiACs52Udid2d+btPlSvwP/Ac6gLIG6mMy69Jbk6gz48
3dJrUzO0g4KHqXX1fdH2IfsBod0av/AJk/Xrdfuf2xndQtHL834GlKH3N3hqP98OxuSqF/S0I2yz
rFQDpyO/yqcyDmJmwAm/o3GjIEsHn4C+g2foN2nwcZL1zXx4DsJpnzBPlE4UWCc7Qwvli5Hh/VeR
Oq09lltIJmCp+cR859pK6THSuZd3PctsO1OqD6WJTR+H73/OIIcyxgViW8SnGTGalehL+7UIFLkx
QBZBGpwop6Z+LLmV2v7Kb2OpPd21nwfH246b8BGC2vOnXBvM5alUb1zypF66xnf4E4r5xcrUNGgl
b3vAR8rJsNs2l6JY+d+LfRtJNF1y8szo8KyXCdlhWQkBspaCYzm2+wuYnbY9sBOL1iAzBWy4C5oG
4i3ANMYdoALsCintXLi6H1a1ZAUEzyzokxRdr/68Yb4Ya1sTw9OUBshAUhal2MmE0zvpupzoUa6W
5bP22/9gVZgRZEpn2Q7PXFna09se8XZuj87zSlNhV1Q/is4z6JX9a0VIM8xi1ptR1hCO9xqdSqzV
VCyzkOt3pBTmjyL/A+h9ipHQ6WYQkVUYHbPReavlEeobDzKmMI0yqTcNRbhMXUIA51Z03XbEhvNP
Dsbat9o7EVaF+f6KDbZIAEX1C2KKpS7cGKrng2wT7WlcT3pA7QqpjKZXMkRjW8q49TZQOyWPkGve
rlPyiw5wAuZ4MlKeegzq2X7uXYK2Qcu7aBbpm7jiHJfUx5LQIhSFIRyMs6rEZ3Dsfbr+snQKIPSS
od6iPtYwZgeW7zpgFHyncAVfXyN1rFBELVHlfMVY/qUDuF2XjZZmGqTkzXQAdgIS3ofwQWcMLPpZ
zIF43PqiJgJ5Mu0bRoVYbpjvxjKs2SKZOQJ8mpAlMzbotCNUqj8AyRuBoBMJaZZky+PtPIvvTXNB
coCO1q6ahe7Oq3vD/ulTusQ/CAxH1ZY+TU6A+gZibdpGq1Q8vAQ8XCSxW9mOPqsXEm471KeQsvql
7uLnDscpEDUzDGtVgUrTii8dO2zYHhgXFHWOor4ZG6/mpR2WLClAnO7MTF7zMGQXT5yO2BOJ6+Rv
48jZF6X6uEY53Rptsnoq5g3Y9D783XVUPfGnUz/JqEJOV2f7rnai7Gkf6vD03eWCDzAjXTl6aNlT
LsktArPEFVcHIH7SnikitiGWgiVSIiwFcXUKsEu5BnSH+Neik1r7KhtvYr9lLts2kbEKjujgTGp3
ZGYNjN56enEpBDHUYdsUnQZ0ARdin8XJZCOhqQZeNiVXTHhkg+NllMcqwCsBtw5CaZzlPIKqpxaC
7GdPDTaSOizRkAU9r9L8RzZH5W9EeG7uo7Cy7737YruJ5tNEOOc8ovLHom4QGZw3ARpZSgTemEkX
9V3zUIRiiiBiOFC/Y+lEKOBpmw5pmhprHs8y/F/Kk4PtaTFtlvwfQdPShlFyjaR1yxHu4WExKVBt
05R85/83KwUIZSxIUyvcRuVOZfZ3O4xdq61YPQcN0KF4ZBkM+oAhOtZARkS7eSYGQ70wY4eF+Eh3
4no2FFAVLV5z366bh/Q1azr7wvPNAwlAL9N5EvEdSsNz64pPzN6SsXSYHYu+yA/diQVc11Rw+wdQ
S+b978o77rKXPprGIjB6Y90Ovgd0qa7LUoBxAbr4xno+zJqL90NXi/vTHGuUM7zYd7CaIGCvs0qr
lckOJ/C/GCh+dqbfvBf8uwijxX9OQtaptI5ZssBXpeoqQQRCQyBTgLa7RqblorE0reQjtX6uyhp6
VaBS4AYtvhZSBMq/2SzEMJ8o13WDj7AWqKxn+8D52qBR6ALh9ZIpbAg+OwLhvXaCwgc5puqRsHKt
sYfbpqudsbCjflZep7ndxu9Jws/oRSOMa86R8sJKm/e6s9TKPZ7S8B/XUkApFuuf+zCBOjY+v39p
4lt01+kFVr/tS0h6TSzypaQ1Val7Sxhp7wXqaLbqRtPwkHZK60fCM5TX4+Mx8H440W3MmehQclFl
GHyy4k2LCnjDT8M/3+ELVUCRuSVO1hzc4bU/MMwsxdAoQHGpzvjhX5WkZAizLYJFRJJ8HAQ998BA
mKgRDvf16GIrNvfeQVd0hBeIddPMokAWifZ2gvzF80V/1W7ys4XTYq3Vi4HubAZiqaYzZgPX75Fg
KYZy9Yp9wKAJIGGFWZVARcfV3n+6U8feZNC9xsPYO1+LWk9pVeU1gST/K0PrMVJe+UfNzENkyW0S
LHGm1qaQT2Qs1uygfsaUIK0KSubGUW2bhGnjzCUvLjk6VXSGBmUqCJGrozNmyaFkch1Fcxve4r/1
+NzDSkNWoSUyTjzE3LMGRU9UhYES8XErkO5V/AkUrYBGjj8vMMWXbg3ym51gZ84j6DRW2fPmVYgi
gCwxaIxyDMJePxkl+8EzaB1b20tRSQp5KBa5muUrqgy0jg3vQDdGHPNkKJkdawcMR+3cU59GapYR
elM002Rah09YakSQ9Vm7K3JPwZnhPLUolz9KYv53MgXcq/yuvhMKlyvVPDozzaUMUNDggEUq4OsR
jwVrYJvv1ysaJTfWABd18CUkxPoAJyvpjfx/UjgenYr8S1rlCDB0uxUV8WK+RlLuJrCoSDgQvB2k
yUwx72rOLOVlIBy1myPMrF5VckeAUkTqnxMYSW62ub+/FREiZ049WAnxCL9Dzd4GNdWwSS2pA6ct
MKVyA/WkQQDGZNm3tJAed/YNNScdClmvuQbu1dDYZ4Ecz4nSbBn3vIec4e+8DZpXaAGb4vR/EWcs
ZluwAY2kG6lNjwigppds7gqnILk7TmysB1miBlH8YuQcc+zuz1C7/qYtqp7dyfimO9QsHRSjlwC7
YezmGUb+WOQMey+zrEfFv0NPrtRBD5DNmnfncqE88OB0d/6sCpDsfdbrb3lr2OKO+ALd1aOtugNV
50Tc44S3V8fdiYfV4Piu1monRExR6c583fJlQBuD9kJur9EA8sTaYe4q37JcVhXvSMYzZU+isIK3
vRI6Z7TihlhqLWbuUDGrzK+k5mMSTT+YV1Vit9q5K2FXMqJGgH0urjIAFT5eTS9slEY2dAa5xSJs
2NvVl9XzC+UQ6mmhCQWu4KrDcysTg1KtXFM2L+XvlkyQRHy/feJMxPzQq+eVscnSPBpHTxTi8Itl
5rhoBY29TRiUaLzJTZhwUnC5mgoV4DudYPYlIpCrex2ltmfN9lcp4CBRMYO+NC375IB81AFdjSkw
kJaGTQnEosXVmlzTmiodubVGIQWK3FqEYGmFm3CqQB68DMSSjdIM5tWITVtEbzSPW4iYtl01iatK
VktkOvXX/H3YQ05VY2CWRUKZwQcI7gAazDMSgisymKiHp28MZORkqzHXtju5CYTYXZffrhUNLN4t
uSWGJB+7GaQ7n3rqMUTa3D/RilmAhpTKO2WqMJp6iGK1d7e190NmGLugYcQS69U+T3/xHwmjjkFd
h+KXGrAJa8wT7SDLJWVgDS4ZLdB0VHH9801/Te+6VMnLe4+7oUSZMCCzLbpEtTXE/H9lmlBRF8xg
v8OEdKZXIp62CWlDXrSTEE/1GOKD6DEEvjqXVMB8hSkmgukGXFMbJora/zCRoOTTPQmxiaT1yyRd
hMa+ANoPM3ebiKVDkYAsU4YtvWlVYx2HPTw/mqps1DpsT5XnQ6kXaaIT8EhJG835WgwwKHsAlXhN
4+eeJWe5MYN6Ob9uPugCqmSOiQ67rLpocFezb76fxMh5KwRxxtAKS9YV7gGvvh8vjRDQwYf5kNQR
KCn2tnVmmXKVTc0/Dsum5Kft+CAiLR9Xip6x3C2KRlnmKImA9kKDSpRxI5uAZmMZDzchvB7Uo4EH
ge+PMVLqf0A87OwPV7JYZTRVWoAavMUQ9+Y99JpHzLcJ8Ege8V1nndXS4DHiz3eNK3Z1aFwSXn9J
huXJfRLNSg0DB+m+rqyNWpEH3BM/DRtsFCVdcpaFMOwDDKAkXC8IQzyioQaYNSivHfuyxvwZSBJ8
eAP358BneHv8113X24emD4+nRc0h3BLtPqj0yD7I/93/kBVozQEYL0EZFysIyJJvdqKvH2PDv7dI
yqpaHV/ghKX5VfjD+pDODeqPTa4HQsPwYLDJqfLzY8vrajJ72tPm2O3ahJmv8hxMLA0rrzn1HMHd
nIC3js5Igs3diNI4KOd7QMsD18FtdCmQ9BCoAkRENwPB7puHKsuc+Ddx39TvD8+iBl8ZlqG0vwyd
73HX32GGDTbLLincN3xOP7fqzwauaenNzGgTfpP6Ra8wmik9UuGcFGYo0zHY7f6z6NbNNQ50/9+C
G2B624cA5YLABJxTqjheadDcPc6Ee9WeUUbQ1Vehqdyf0jA+EYJf8XFAXaTdF4GjEb9AgbhoH93Y
SpVxvsxN7A/D0puOYXV7ekjZspU/VvGR598sO7v2ADXOPKaqa8REr9pm8Q/sz+oqgEn3DDohRibd
IONgLbiPC/fGJbM6UNIv0EQJfZkJlc81j9dbFEMTYQREJLaYy4BLfIiGqK0EEXJ98/RovlJ3RjF5
C6a/myIvIEQC2HNDQEKuUoYSJS/K+CgtXV0B1uKnAPbc5e5P0riXRExzb//zGF2/Jsp0CEyNw8N2
omU1sKj+wb18pFDlnruXrFhfEhJs6EXBMibQfM+hdqR6itM8rdo1iHdGbbFOtUD3ZQwZg4LuMFfx
JDX7GRUKLf5pPx7sbO0NHWO1wzKX1sYX88lrdxWVKP5v2osfBQRnLEOq6nidGwwEe88+c+wbLq7d
rYcbPR9QY9WdPWiRczE/GJk3q0QPXu1e4EUt0GR/+2q0d2Y1GXlBdvJAF4cn8H2r+rBgREILHKyM
5C0n3fb/QzaI7b2FF/4/OKYpNSL960+geE0RrIeMyFYCV2NJPnGvyfik7eS8cbPq5jFKHsNeJjm6
fQQWO5sqimVqo6VopYLBIcWRc2WEKOOdm6sWRaNQ5vLbfkHKkt5j5YqU90Zub0nxqswi/rRuerYR
OePwxPEZ3weuupiDlgF+Qx9PSbrT+V7xuKAx60pyDGpAdxwv/KAGG/HL1nzcFYoeq36my97WpSSZ
O+QezXTYLECd3qp5MC0M+8Z6hMd2JKuRWu3yDEjJxA+BAE+ZxBuit5jS1Cta7TJab6F7taaIy/jy
oRHosSNB9Hv/mtlEjdsKTYTpphEU2VZx5ivPpCKf2Ht+IaBWPZKk3Njk+TrPkBZ4OyIU2pEGtjtr
JYHw9jF40nfN0Khhwtsj757yB1nKHgEbXaR5cEil8dSntbGYeYHNM3ATzuByas0EKHUATNVPpcca
Un0V4hicCSzAs6cKzHX5yEzVAYn/hFlPqyj2CUPc1VFJK6yl3NW17McNrc0mwrmXs7xMWksgZvOL
Jy02gSM3QG/TRpgnm5ZsbuEoJpeaq0n7VRnwOVkNhOSqmE/aqHLHt8XQfJFLJrJHVDvQXf82y+mg
d+7T7fMNNz0OwRgZfUMCMQOvqUuiSk84hLCE6y/vRD47gfuwD802oWREyGnU2QPrcZc+hUNvQTIL
chx8pBu5KWPW+ccM19guAX3mkQ+0rRG1sXBE+vvownY+gmYeW+JX/O2hagU7raSSfgZGFy5qlRd3
H48J/NGlsSU7XPLRqWn7nNJwyTxBkgLJV786ZyEgbiyxCIadkG4b0JtM3aPKJzRpDlPvlQYfXqdW
/w8muEVbUrb+CcS9lrVqn1pzVhAGsKs4reklphwfYcwX0UKm93BrlGh8BpF6Q9kndssxljw+ej9I
fkOiVJm4ALnI5I3qVf1hS6apxS6vZtk0NQCfl6lROY/kbAGya+MfvBXxTirUZH1kILHSur2S9Xpp
zaxGTSbq29TT6v+ukbao0fyEDAtgrPlDeqEc2SCtaz1otwF1hYePzfTT7MBt6+5bMPwJOYjHtEZR
KDC2Jlq2Q/j2IbRtZPB2AQtgscCjgOwcNd3XEfCiYfOWdJ9HMPUHtaA9Od4+vpdQzMTfHTXAdWfX
6xnWuDubE2tsHEdXEAoq4/eRLkayet8K9mXZp4pzDbKPxGeKKT73COnxrWGQ3/gjASzUiOmuQsJ0
CYEVAmM7dH9tVkprfpfBavpZHplX+GuQShRpZr98idMys/DtXsS4EYj0DRxXDJI+XBChUGD3ltRI
39nv5e78V0aY0R4A+ett43aVkJyfke+J15vN2It4PF0zT4Z4gaNVfN/58EVnzleW9FREnWgOWT3D
+NLb27f3T18OWc0UniH9MGM0UOiz+l4CGlZYx3KGKxnMHO3HBBY9app9SV0O9OVQrzIjRMP5E8aJ
20OE8aKnzIq1gICNHs1Ug+EEkGUx6XXQm9TiD7e0PCoOw7nCL08to6rZjTD5GYTGqgUN2L8t52Ue
XWDeJJCdXdE6AzdPlxoeH6jOqyAVrQivdX0zFKqvqXXrLxEveIcBIrkUFix/wpWFqmA6Whql3B42
2a1UkgAGZjqFluY8L3UhwRkj5FHI935Jmin2lI+sjp2H7wg8A5qYOxkd4Fe+CfEzavxz/QjDC4oB
uOGQChuBa5eKoW85t6k3ZP9Y/cbVRRTg1p2g5TjvEWpH12DUiZ2aPCP7OsaprH/V/dmAapEHOJWM
z+WDLh/2S0IPKt81iwcr9XhQDMgTKczUQscotTRZtVWgRyrpyuJLcuMk/IUkfs1r7avBL8jyt/U7
vcb+6+3QsWArbAWpNF6FQMEXQ05nTR6AfxjM7duJ3pFZc4rd4c9XBhDljdmgg1n8kdpjWVWv6JWp
eKdBlwMTUp1/UbZwDDJ1cflsATXecfn9GAMQVe6CdKgX6f26u1kyUdimCYk2HICIvzsBzCw4Q/AA
PH+WF/PR60c8Ik7d2nC02WYPd20l5x3Yd+nT0wAlINRXwjWM8bskShE2DGzHLX21SS1zbfUSvhA/
b2/TdFpm8HD9FNSBga2hzPbUhgVSxtf3spRgA1GvPeVXowza1YDDWeLpVpkg/y5se0Q2JYp9raY2
ApHupyztVTfWCXGcGaqWumET7EQ4gFV8FXID5gE/sFFXD1PGPPWonZnVNaCUV3rFq4XjEv64WeXw
GlnYK70ncADYqHe1eNzjVbo5+G5w1JkJ0ihDG/Du/sie6LMC9tFa8ClSwaZZyesHDygq5TJMHLZ/
dtLqf0eeveVtSfAGOL8SxCpE45TugCUuybFiiJRAcGgZ4xN8IXsia1YQIrzOtiAnPoSIOQD76Ok9
snogkVmZTUfoI9fnuVZoBA3RLB+8n9RJn5XXeh2GY3h6RG4115dmOThhNuL0qaf+SO4dcse+Uq0h
B6RfmIScg2B+ZDaHZL4wF+CkMLMlwDTkK1+l20oVEpfFLHNT5y2hzEoza9hOJ8C0cO2y4rItUoZW
tzZBGDUL+oKpTt7V3FD0nsiEugvBhsD4CDr9Z7M/otjPHwn8ha+S9+Pdz+AxI8Z62OvXxRPUxs3S
ERcAGsTRLdoyFsqCg5MDCZx78u3SAmX8Fdg5tvLlY1kpda/rx0q6zm5J9/S/9ZRV0c2Zxbepsxcx
n1vatuFcv31gqkGgspo2kguzGiasmxF0Pam0K8vE8BhF27lptEGRqq48vUme9QZy+qgAw5J7hS0O
hLy+AQphIBcND9+vVde5hwV8UodSzrWvcyHynavEDXMC++ybw2ZTAYog2GW+WtAui5e8MZkg3Xig
E/9g4/BtBHxJhgDGxY7n8rCZNjJfhetLO4fXot3N9idC0h25Wkeu6Tcz8ZFe8ts5zRIwEOEQvZg0
bEyH5XEjDh81aKWfEDVSD4P2XbmPyUFk+F9OhtmtnOgrAU+3o0E87fVuCcxSZDhsvBjTA2x2U7My
sFQ7xmTcVbefC6gXrk7Dhuy0bhNgpaSpxMfAXH9RrJcqrm98p4l7hnFzJGdX+aM/2HW3/PN35qg1
Ryou2mXZ0go+Q1tP8lk2dAtAPW1OeXuitspNPP8zunnnEV2oCAtt5AnhCxhNYpRkstnNmberXdx9
VPw9P6Fpzsf3Us+La0M4RK96AjJG1mt/Ffu5VlmsM8vvUgiXDv9AL6zJY9ugEIFQSiWvUWapfYWe
iYv2YEZxmrc8LERdUkhLh5IV8gI6FLqdj4d0UQnlbLah3BCl9VFR3LkYP8PV4AvWIpoXgKYpevsE
3+9u8P9qhs11O5Nfp2UNXnEw8MZ5h793MP3D9Txd4TiC6tpHdbjxOT2uia3XzAqU4Tcd9ULDcaMR
3NRg4+8iQC9V9JHYUOm+t4zvwtbXu8fVTJTqG8eFTZ/FqR0LOCFOTNhMG4WerCNlz/R2Qb0vQNkM
MGgGYkuE/EAPSCOkiPlEqJJ39C2aY4HybTAH1dlALfEnnVAEe9NNEluDg9A9eO3Wp9gr0i4Ee8gL
WZC+dS48IRbDRjiDqjVxKeRgWkao4KXM+w2e1qg1qNarcGF6BJGqqioxz+HEc9luduC5m9QhraV+
H8b8+NsbkhBmeMXd2WzF9HyMeKE8Kse8x7NeFj6bJPqHTvjHUkOTaCxAA9Lla4fq4z58OjthuYJU
6u6ixCiFwwmNU9dPKN4DJ5ATe2XYyp9dDLv/wzg/aMUdgx4EW/rJ2VpaCFP4kSjV+XVz1wwcrvg+
AiCu2iK+3sVc3iIkKx5Radms0OjPKKcz3C5L2ZJOHO/OCIgYqSFkrYvwmzY+0CSrBtUvmaymJrp9
B/sPWCq0Cq/PfV/0Nn/P4ZeppN5SzSUy4P6v6GVfRkI8L9vS0tENhHxXQPIM7kGbXdcKFt5tyXac
oD2AqYg/3R9At3/JqJCQLg/QPBkB8CrfLq1YMkGdvzvbdmoELbXCR4gC/ru6tjfVM45N0s02qLQ/
/j8+oHRXwhiTgr+9VXqNLLbOCF2IKaqmzi6VoncLri5UCfOAaUp7DWnpXrnU1d8SyMUSf8pvvtmc
B1I25TcoZJyHZAY2AlBUzklPzfIX2btrs64CZMtji3ehNbrJMz6A7JfKQK44tTk7Mgw0eYkRMaVQ
aHRTw/Nm/bZh3tzDUlCsbE0GR5yAZbXYH4wd2p1MXSKx7mc5UKff7TpFpUTxZ7IvTNbXyv2jXjpG
iviIwElluKzNRzEg800yBR++/SUMJo2oNxqb6/95ST1dUbp2+IoBZbTw664WkkfIOI7ViumFTjDv
hWBv6ky7zW5DksDm3hv+rH1wiBp7H3otMIP7yJINS8/9EMEEl9afW7SKPuxCsnF3/fBhXxzEGekD
xfe1G0tvjrjgQN/fK31q45RNIx9vYrPRsTVlH/REmHWZINGfngGMzShrU7wTNyfdTZskZ6E6nYFp
+6rC9YkDK+aXTT1SmdVJEl9gVYiZd4Pr39na6Kzn3Mdv2nY9uFuaZnAORH7FVhBpk2onWd68LWwo
KWdJBlVQ2Dzl66wtRxOdOQ7caYVqFKS/titGSycyv33luEtVsF/TuwAinHCDpV/P80iD5VFOzvTV
nnXFJ2pjXX2rgnvVKQz+1dCoLB/iD2WQzTfKrGUm8xA6NEkmtR45Y5SRj0HddaTuRxuemYdilAwD
bUAp7VgV2PxjkyEA7k/KPSYLgvnbdt6vtfXsc36JZc3bryHljNFtYCSGpqUr/XtMZ5oPbUw2GtII
gykEtoiv3R5Tyuhkk255JjDkWjqSgPF6Fs9GKbaI+6JXapQSCHJYe1A5IcRpR3u0tsgrr0vNAOOj
fdURHqCdJrP/J++u/g1pOM4wcTT0LSGHzSJi8y6G/QvYU3Rnu8ECvY6J1KppimMWrXUkPD9IpMEN
gfwWfNknD/3ZxzOqgnmfqukL789Sw0gsG06P0sES9ZvdlDooYDftR26cAzuf2QwD6oPlCP9s5cTd
mzSSNQMu7j6MfbddY5f+T/CgJJ/DryuLhGlZJKU6v8VNqv5tY91wIba8jLnyozVG2P1rv/jA2E+Z
as67eTfP5jDUo0kcyX3PAly6KechzNrjZJWlKsk17q4FVSQmagIAH0ZDh69uTQfV2Y4DWHlDy/7K
0k/L/0b5jzsb2TeLsH7t3jnZYBZ0E3BPyHQeb7BE5/u/naWVWfdZ6IVTyQ/jO+04tFNVCdMc2sfm
rybGw8u4NelzlpOMq2bzS1oovjRCaFEPvoo0eou2p1MXLuG8NFWXbImZlq6w5gGbxWyOlrG7dwvu
boIly2r0BECxfLcSP2Zx36JlNrjtX0Of9TjXM1a7NjmB9/+ARdPKDrjlzRzOwDuIZ+pUl97xRPP+
buoOBSUkIaSSWeaV6PuJlaFY6eHKKC6J2QH6Gg0gBZvBWXW8PGauu94JBS7jGO+eEaZKNMbq3VWP
pXFPMuHf9BNPHmw0aigeBuBeiIJ3nA70OKJTzzVI8xgB35bkH/VCikW+foBY6dQHL6UXNM8RvRMs
P5mP5H5vURJgq7iQRKfGlTu0YBoyXRJPQ2Kfe/8Au7qjA++q8Ogu9SBoBPWpgLqTGjapcP2NXDxi
XKJ1w1n1+Th7FeUcEOUeUBVbvtDABVIWacxzvQ6RpEw7Wa0yO6o9fXyT1q35NWwWFoBleFSeLQge
21T0pbSxTUHpPi2bdwgt8vbQHmUta9wcfbIRx08T/V4A/AkwXho8GCgXD3Rp627fsfPZpjI45BW0
sNT3vVMxQl0fJdcSwlj5TFEheVhH5Zz+0K5qZzYV6NbrQpn52v1HEEmvwT1XPt2f3B8auqBcPQGH
bI6naWxlVu9Vvt3fZCi1gtdKuHE7rRF/OL54MlLS5leZTu8Ikql87Ky5r8BaWplcz8fW+REfdj+O
c1tq/iwa3VEQiB1WJJiNXGVdI87YqHrX/vAbE5zXI2Qh49n/uUNy5CwR52Zntgx9I5P1QRvfj7P8
CKZ4V1+HJXB+WkyaWMKtq3TrqNIcoQz2BFjViiQZzjSZMLlKNJXvusK6HHd5629/M9qr1BYkcpzB
pkch8iGKoEEfqIR+wopSJhB5FcDicY2wWRhnFLIA4vRyT3OwnVehgmVHcsql7aFtjMIHjK3NLiDb
GCUbaKNmsm6iIR4FJqqeVNNHodCBkl2DG3KofLBsw+/qiAgD8j5YbrpUsebK3FcbUZuNgvlKjgnk
3ZjttjCmX/pdIzHuZ1KkSXUpQ9jUQLxKIvUM3QtaYbvlpB2QkjZbKsLgHkMz4qSwpzdXuOYZ2+wX
wqWhrPWkg5LC3zAjFodCbODPhASKSyEdMStSLr2RwqXkmx3thh4yi3Y4vygngtQViLKVFYQ5EY2F
AoZH6aLDFLwMysM2/JOyFtEO57oUX1pVQRLXehmt0Nbledhr9lFMydJcw2+b9fKUAUd7hJaC78vY
CJRSpvILy3fSJ16TkLxI/chzNQuJcShl11hmmXa3hXy6DepvshCPbCh0W51CcjkgXGoLh+38FJRO
Q6PDkf8B9b53oc/STIHd8vnCE246/xhAcrfFicuizDJAHPzAPA9IsiD0ehdFsOAfMOOPehwlBP4X
oeKAu/erXAOnNZ8rHyxJMnTYiTcZzaY8J309hBrjrIm+6A+rPAYCPIDftCVpf6l3IbHocOmKVRKO
inQciW4mfe1klNqDRFOI2pSGC+9cBfNS/BSoetg8BSoMPH2At/m2O2qq9XfdS8UDmWhp3q23gltC
CeJSvwQaJgMUZRVLmkHyhS/faSDP/THtOzkqnd0nHW3WlRxbv1ar2P0DZYrGFZJbiW1FnrPogx5G
AE5IYY9QPgqi84ddj4PyUzV0JmNHkTvEkX7mLTS1omYwbSGNQnWoEg7SzKnj7Wq0Rnm8tmB0rjzQ
vGEoEoCGSQJpimPR8rg7EpMkzHtAiVU9ixeRUi2BtdlDfAxZBFauu9gdTjaQS/6cUBsYPUUWcAAv
9xZtuX391VX3fUkZK9HfCVpHminXgg+7fEpqNAErAIlHWPBTq8TG8vAj9U5MMtknZ3/dLiVP6UZ7
6/npOd9ViPC6v+iLxeznpC8UqkaJMgWk9K9aRRduNf5hcQDJaeSGV3AkQA+4SOMhNH3+2+L2G8zq
8U7rh3Y0soGILyCR6voeRHUxAcMyxVSBun5e5M9yefGUGcc0nBqsUzWPM4STNrpZujL5PuPZeY2s
pwUFWHsmT7vwP7m7r48sBL/pEgzDxZDat2gM2LwQxjLJ88wOicAiO/aDXSwxACWjmJiMVt405+TP
orczzZrpLhVTvHCNGCRVOZ8bz78PRu+TW8Xb60cwLd736W4ZmfXi7HM7IEqpcvuXLUjaivPd1atH
cyvd2zxegyRIvXq4ZEjui5RU5F6oByYmFyg/ZaAPWg49invsl7+xYnw3816w4FtpoQOcoDpM0d+f
2WXHlJKi3oNdWDE/fiewE1r2XbOD3dlOkYHZu2HUw5X25odC+OdkCsaflPcJ9o5lvmdeT0yYbmnt
U3FeEpEq+UqiZ4v+5V76E1j4haNvAGqXQ/AaxdXDRPLgxSn3jDJYQHLqKZmgtLru3bVOv0zkNuhz
ppNXxZxiVMYbBKhCT2T57a243QBPaad8mcVyk/lGu8EWlJ4VlKq0lpB3Qc1NV0lpIbK3QwIVvBR0
oA3YcUc2zrQ/1QSbFgTdW8GcHyFxl8+JOqUTwTIJ7/f4zF4mlgJKa6EvD3Bb/94YvOgb0UtkAtZB
95Imag/Gv6Aidfsu0F4Ey/DKyvxccXjMSWviEH2/NtHdlU5dVZdltc7CooZiRvPatO3YNONe2658
L4kqf8YcxfFrYRLu44ekwG52Bx8dHGM8fSddgQtEp3kw6+equNwQ0QhZLfZMxGa/NLkwcIpfZ4eG
RxGP5SUHll+NVPIbS0fzkHDHTsUi+V+Wh+s8HSEE2r3MExRJCZR+EB+Sllaq9KkE6EO1WggHqAkJ
3EsBOm07I/4KT9VCJoxtgYti0Pu6OMwtQMQjdmgLUNMKVj2ldG8ve6/8Qkpsb1OZSmMPb3DETxNc
7P7uf4R2NZ7APtMBR1Jm2TFciBahB0QpZaQf/8cH5rAwCajaPl/oCeOWVvszBoH8gbXxvBoaODEc
M9yHDq5gJSZP1cVkXYEmgJqMCt3EiOjJbwBHNLau3J7xwGxTTBP73BU+UlMM+Wn+NqLjVIZZCwxN
tLTRhYorpVmu3FuyNYRmis2T8ujOGqEyD0PIgHX5v1IAfKxVH1KhguizzKSYBh8aIFWvhjCTO6s4
Mv5J3NS2W5m9LyPUAzD9tst5E+A/Ouh2tzHFqWeT7gg/Fo4MPIY0FAz9vW6vCEvyKuqes/cs48hy
ssMiMv8Re1mbwHa/eRPS1FiZz7XmwkYt8E/u3AOmfg/f3iSzmw3BRh9f1aPG6fkpIOd0QfLmzlmh
3LRBEsimW2hu2MCAU3bBg1VuXeRX3WfXVtZw59VJ7pM6yhGEW3uJNO8BpLmYhDlS9v9dyghhyZ2Y
tEZ6Sv5z65BhOJX2L1W7FYTt2XCcZsx5fWo3oUew55VloHUSA1PyOSMVucqAscK4ET/WulYp7QKI
mUeC6QNbqG+vzNNYRpW7XvrmGSdKYdU3iVNgoCtLG4CLs14gayMYr8wK7tcBg5ZAd8vJeCjJiGJG
ZmpRoYz+fAybwhm/4GjpgAAAS5IV06kWHFJrr7QjcXfm7t6c+OZ1+Y5Pp8TavcCQtyiH7XbGzkwY
GMBOxjD1Q1eQnX4/CdYa7c30e543NnU+D4WAwkjpjJ6XDa6pDeoybnvXVKUw17Q3HV06inUnzZQO
YwQ1Xeix5nHh9g/Xjzl1XIZXClTIAzF4mwciy4TpRvUh5dI8GPE5Fv5fhKWink5pn2pLhDCZoBnA
SxspkT47Nl+BDq01bGUyOwWINkXieH1p6nw1WBsKznHxowlkrYjbfKjqpNvDRJVw5vnhAoeppmkq
PD+gv9DFu5YyEGZRxk8Srq2+SG4uqDx5aT+JYf/xPP6qP06a1lMrV0v0N9ZKDG9s19t/8dTt1nHY
1EaA9uRlnf6jcpSf7jVBh/hmgRmZoNhArgMuie1ag43Gw8fR7PwDqrkIyS7mOqtpfF4lMQVvgKDf
PBwUbl0s2oFVaf59b/XzfQvbq8UaBRCi9caY/RZig84FF1NnHP3m6HXwLJ9npFtmb9uegL7HdkYR
9lLplz3p+aUPshtyBoq4uXK/jKVuxKUnBpDvN5lt1htEW001lhHhjY09QB3LJG0eOhY2cVTvLcOY
AwOuguihpT+ltL5kKuVHUAIjYv2BBWz7WgMZx5U3v/rJzJ3gF5n3/P6pxmdnaUOgpiPBSXZ278Dv
v5V4ulUVsTc4i3B4ABFMwSDaggC+5s/fBkFSwF0uM29c9loN0e3mVzBCQdZipt5d1a3LmXGXt94O
oCTyP9TM0k46g8m9JxKPWyMKNDqX1L1WMLw/NtWtlM2NtRya5Q3pubKEgbyCjWQKvHSyxJz+ato6
UkCTSvKo7pw/sSM2rCGhYovVv0NohkWqBFfvV2o+aNwGqqzjUEFzkON5GXg5UN++vyheHxQ2xYCP
iGVQxRhrD0qIn9qvBZwosUinIfa1drFPECGhJ0kwrov/iiqyJxGfb9BiPt6Cg+J41N4w++xHzdWY
hWYAxvkv/8cwV8MJ6OsRH++81SGY+KmCOSXMcsP4e+Fd9kJ39dYufoYxHEX9xUt+PW5oB8eAdTtA
j7hGTMjN+MEAJ6QuSatb5L1xsFVzfC6i2KI3Oy8hsCuORhYmDWpLzyo+3Xco3jDh7Sapw3uJZ/hL
owmxG/oPIYGkKRCcYkthzGP4R8fx6w+B5bNHNPHxEeZhkOYi3guXWaf2B8cxK+nhJob8H1tIQqmt
iAd5VnqnPNdzW4+M7EGwYlGcQk3LS52n0ypwZQFc/4ZqPM3QqByAgTgdX70gtQ1MrT0K9dPwAOY1
cPtmJAoIr0oxVfF8Yx06DDYfpLtzY0d8576xeo/ll23XAbu1D8hzJP779GlC+41+E+CHysrgnYEz
YcvKrxD7MuMv2dnu0Py3F1rQIiS0cTvoWXJp2WDtI+jzefFCJHdOScQsKc/RDQ3b3nnSY/tq8fjk
SBIchoD+13DuJcZ9EhiiHpa1UD8M1UocLvi/gUbyL43hnNV9+1sYlLxtje06cVRyKaA8QcHh+7YU
d64fqM8A0rxPpKMjWp9Kcas7PLCZ73qjgVM9Jcyv4UEcNNCJ4hpcci2vYfELstn50OdYpNdM6z44
UyijCZLnq6dGQhjY+Ur25/K5/U3bIR74OMZUIoCCqWNanakq/8Tv1RHR32TEwjBySBl383FRAcog
I3Cd2c2wZAUjUacGEXl5dC7zNuFRFVtuJ2h4SXw5fGXOc49Jh4vylsuhQdR/PQCKnmhOqI5oO8F6
n15LnVvAQKN//OIY5UwZ7CvXDDJaYlGwVjqYsmuizmL23dD5khPTZexql0R6etoWqyhUy7FBnsjb
y3U0Na6i2KCDYu5WSQKp/1dDuIIE06UZ9GAmzWtmuA8w3Hry2xqxqI/mjKrTndHKKis1/nFhnn6T
iYGeU8STwO9icRTcr1yrhVSbzH4HiL6hvlDmXY65jJ2CCz6Y81qbylwZQM36oIaSiRHjQ2Ev27P/
V6TPDe4inwRP5xDlzFWAHT2TbOiXWhRRLU5sNJv9PqPe+VsDevfkybXMT9HY+urhnp5X2Rb0F6UZ
AjMzTGuFXPuE7TPjx/vDWXSjMmDHcSZCVNXReDLSRRMVYopbJm7bAiNHRwYFdo/WpN+ER7Oel2s9
EQXavovETl1i0zbv4F2tDJwmhImxTUzrsJWK93OtncxZEuMS/I/0vv2nwNb5Nx6xy3Bb6Rm0EjNR
I7IQkGg3h/NzxQz8NUlBCJ+xoIGJpg6d465BtqjUDt1mZhyHwV/HLNrBVSWPlb7kykYukh8ewKvr
EukqiSrrNSXjZMcwEimMPzTXLV7tkh9TgHPio5t0+K+g8KCtG7S3d581IGfHCMX7vWWIB6gbbZmi
P3DhuwogYyNGFQ129kV/v2kFn5p3AVY9QesT5nb8XFXFygzWPVeTj9VfYG93TvP/9f8L9LfvkpmG
UHGUNCF8iiK13UA9aql3PCJXe1JRhPBvq9AKXwMA43iNLYlw9HH+L4DWvbq8HS1S07fai4FXh4aM
Ba3+XugMXO1YR69orotH9+nWaOGx83uC8332o1tvpfm9ABm5EUMdro9D7twQQtv4UI8rQpyHQsLG
vuB9bjlc+VDtL+wAW7qUw4HeQ5qY5zBLbnKrwdBtgW5wT7DFCNV4KBr4/aCZZOJn5MNSUEV2l6WE
MfHyafOklpBsh4n+GJqxSsiknNuVG8nBsy+yARkqSaHCivxHzbkADedAexAMtBQpsQPI/epFJY3s
H9/S1YzWltHzuTA6k5JUxCFFveIesOepW1DAi7bkYnVqCXsiwhs93SfTt3LEqazkHCPtgzbIwOe7
Qodlg8jr4/SOBrOreVhB4v5nabXw/VTVFYT5HRdqJUalUg/KVJ68BdsKxHPSSRxwWVzaJBsJ14yy
3T23llkpLujOU+1yD1AdzSzmJkprskR5EJbWk7Qrfrz0wchdLJ39hYPPF/eDF1XGjetiY8OBRzRf
Zf7yiVjGe/m8EhYzSWsjMElbOkMeC52LLDG+OL16YdZl/Ev3Ofkq+tsjj84ImZbVW8S7aV05BSUs
D4vCLkQqOItXVO92ZY1SMK9NVOClpdRM0O777z0jH0kF0xrFzAxySuTMGHGw3/oaBGH+bNv3rO5F
5ZgUNZZobi5UliWEqY92b+oEggLNGy/jCI2gQadGAyMTTkRIi49Ed5kgjuXZGTwKB1A1py9zAAQC
+/APcKFSl7JIjv9WRqLEunKz1/OfsfERQp2RknQtQGHRSjcuFEzhPLQP5iB7xQF2Vp9BRtccLrYw
Ec51463CeouMj9VgRCzGk5SCUFOjCwDWpm2gwe1wb11va4IUfacZudtlKSMbNgX5F7crjsjM3Q0/
uiELKrVHgCS9JFwzUKlC8BbQCYZF+9C5nswn/8LEvhviy8s11rMbQr4+gDtmur4YDaBIlcQZlaQT
pN+xaPMfGdEXW02imjumBHEwuvyKjsub97dGqzea3CAPxHJf9hulrxlARG70d54w48LHc6eBzKgx
GNpTQ0R7mCpfTkY/XwFECePTdPzjrA5cJvOvpNaLAstYzYvBEaE5GOr3zMRDgcE6IHIXAr2Oam+s
kSc9MlapasoRih1Ha5NnXEMmC+swPA153sVt4YpNKk9QDFO5Kx2nRmzhks5w+gb+a4JPhURhD8fe
dXpfRcJn62Zf3srKArj4Fp7Kbl1p5jHdL80T/3Dh4+XpLxfK7UAZ/K4XuHzKS1nl/k8IpDwQkCKM
Cj4D5gJf8i8FDLDeroxeC23eL1Z6Es6FLZaqVOeH3RoblWAyMkfV1kySKj1ET66ABhgMXplwh2sN
W+ca1GqLP9I4Q90ZVl65wdq9q1oXf9z69oH8z+U4Wd8obaGgWbrnbjiDWr1Kgpu4uYMBGcml6DjQ
mMW8AMwDrKlHjVjol2Qu9jNyD9SFwYgnatmDNKoxhkcAoj/o19lx2TxdK1dtQqsJVHSd5EkWZt/p
x/ESEdLrGE14bR/LIIJFrl/0e9hxX8Gua3C5GpKRYJsrpgCgLRJeULdP3AqBGG7KEbwyX12fx3UT
cLiAiTgOZ9AdZCWve8TqftCDxnYffh/US0iEOMHY5BFBTzMnKxox2GJfbKidxhkYb8DtX/mF1at4
203LZCUzQU5yRz28OYMHOfcWu/c7Qq0sVNxkVqqirOCp8B1nhwWhpNFrhCo4eXnZtMhKqcyf2+JJ
NOGhIIg98UNJsesFpk3cEppUmj+En7+fhpsJg3INB3TMoLJgZAZBLFkS3TBCTux89ums2FypIe2H
cv9i+FsGgK43oZpwLLgjwIcfH5Rupfjhgfnp5bRIwTUsbZrAEACjmB1MIjb1OUWDDrUPVBz6fuU4
vMxKMmnBzTakA6nnHtX4ImSE5zQ0crEVZVjQaLwjY4IIwSG9lpfdWS2Pb9q2ZI0Sh0eLBt582UWc
lTtdKtJ5Ya3CXozzCrF88ZikqIUQWDcSJmdalev5M84CGT1c7dfftIyKVRR3sJVJ4ABpjVBHuJGI
OfVOQkTNsOi5ZXytnMJJd4dK6OF2fdT+ZgiRaoldIm/AUVdyHs82jiva/rg0MKuK9gDDSMahO4J7
VP4s1yEbEwfO1WyoF4sTlMwz69bQj9LReQwOuVkwf2SoudU19//ZfMQDBY2EeS2Jx+g6cEmnNBhM
lJp9eeXPkIKLdJgI9eAIw6llmLh0c4XnietPS0ksQXkiwGAI45WOJXMLNz4FLk9gTq7V74nUpq9J
pX32fslOz9YQuFT3C21O2cI9/yo6asoOGk2nyjoN0c/j6XCo0ny/aB8IiHsBo+HN+xQ6hu+5WYNU
c5pRa0IE+UFjeo/GagPqMLmgE8SukoFNGfrspvfSy7Ck7DsoDRtB6lmhB76QswitCVyP86VPJoJb
xLJT6IZQAI6Fb4kEwME0i9owxnk8XWd2J8vx0WMWqtub0smgCW14mEzgjknFpUASeuF5G6KdHuK6
69/CbENoW/aB2O/fygmSUaKkH6m18kwqkiH0CnyulVT/bzzkluR2bWrj1fGo6B0zQ9sR/wTGO5hQ
xEFU6f+IU/IHLR0Vik4VGcXLhW9zGItLVS5C+VqUr8PPG9VpcvNq+4jIM2Xd7ULiKp01TD7femZr
swsjH5yx7RXtjyC3buJrKimdfHt8vysOeR5bl4YVscDlbmBNnAL7NJSh8UMmq4476cneefHsMw5b
TJV23oaXLQk8Kg2noxorb5cx9xpPw7E0WzQrG8eKZHsWd/tx1kcn3dDkGBK0ipW/ej6up/UMN53g
N592QM4/sjsuCJRVT+TrNtmEA0wBY/SjCvgdgdQKLUwiD3RiESGZpyTwJS5VP4TfETD3bG8fI9ck
plGf/RUwJLCnklHWN7BqnXov6Ped2d/2UKYJsEBF5jwP3d2AgYvQNXaqE5pQrPNMqhEY1kGDVAbL
1qugfiOWpJ3T1BSp/Y9ys+I0dPUlNS/4h30RH3+WeUWTGZpqgNhYnEayL/wPwzCIiCVKehnLNMHO
+ey29tGIFGcugaL0Ut3H8R3B4moB8crm5Vx0EFdTtGNRe2uyYeQP1YPMAi3gvqPMOtD237ce5vVn
OTAmF3qfj3dqeyX5N68pwoPyzETxgHZRqf1BTgP2MHzv4BNaoDPUpZDMEykPhBqJXlQNWN2L+UsB
8dXMFbqYf6xiBHeQRB7d8/UfD1zimQPn8aXhWrJCD6lqWJxWiz5ycYMyD6Q6/jwokEstJVOWJv17
l6itejPeGY0BmhX6UYq9DJWKKLVMVSM8u9UxjXkK2H6vkxBbN+BaTsB4hlKDkWXNBTXHqbsq2b6y
tJy0NVQDO8e2yMninbCOf+Z7PkR6nZNASCMkyDZZgZPQBsQ7MveEpqG7jIAcnpTYmgAzO8mgwPjk
+78Yaj9KQwD321ADhB4lkx44hAJXKQHvVzREBR7hNsui86Sf/rQe1u0xXoiQMmYFJILy+EjwXETe
x7AxSSgfpA65y0gM/oVKDpqyQqnlynf2hQQMOOYvGN0bNONeYd1mdm4W5CgWJUEfbpysZ0hU8VAY
+AMqrHQd6i9Oev0SuFBAlg0WeSuoW01VEhjGE74UF+uRFBWJ7sCeLrPOWwjTJH0QIVP2X4HoZOdh
gMIApS/ZEzzmDEYBLkj3LiiWF8IrkZQqTvNvoWGDmhFqJAFPeT1ocenh+XVJqMsGmsWekraBF+X6
C3eOQBcJmBEPQDmmoboTq+AG+Dg3WxWQ6ZA0QBEsT2L/0iBLOF61v5tfP76mdYDHMX1z7az5ckM4
i/vgBlxYDsIDx/g4p/JIUdXqPbI76t3Oe1RShWygzgenHZDEXTqqflBgsKj+MJ6ApaZfxf48F9j/
XwSS8i7wC4ejuapI9IqUoZ3RzZsC84uLd/dpTzdcsz8WwqiV3o8vjs/mGpeKof0dbBaq6vjI7f6D
C8kQPVvTQhf8R3kVEi4MFFUw8iXzud7u03rZR02PGLkBSIF1GEjVG2fNIteLDUjq9x4UeYWi48nS
BLzYRctTfWxGSJHEG3LuBv2+pgGiQ/6jM1NQcr+Al18wMuzSVxP1FDkQncfLd/t8fldj44jtkhSM
+/77wfhH6c0oRG7eQFH71s+36Sw/g+oK0p3z5OKoZYRKS9ZGvL80x5On+Zg2bReU+mhfYJbn2KIk
U1p2FiLWugvEAqOc1XdS2UuUEaYhS5sSPYqw05KhWTXoh9lA2f6HMCt+Btw3rVBYyhU4n5HAJ9IN
29uidVypjoqURfvbX7YvFQNZNmFXIu+KhSe+/Jc0Q8/ONLpsJTvrT8LUH31mB8nsBDeI3GXXPOBS
jgR5Q4RhmgB4tt4tlverlULmt448B4HtF3VAz5bmR3pWuLDFqaLVjPzc0DQ5bh11S0GlnOacHB31
qXKnf9D4qMshoO1i77pxAcmwVg6WFmq4pqJiNCwdNdZNKEAlBGL+3StHSP6hhHl8BkuGwL08En8o
QlnojEVUl4so5KlYQXp1pxh1Os81ivEF8WYN6hlXohhsX/jN2qH4ZMuNUPs43IH2Z/zsz51CJ23d
re6BW9Im+u8aHTct7w2HvICASCD8pfbgdi8i//GEK8UCT3SWZCvKnydE1WzgXMUA7SBWRuvzsNQm
UfIiytimGHKW5hFval5XcToJMlgxpjfjGvHnm9gVOxomTVZIyUUX9CE+6BPEzU81DknIpGaIEzg5
/+YY8dWy/fimIAdYlVQZM6SgdCQb3ZXUQ963C/vVk66DctHfgrQbmx7Rh4WXjIj5NsjGlcoJp1fv
GjtJlCNyXxzXh1GgqOxWzq/wyxRDHjv0PCoFD/9n9iHw+lFZDSonk5HqjieEZX4oOl2VYxcY3tMQ
a3KZCE1FUvQxjgtP7GhL8zhmYVMBoMHhGjqg6KqwMmx4kacxeK90ToSmIcMcWtraXEb/+PRX3KUu
/rwydNh1c5iXo4qdsi4oHrFpkNGD+A+mXoXBBuJ3G6pNCa5GIVRkKa0BjQkLFyYnfHIw9ls8S4Gx
25ikCvCZugLRREPbR+RaUZ1JK6QB/PGsLsEa2VjY3ADGcwnxMeBYmn+dRSHh4NlMguqaQni3mNr/
LlWgjqGxe6adYuetOLopGKmex0T9WygxY8KHTRI5nfsgoAR/4j3o2THv6+HNxcH+OusJMLkEBa5D
rCd5XZztIGnIcUI3H3XQZ+E9ihIrjhqBFLt+y+5chD/MjO5AUV23eimYulxaAiowm+U3HuG/jYuG
eSTzIbCGNXT9zLjw4HyPYPYJlsgJu6h5fbvWZocl2KArATqjGDfacSHKSzufqUoKuLTpbFLCpmma
a/PnRMkaVcISvycBu+n7CTtnavxeUIN+CCjIBk8MPdKzv/Fen3GKcoE3zSVZR/Dogu1qyfVTQsJ0
k5KuXpLJZOCVCsq6ZPdzSHsMyoY6corcC465RHg4iRbQeWfPGXEVBr9ErFzcD9OYqLXU0SbzXKgt
1oTLWd1JzvWPdmb9cvEMObEt6LPQUutqjjLqTW0S33kT3ZQaBbS6hObgqQGr5zwqxcRtOGIZEaNH
sHe04pxtW87ISeZcl20nsABDPGtdF+FLTM6TazYoz6p3lOO/Uxy+85g5YjkTy/bNhWZsePMrDwvc
0+0HiahOKT841EHu757sigv8Zudn9QzsTqhZyQv0uWuGcDzQvzmPwbBmuZ29F7SmrrD8McLgf/+m
w6CV2NpDlsHt+6yGBdTGe/mEaElYMVHxIf1AwaTn6pilLnMOVuL0bW0XCeq7Nm95qGms0tJZpmOw
w1pwCyz3KVc3DZckr7Cwcp7GEqG0wR+V2uiyIvDemDri/p0qHESpIVgrSgm8uvJASACNx134w3u/
80Wa3uFfc/5AWowu9oSqBZyHgsD6YrbJTaugtfXAmQOGzTOsD3BihzMrJkh9/P2KDjRByeHJ3ruQ
KaZWYuWoGuDSDZZz+StZfKrlkkkxGqxW/sZkDmTf3SIclbG6vJGeZ7V/f/eeasxeyxE0mB+BFOHP
bsX0R8lZBwGHKjhW1+YWdBpOB0beuW5r9lvz0RgCK++tklz/aAMZ+qelLdqEqY1n+TLxF2H1hHzm
NDMbyPMeMigGRLwpOxyZGdFxkowooHuMD9qcsj2TQWPqzMuL9Zn71WESe12YCPNPCz0ot7tUCYgN
kV1cx369aE2Mye3QTKnj453g5AL2QqRDVVHxOjXyM4EUigTI+pvHEeK9zXnlQYqVS44pqtHw+WIR
+mMS85DUqWRGoWao1mkMRwTQQhx8dqYjbUu1OS4SwDDAfirTH+sV2n3M1qSSEJsFVWPI7aWE7fTQ
q3KHFQxh0VW/aJwzMSvp85wLT8BgwgZtbCURSAfUPFF4F53Dag7rK0Crid7EWzHa16+D69NRrWon
S84cG0NZNLs8upfv/KIQxaI8BezLWs7Aai0XlLxK34kDVoXAnetG20nc+a9gYtN0/sYsOpiXaoeI
HG0P2oM2u3gID3WZLjIk6PXYTNyxVFk4/V0Ht8wBDNPMBVT7nZHWIqxNF+ThHhGCSuvQ3/Um1Alh
KdsjQmaOpZy1gKmAm0awE/dfBY3UYa2ZmtgvH18qKqEWwzCeDlWc0a1U6PynXELzOcLbxLvnz0Nj
jXMkLMQMumdrTI7PVdRkRPcdoRyOsinEqYVEso17kesz2MXZSoNNEx8lnljZR8gx2FJGAXd9nsNS
+mE7CqVG1ZSPerU3iR45v3u+KsQZwzmEPqdSmiQCds42MLR4CQp3KRoM3xsQWwGAtH2odJGlsiC3
858XHEntzcK4xQaCkX9tYcLCgVsmluWVN/BK9xG1GQP0+35yWoqYTHynLCeBZ5WHZJ54yKclHknM
ZYtoIGr+wacQYxgp0ghGRCNG83fqJXsRTDVvlwgf3WfNtYsmo9EPxMo2vcaHieMDHVgRPqmxS7oJ
skZ07mL1Gdl3Be0WtE6M8A+leVvkMRjGiCu3tlQgnZgoZgaOr3QUldZIzXo/I/9tLk2zmLsbbXWX
2UVSbh3zXd/FW5WoyINfjj2k3aNzIFkBwX6Bwk6Hrd3+WAUMZjUfPfv3bKww89Q2hhylmGaJJi8O
UsFtOqY/XJ7LW2og46xgJZFYlnL7g6wbRfDQ3XI8Qmi/CBaXwX1Bp+b3M0KYVc2lKx12kKuMKYh+
JTx4UiWUQktqNJ3ngbjYY3PnT+CvCMdwHxPCvNnN4M9P5egqyB31kOi6yTRJtL93jp2KkjDSjfdw
mfcPMcahPTKaHstiHdVSvYA/2CiB/o4paoKzWipd9V32pWq2zp+Xt98qq6b3YdyrelKu9LZOAVF6
buYfutHSEHBYCQU8/iY/P/YW3OVzmIvfWkmxI+lhoo1ZHXTxTESVkuVBxmbEoaz33CQ6t0V4TPAB
rkPnDbv8L/An6z50BqSKnSuua/c0EyKENZ7+h3wSNrQX3VAMzyzJDKnOTnoQkL4fe2mz+fO7F4m3
DcI9XjT/z1HqZgFM5XzTm8p6fnDpRKaA1g9oHM77LDtgGCQjop61eP0yzeg6cDp94NyNX/X8ptMU
NwY9eFB3s8lxrRF5Mway8DYDKNjdgHizJdciBPmjn8mKEEdLKE1ACv1E+krAoByhTwjHxoUQ3DSk
hh3TEKnOFlEygmxP30jWP7r94+yQqXh4bAAoB5d3wOY83kveBiCZBJ8laZJbcxjMUbNiROMxEf1X
NlM0koPw0vq5N3BPPVeO81SWGQgRsNfGp2TqZnbwn+Hdo6v+g25ZMfa4+jEmA25ngjKhZwe2FODN
w79nqQD2nqwm7WfGUiXqgiT/G89OkR86VitnROnsOXbNGBM6CqdG6O0K9/YiSaoJC89AozCqF9/P
u/NhqIDl9EejnlX6BQHM80zLJRXkULA4UlgmCyXFBPCW6yTmFZVvKKL+DaTSafEad3rpoYrB/6bl
91NeuzDuAqng2He1kzRiHofxDkaU5qlpVnor1RwFYC1jlMGoffPB5XrdP+GohGY7buGMnHaUJ6Fb
mjrQvAZ5eax4v7O9T1u8QIk6T3ffqVG/4Pm7TBZfX5xP/5I0/GO/ONDSZVIJ3fFfHDlJmJ0Ajg6B
sNACKpegntSB3uKHz2OSFNpWDvdDEAZDYPYbKntTrHWJf/9hjA94Ant2Tesm1OxmkDnKUgrTqT9q
8YH17XajJiXTY255ROvcfRsiP3tH+onS88DCl4hucd2SXaQeKrJZPJ7w7C6M/nDPmmw6P6M1GG1l
X1+9h6rA8FAAOpbrS0P/A3ZrfNwHVtr9a2YsP4a1FwNOQ9RpIHzucLYpsuGxihtZInymQzvz4iBz
/gKWAGE/HQYyBzMQeSOvo8YZdbTyhZtMmBhTV8n/59yrRf5XIQFBU3hQZHOVZqHqoCxkOkrkvTr5
ntEN8cXIQ4TYnr7xEFQtxRQOIjMk5uyibIO41M5ERkZH2SwKvGwM75AXW95jWJa7PSPMzQbssCw6
2lthX5PDQmb3zjTa+4RigXH7q2Hbxv+O6gXvHN61GJrKs122osGY2Zgz6sDiyZ6wZaP7dbDtIWZS
yWPPIrS/GFtmJ1p7YRHRxMKzpHBezcZ/XlhtBGwFaUcGfVlwWIsjFAU+p2HxG/NkPL4oO3Ktnk4w
HngVJSTcjNpgk6FCmQjHZT6LC1rXpSx338MZqziwTUrymF3jYzYyrTIER3i6iMeJ/zd9Kaxt07MA
DeSgExW/gg4MyzdDGgtugkm7F7U7CccLV9GeptbNz+QUZmHqLhJ49b644iigCuRJoH4e5NrJkLIY
AI0dK3KG5r68RBa5zuVjX01J0Ozl3Ui+dvgfhIlvhglglvf9QVZ0iqVy3xkZfVD9rz5NKKufPz/T
wipWoN3GxviwCFAskfcBsJzrJ0WMOk1UzQou1KfpNmZduioNAgC2INimFX8AWARwiBMRaus/+jSo
yFympGT6IsqZ2r3oEnvoj286KiG1fcYfUEeFhZVxPYDiOZKEw8o3wNmtZYKWDuKCrVF0hx+h2l7z
Tcuy9NzMzfrejwh6qac1eVYxXaKiB2J+JFvz4FA8Nir2xHiooxvOZEYiDm8A698bWtu64O9Mg0aH
PqW8YB27IYb0HII/QwIYQija/N0pN27+ur4dalAD3YuXmsW4jfhdY73Lqrwxd05Yva1k3qiwkmTK
O35++pqt2Sn0BNhmPwn/oOvEN8Ul3POyffTmAZCeedzwvdtPR05AhZQt1kjMMf0SzaySHAPfRGRb
osURNLFIpOI5SyJ5OwIHVOXwjkm8tFs6Y73BsmcVp2JQDe/4gTcUGpp6CyRYkwdnQCxVpYOyuudc
RNMRk2M+1jYkamjRP+TdfacphrJgUwrlPzJ99iOdB5sjiInSSus2/f9RdveeOJv9ZL6cmphE8DGF
WdorlC94tsDBmG5B7I9zvwrx5MN4M/LKPK6WUqsVCPI9R9Eg6cSVZo1FV5+OWDGGmPj3yfVZwA2g
q1A564f49893Vk2BbwNYiZIbL85W/fleIYzr1lJ9Stw3xBUFvQ8/aOqYul1UejlJMNJlEc44phi4
C+E87F7A8aX3SZ4sTb93z//A1Sv0E7t59/vkZXR6pKbIw7ZYxbbLsRXXjlGqKQUu2YTFmDzf8lrU
rlPS6m0YBIQ3tB6w8N8ymfjs/P6UuuHi2r92aDfks/ozweOcKOkciWh1kfAhB9IEO/cno46Q0L+V
AhFYf0iN8uChHDmBzvCaGUgo9QO4I9SZowF/O+kO0hzze5+ky1RrepvfuJdRXUkUzxT51nBdG3j0
7P+77KyZurutu66wPzj+N1M0r6tNcQU8k3M2lEJlEyz90vFyV9YafMqT+8tkULIs12yj0NyEwhuM
JgAwdnTyt6lQ5AcbStngnIdWBA7E8F6aKUR7rChP1uEiUefJhFoZhWJMlegv9nHMQl8BXYpwD0eE
FduAzXGgErdXlVZX1tWizakS82oYjEpSy2NKUuj3cz4emyjuTSsU+UH1Asr5E4xCHngdP/XNb3DW
p1tOL5RNFEuB4E6mJhyi+m7z2fOvZ49TrgGREJMGmjym4hUMQ7vSKGpTvpdxbwUTrpZrAvkFQ6OD
rZ4/tHTMsjfODMM24a6oCjwV8KaMwaU6rauI6tXWAoPRnR25JfEdcEdn+GYMVsAeap15moR+ldSm
N6fhVB6YcQnROAxrY3hCZE3bB5dwRFE3LyFwFQMQO6Pyl3CFmx/z1eANRFGTwfTvCHhUlGZwxIkP
3pyLI13luHWPefbATzWJGGiiahDJ+rwXsax1P2hhd9mBYL8Isxy4Y6wZTjMBPkhhnnXIQHeoUSO1
v24/+99Pld3v/b1+JiNGOyxjBrayV5Cd9cNWBsnasHclgFcSWB4A2e0lsHKp7YqMfYq8gz0wyJL4
i82isl3ktuBnVhgAff8y1Qz3jGEQFFzLYwArm2o1Ma6ZjNCwJuvZJU2d5uynv773ZMBvs9hoSDiP
Lv+XstW3tLciBkWn5QhgkASCh4zTg3WuvOIoGhPFg3Y+8wA4J2XPNg9tCVl9Yy0musqqHZPSp/WV
n4rh9TutNn4gHQ4yoYaPXaTcJYz3Ord4BKiBeyPnIWBxJMdEDUeqSUoC9I5jVggbiHbybVSTrEAc
g2tLBTeNyJmYuu4AnHzwZrzdarrwSSSPc741K/pE0kMLt0S1m8qZgJTaNVZkqCIKpGu5RSB2oSok
s+zHReMgYwgeETw2kAPd1oMYF3rvbF90r7xKQjLcoWJd7SMZ2edZdoI+LvWWjpEl1QXdYwP3YFVA
4uRxj7G6PDv6D9UojliFN8ss4c2Vdo3YoDc8qT9WUW+/P2UWvdEWxdRaGthDdRxK/nSyWLWOvBBL
H2cyF9OFWl2FL8SeAmUCR1zknSHA+6QGmYxxAChFCLEbjSqY9dZyqENODsq3NYHifJp/BfYHfBSX
O0LrTBwVUqxp431bRFdfTUc8sd2o7H4DicMT6Hk6yTIFlqXSMW1FPB+lk5e7iwZUk5QiVlc4a0nx
4b14GnZvFKr9rkoFovClau1egPuNHp9uYlrszygdJi4zIpL8XFmFmqTRilZzXC057vyroj7r4gDW
n18qIsWHCFhKZSPXShQQM7pl25ztulEICKg5+NQxnJEMpXmTfszu2WX5UKN5Mt02HakdOaD+yinD
e3bGXWHwo6RIjpvgjm0ks8xX5fFpfW5oPu/7rWezSHP5Pd3SsMSOhydUomcA8n29vTV4Au/lbgPk
wjiTo6otlTZQe0jicHdEns6H3xHnAzcHDlA+MUFm6VCIkugFzSZbKu3pQDnsYPAQ0h5kd9QDVT8J
WF5LTA7BQQjlHyWcFjar5eg+M4QL0XYEiK9TMal/26PdziyGUjWjS2NSvfqUeZJxM76EMWgwCjq5
xTQf36H7u4sj6jWV/I3rIfig2MUzRlDYJ1MVJfQqmSMnf2bH+dbcx2daCpaZqJXoDX6MbpcNVGhx
IaPFe5i7GLRK01hfRKPD3OBpsGrOLateu5VAxNgfMeg58ys4Zl0Tq/IQclStvSmuA3FoZwgBVm39
pdIscJGv4ZlREPdGnQ9HHIWmbTPjUdVTCWrfHMQsr6r0Y9B0R5REiAv0lZ13+oBQKV7PNdRDF8Bj
KqfXgCZufghesnOWhnqaXLuSH9PUCuNjaufEe53QvYXFZPhjZDn1jsUSsHOPw0yHcizAUI841pHM
KPNbz0y08hBcPjHyJre8vH23+ajo0++qNM8Xz5HmrRCO2v/Ykrwo5dyO//gShFWN2Wd7FTza4yG4
o+BlAAs61y4hc4DI7Vmh4O+WOFR+zQT4ayI56xYfcvQ+vTHMrEhIyVImeRwxv5xJTKL81NYLmia7
fjmUjGTXm21uzldUrNNPMXwJ7oFGPS5KcbTSovxl5ioSPP+A9OwW1RJtVv12+Aoed60liSonPtaX
AcdzKE3YWRchBQRRiq93D4EfnASE2WZDUbSY4LXwx4k5+CxensC7wSo1cNQU4lOhQJeXhrT5GUbR
mFKyQdSPZao6pEs4ieg2068W4b06L0NivKL1FCz9pXDA32eGM7MJrVo2CQMGKSBEgp+SBClTpmua
mc99oTZXapEULCDpiEU6yxXHe+t5/s37eZtNZPrvTqH2CG8/cDSUMXxeXLJEHfud5ZpbmCEPUwjq
Fz6ILR3L5LyzyCNXh/DKYvyd2dieZl0EzYtKS1uw831oD/8nKRJigLM3cDYmY1F9emAeXNyTpbGW
VX3YaP3k2HWBQ4RtUAOD+EldYNYCg80fGaQG7eJ06P8CkzPwMgD3OI+GSRuCs90av4SVZvJLkzXU
FZlGNY5EjdxplSJk5i/iRqC7yLIJrjP037GdWCxCKlzhAKiF/F8cTjWETrN4t39cacs5XAK8R6Tl
GXWxwJQv+cCksgC55NJY8bhA5F6IFECJWYK85/3QrXOX3EJcQo1LDkuH48X1c9dgLA3n6eejnMyd
qLrkiHSrNOf1mp8nT7Fgb/+bVBZNweVMj+Jp3MJXyDXCpeZGv254L17Zwm9Mvh3sLKYfyoI6cMjK
86kMP/TMLtFXucRdZUTca0IM65DZjt0wPvYHOOxS06OzrpMj23RhES/3xYJ7GDH1fI8SeBvPC2lu
eOZ2+3pQ/DbQZJG/7zLHrebFCsx+B8XyDypR8rv/kOuFi9Gr/XVwKujAZ5blofSd7RbYB0tSB1+L
pqCChL6f0VNTQaW6WbAfO6n6Pad1tdNbfDKVE6a/DexkfC0v+8KOjzlMxGHH2LY+l1+DyzRd5wgS
qazYoo8qOwjcSvmKAZ9Y//iSm+zGqoCUUAl7pw3xGUazPZIoVXcwMVPL89yfIs6krPm4JPba+CKj
ZOzSvnUAC0EKLw/DfX6gqvbHoX0WUK0SEJRuulAriX0xS8C4iBKvKQi9qRoHFN2WtEY1nFDKRZYH
U1TxEL7lguMw9SVo8nMsktyQ4kKkmyM6Dfq06JQowp88PaqsDNipnG7ES+ZGts5FUptlRundhTkI
THsbEweZxpOeyvhClxgydFJP26Se32LDPkHQMsNwlw7OBezz3wP2KEgLHVm/lW0KF/VBHD0RlH83
ifkL3our0VsGFsTBCp2el+5XJ3Ud0q3RA4hD+x8DqqrdIXs1V9Y+kTbw7uSyLidxQkHulUgQg/Ir
1zpVoFGC5gmsDv4Bc6Hutd6JLmUiJegXEHebKseVfJl/MW5K2Rszflg0VBWeLSLZVuLK0ohmskcG
n5FaplGig20zeVQWOuVPFEQgZB612+70+yuNZ1oiATZRYJLjkfGYHc3j5SBfSccqYM2Wl6t7D6bV
ajECDLldzhiMdp/2IDa9x5vJVeKvNTrijrLYnkQPDBgsWKFU3IelbzgQ5g13t0w8GSPJ5yjj1oja
mZxKG2WAMi3f/6VklYVKYJFNpdYnHEicM9Y7xs2+M5EvwNrLokkRmHld4b4idchYn/3NCOIHbLnh
vizR+As0gsUls6TQmz8L+p6Gl5vFv6TYt1cyyERVs1+CWEsT9XdnpG/JZKgflCTguIcOlpxetRX4
VPK1aLGaLdBTCWATJRe5bCamyad6lhTtD8t670KoKbTdmkPqnhCMoGw27fHFMOftBSjO8Al/84HE
JB3PjYlHMFkjpnfnISC4iyu0UddQ5pUGZzSseTth9FPflejwZDmn753v3QVq3igh0iXOYZ0pJQ9G
cm2kU1PH9FC/xAUsIf1xJyGZt2xyZzMmjp5xp4NswszTaSg5DVqT+vd4akOpyC1kqAivjYq9LC8m
WTE3NF8omm0VnFRBp9VX5UJIyy9l8qaTUOvE0bULPGHDF12K1Kn1aE4FDlS83EZyJqJo/oT63mEI
q7xv0aLPKyPdVqVK7RnSXgTT05cErGSBM4rQY629H7a57UlOiV5rdmiqIENpTCEXzd1WyC0iDyko
kmBkwVWlkTwzlG7kDe3RFCM5vBgMmchjK8JS/C9a/SJ30xU9wKCPVwUVH4Py4SaW+ilxQgRVYrSr
qQjP14/FiQRvVp+RZJ4qJQmqpi3yWhAWufO2wbt08XmpDUYHv+hdP41ZnQqsFUC3bnxSBad7UuVa
/K+rwCCio1fXeAxIHjuqu4I+HI3rYq6CT8SJUm5ZN/SNAvotWy2b7lZZi6zyT7ATve+iHkrigfEg
kMkVsFPLwEtX847hH5qXJx9cWQXHdAm2aapFtLEPLZcmJunUfYUvQfwA5YwzxFBZWzV4fIKyre5I
y24s6OC8AI6vkDaIUOUzoZvYLv/itXuNGWx6BTt9Nzwk5AtRJQLvx/tATKoj1s0oanl4xOKynyIb
kS/AWTWdv8gVDgRcMdZ1Z2ylYo2CVcnO3g5Pyp8WwzMpC1vUMrlNmg166hCnXD48E2cBoTZ4N/4a
5hkCi7DYdcSlardONA4J5PpVpzEXYiiCHuTfs6YfG81Vt/tcZSvh4hHE/q9VN5RHiIdRDiZ4b09x
IhJNQeKG4FlFFfQV1aLQd75lnD0Z4COQCn3GezuR1Szxf13RBsr1C4QMG6UodYThNTXU98VqIHQi
zWwRwkknE72tOqBIHb7uArGK5DWNX8yRBHaTVJIJZhkIRDUxKYXDA73d3jFmKgzS3TkE2x34rJ1t
NDMfcBIYMuzPRhVayvB43wmIdIfw5GVQn1gbrxxpRP7EB14zsd1ChLR7S8nU3CCLQrhUfNdEyuPJ
jCDDfvfEuuCMmPDuNZGFouyH/awjRYvWvzgKiD/CI5UhSv5mMjbx9vrYaugapvq1zri7X0A4ZRAc
wJAGklD1Q9MikNseVICqmXpteDxDZjHZ0woTMS8vsX3FUpQ2J2WFzrUcE3OmMhaBwpzUFllY7/PA
iY1Hv8zyPVeghYwoFsiEeIZF4WP5qFrfqpXG/2G1wXoHNq6yzXahngQhjicjNbLEXNzS7nzj65iI
jgbMdR0Q/iyTLrikH+76vmR+skMx+GVBGXaYv5Sb7EKu4zEwS1zlCcY/fsLkJmhab2S/gKDGEbMz
fJZKLJVgo3bPMBhrJSZX0f/qS/d+PVguCuzwSNA1vFdDMXJKVMu0j7wL07aGaSWDZJHNujn2PqmS
Sr9LoxaavK1FuQxuBaM0A78J/l1po97HlssOs9k7CKKiInaZf/hKcqwVuSbD1Vea7JXOo9DFnRip
QbXOoZvDryb1LY2XUHeEMhFO5rEEt27olaEdDuW9Ut6X8KKCTkMWlC2irZeQDhwWhmJ8dTl8uwwe
dJF27jQbnmdLsMFdd0lYfpnwk/VGo+R+JgNygbST9F2WALU/IL2U7P9dJjLG6sHLSuU17/4uvmsB
8boYD/yqRi8My4E58zbahGJnz6HQJ/NtfGU/68ya/YaB2hdHuXhJg1kB8eMVpXH/TSAca05q5fJo
f7kb4spg0DSHz70JleMCXZ6NM/iAw+yXyMuDKl+A0m9YgndqYw0wmFj4qMlUUg+8C5P16+4TKMUQ
wH7giuzGFHAcfESufGI+QhxFBiMnGLc/gUUT4/ubsVL1dtkiITahCJr4Z5GBRdTsJCaXPvuMUghw
dWW92EXemaZ8ARUNrbcsR6g5nzKnJ5MLYdFZvdmeauyokREcfT2zfWZnnGKnriEC9SG3HB4X2VkZ
KGZ5FS/4nNnXfGC5lbmLdEIjrxBRWfrSaZsfEyiM9l3+SutdoabDJXsbcK5U0rLSP2a5o/xnMpyH
mhxqta3GuTK11pHe2+k4Pt7jIuWCggkqdqex8E0AQyX/ksAMiBfznz4BK+MPw5ohDadf8cfxL5bL
X5uHiOBbQlGLckDEPtXOZ3BvD90EH5c3PYBNtk2QAy9cpLhLHne7R9qnKRRhHHVLb44wASjqCE/v
6zpz/LfxvuIL8hWoNClhw3jq0aneDz7tIiEPFYGY80BxU5QTMHPpmuVWJpKD4WRQog/r2VLfWsja
QmHHOjesrN5WoFkXPc8h7nvf6QoF+2LFon5PYdneHee26DCC6Vn3gsbcp2xen3/gttc4mPlrY/RK
d39Bld/D/p9/Jqf86ReoLWuctre0NPGwDuxCv79QTkytFkH5Bx0zN1WurWtOKUFY3d0DAvR14riP
aNsaopMRxHSitrZRKzNm+nTqG0ZcDK7IqsT07mCQysOTFgCnTkggBjH0mjD0ejBHJoDpxaOvylIu
rrt+Lwh5h9frY2inko2rfBFZ77HKXdOO0XqNLFm6CMBZKgzAvi3gwvbz6mafRiPjJI365aw/P3Kf
E9IlGUfVu0FqaNFCZuTwI64+1+zAjC+MIvjW876AOb7kghFljJnvR59Xw62gKFsdoGypxCTycLsM
HmPaWdju2IeWcMweD3t0+tSm0XahWhN2oPnRhmwXtbmCt283Ukrt9PUNZ5ZeNgWDyc41S18wU0dr
baxl4SWyIuo6qfEFsbNrFFgpzo4eEsKAf/NtJQeA8rIcSkROOfvYhWAc3IMsTZIzmAcHptc10e7M
0ruWshIPA0Q1UXuLgvKY5Wg1kdqaSk1s0x9ug8USoSbWwdsOGTPd5GPS1KgVtLGX1YZYWS89jhKT
E4We0nkkee11oB2mHCyz0K7I9TeLltpCl2IJeADA741COLpJKOmpHgCa43PWpwIWC/pW7EtVbjHG
TQYO3Vm4d0sEMK5ptoVq0t1RvRmFFE/EIgUeEdeRO5iJG0WFdgHNjqabTahBzaYsNTY1yC3k2za3
Nb9iEgJE4v/x3I8CT6MsvXjlAYw50y6D+LgCYMkIQtQqeHI8/p1nxn8XfT84laSoRg2OjSu8Vdkq
eVQPtcU8Lg6PP4/y1dAJwtagnvwqmH6icbuQTIC5dFjwCS60d7NpauDXbJGr+6YOjEbZ+wjLmjnu
lEleOdxqxRdSmmHDnZKBZl8QASbJz8hrHlAmvKzM5zxBV9cdglLkh5rby5pUQ4cvFGqn5XtTg8ue
T6qzCD4yVGWBiIa1eq4xUKgg8Y4T6lEw1WFQu89XctFppQ9a8JiDY6rQ7nALZ6P99Hbz2FiFHKh/
ODCba5v/0WuilIjqU25YZYHjbjjmev5/hca9k4awCQQPW8bWfQTFix5ZPFvyvEg7flkevQtMBOf3
lkLXw4jrZssJln6HRY7CIQca5wXbOloBCMjm4XtSuWspbaRxyBU9HeKhsYJdlQqar6kqI1MDA/zh
WjTQ317r4i2l8sv7Ks5zkmEUn18b0AlFjZnLipL5RxWSzWlOr+ODOKnQI2MsjnTpL9RnJmCTgJvv
YnpVtvUAyBO9iMZuGZSX1CApqdxYj66uyTpZRhIMgXUEHfK8j8BW41stm1kgG5F7e9spmrZFHOGx
bSHLgmnX0R9ccWoehVTc4cbcnPeIBl64Xu9wXMWZMj8H+L8eGbnsmIJOC0IuNaBGbFVXiaIs86/n
2zCv90euvSnt74xhXwminTWDC+8JXHhRlBtmL7SIz4FrKbXjMH4AK1OkeSfrPWXUOvisnr9jkRfU
c/ZXmDdby0Q67BVWpqUtUoFU9xV308AYATYvU9kGvC25dtR4Ll+nVBd3c/a7idjakxcCDULvIrg6
AqomQBfme3CLnf6uscWIp05o/fesQrZpoHS6dJSqSoWxQ4xKjBmUxDEEnoJluwFbRK+3i9vVdd0t
C/C2HWGD8Ush5AwoAOdx8QaeJNsbCNkkWSeru/s8fKwcbQYpkHQ6VPyMOJgxbQfmBID87Oyfa2gv
AmnJdsEVGnwh3XhROWga16C+aH1B4IuOD+g4S9x/DwZ4BrrY4Qc13yOuK/ozu8/iUAh07QdZRhmT
CyP12VtVjHlXIcDKhI+WSQBxsWb1DzAuj4HR+0V+PjcVZQN01CWIr5ldTRfDeQn9m0xM9mhHvJ5E
0/RyBU+Bl9x7oIep7E6BJe3w2fnsXaPKRadBQffraw2pkA/AGQqIMINBBqG0raYVjNMsXhfZ2VPq
zDYzbzhQcnff7RJYjdupnYbig5CyuvbEfwgMgG75AKyJRoXhQxklxDffr95jwDbD3a+4Ax4Fw6oA
xHMxCmWbacgaG9J0izxfl0L/gTt1rqllgdZCPHKt7wlLJEXiU5nMNsjmB83k9fVUgKh90+/4dH3O
HPfmy5R8YHewQU9a/STZF+AfaAWKWJssmQOPXhPg4d24c85nOQTUY1NN7x09Ikqeb9X2Kvrds8/S
L7AH1BJ4Cf1kDeSuoKeXdJKF+sezJeQlTqONHcgbZWLX1lNkHNKKhUu4T1zqu+1Plamy7iluJluH
nm0AzMmT6BTysp3fyetZ9ym+EaQ+QecT97Ll4b3F9YJvhTPDuqfEVYiNiJ/8hnUPkDQLpH87uiM+
aq/0exnqOh88AdjjKO6Zed9bZVLLeQBtdJC3s8kNDDBLb86ktoQ99OjPMWOVh7v1E6hc1uAtIy/V
o5L9DZ5SATVNkC3mhMr5zftdMWZFMsDbsYAhkKrZ36PxkAKg9OGvI2VT1dbY+C5dRHhxo1+F0UbS
fMHTKYc4R/m+wGlAeQAbarDs+8jqsaZOxk1t5mJG13MqRcuv8ZIWFcu4jhwNfgnapLcmiQ8w51si
+KdIx4SXIbgzuGlzrKrPMirq/7vF4nMawX+xNMAsoFnhLWXI92nxrL38BasKOIStiq7RjfNksAB8
AljAx5BiZFaJczWJJVADONt33ebNm2pI6js9qdMBHHcsXMG4Jqj9vMkdQFQJkjs7xNuF/Iyhg37E
ss1jXXOOys9LPN0prffXPZr0EtWFOa7kGRz/7mG3aY1vKrpaipBxE8zFMJhzRzv66VVtHFiKZUI/
HQx2fVT2iTxs50gLe9xSbMEHey9vZuNHek9bnluvqOXYWlK6YzTTHMYYo1/brE8cHcshwtkHCgfy
lMV3ZxadO5slyznxpllK7iseVD4DXyykDOQisC/hI8aSTZivo2BIwnGUvpmBRPNT5OxS5qQaLpWu
ewGwM+hw0wJsMXguCTdZ+3renRuKFJYYYbIqfK6TCQvb0vu31wiGfCvA9+2tn9TMBgY6D16yzcWX
esuCNd+QDYRU8pngYi9/bBHWO2A20CYJCzT6+EoxKrIUWP/qw/AsjS1gUOq6FIcRtDe2hySPxgKC
2zWfVJM6u3odfii22g/FQMppKCH+d+J7vVGX2OxvNRaLczc2/rKtw+1kArjEwuVH5LGr9QU4vNuo
KCUMw6GGU5bxgOIUE1S3pdeK6xd4BSHPOn9PnGM/vIGzYPIfd2S/hbVobUgj3l7kHa/WQ23LKL3m
FlJuNdGHWpEVQdU7d2T0BLBVPV/52Lic9n8ddWtjUKSX0XBjKD8ra7ir0OzHVNDe7oIOQbrJR+aL
opvdiADl1lJLmoWu/sgyYiic6SkmalOp1GGYEOC0+Hf4lRatoiUsBDcHJOntQ+9xvPuZCN9x+45M
j1F4X7QNDYEOm/GJPRooiq7WvlFqRh97G64ndePyWO82KYuHwvKRoiLwibroXLiv8+dj4oG5aVsK
Dse/3s/eSp9X4XssS9zS9jtZjEVHoVUFe0T8udX+ll9vHnlD/333KN86WG9JU9reAZYL0nu5kn4L
nsAkgvWoONTVRwOU560aT4lUex5ZpdmIkEfBHYV7ZBFDtVmWGt641wiaPdCTAw00NVNRK73qxltU
X8EGv5mJDSnqFpaaor5zM9d23fRrroY5I2BhUF9bDtuN2G7jj2UpkTGBSltuLdMo0XppVJWLdcgW
HnT0whHkvehvJ721CptABayIUmcBUMshwp3YWgl2cfHsEZ8vzUhRHeRbEBfAv13wWkr7xfUqCwdW
/BLoIVtK+wxYfce2vge/MiX89j6NhGhzyWseNv0ZLTqJeeDrX2hThsCUdlSX3stv2P9150K8WptC
nhMlgfJzREjRG/ex3mI2hittiLxUiXpTNkgJVBnZnq219xcwg8/xvVWFCLWzolYys1KEcFJ5DT7h
WRYzemhdqbBHMAgyHoPRR2Z9Bo77gMjRh6WkKFiB8N658zWnV7zt1eAYcgBUFlqb890zSP8u0r4c
avtKwMXHiOjgvvMZSEOdOyVR0+Ryfy7uCbTKopwSzh6o03P20VS94qp0L+HaoPcnox/57jOJUf5U
JpNbNtiOGCHlSux+fhsdtr8g3w8/+QRzJwrd28mr0n6e2H0vvHjFnyJxMbTjoW4Rx1Ulrsw4cjrT
tdVa/m4aNCyifpOto5ADVZo6DTp3TF2ilgyDomTB2YAnZcS+hYBf23jRlYxfTI4hwW1ZQGDfTPDm
dn5B8xNmxtMDOrQFDcszEMZECVyWWLBvTRAbkZ9ghJdYQHETfRWyBV2bJLswQ+EWQbORJbHNHNx5
u0ZFcODq+pnmGb0S5wfQgicS+zMv8F8ayCwxouXqyie/10ZRaIqoG1I6lfnNynW3NjDvPNn6YMx6
3LBho9f+ioSgJn4aVUkIPmrZvER26ECQ1SSj+LfM76iUTTWCJ8ZlKK7D9plf7EKsWRAfVHPNWTt4
n34p4Ac6NAREP5BXIdESCU6iGuqE2PBI4ZpgDHxdlfYwcou+38ySrl7MNaibbMT6viTRjPo17sf+
yquSRJcT43u82yBlECzkn1DmIKzg8RXyHTh3wA8B82j6KsSuFnOXiJcsgKNXpL44LkVuo5QBImQ9
x2aFqrW1tp9NmH9VvaLIWfXS8uGCe3AYLP2Dfjd/C1QszZSvsvnJRdl9mq9rn2K+ov/oLFhFsgx+
+Ll3fPED6rdV6paNNPlspQ1qDCfW9Q8XYrVj93Qw7ojlmH8r9Fzu1DcR2onZu7pa9knGJCTPKReV
EFcakLFD+NS6gS1q8wQMHuN/BzipCXh8680dyhw0HemnI3JYAvwz8T0u2OeSTlY+WOwMqc+xEvOd
/h1qSNhctZjpPpsdJOv8zGSil7IEYzpr/2ULGOuAcUju/a5c4y4uf7bYDeqOp9jHKQDzk4TgAFG6
RTrIlgLx7jLjBjMejowRGGwfbp10qtfsbJTUVvEtLE+SEv++tBmjQozNNwikPZ0kuUABNxDQYjGd
Ks0/K7yZ14J3N4LhPcKU9sF8D7ACWh1HYmLL2A3emVyj7/Fn7pV4LC7kkWYeh9AAFz2omzYZpz21
T5SwyIb0YNsi1qmG9TMiLrD5aswzCnNZgPxPIVHIkBqxgwLOZNS83xby79hy0hIGsXUWR2AU65aC
ugLpXcdaQnvk5CTyKVchfZXgIXY5Li0kQc2K8T+G4Wk9HdfU9KHPsfGgYbS8MRFuUPpqZj6rlwws
+pNdbOt8J5AexjVxdknF1ufbt5c00vAQZDEh8zLsOqmQYMRl7V5ZYsP8Qfceg0Fez58KPWhHpbHY
bE4RPDD16cwaTfYi/eLDsV20xpXS/pcpUAEGtIuxcJE3VIr2NRtE+8o6FMbs5Zp/6hqOfnxkXq/j
mYAnZfEtZc/aUNkxwso7f6DaBrF13y1HE9wiU6AYH3TQCxTLH6bZ2KGBbEfo0JBZjTVJgqeQL+sl
K0G+tZbnMxcaZfWSsb7PPJnxpzu+vYxghJ/SoU77yXrL9qOP2uAlNI0t4vc3/CDO3aT8QsIeH91a
NA4Jaq6652kLANlw5I4Vh/NwHA6Ph81lmNT8mObr2JGsq9YYQ5qjHdgGk7/17dLLeFAQQm7Crdqw
aLCC22Zzh6KXA0/E+bzReU8fhcD3v7DT0MTeD4opoTjw1KbOonMAgEtVn0F5VYnUuVXwz2ermp6X
sHxEo17Uml+B9g2m4673I5qWEPbG5VR5zLkUcK+E07aXeDAhxPpb2YN+cOGVsB0j0AuA53OSTTjg
6yw9SCgAP9crr+dp/Z+l38Qq2+VJNRDx2fmcr/BhK2+/hIztHaFbbH00UWOXiqyBR9pSE7BQ3OJW
x3k+QouGFl/vK7OYmpIgp7gQA7T5UM1cM/X0dUsUJC51/FcvxiQiG34ptTauBlEuFWNDxL2U4gjm
b00iGuSLf0zh4iaj6XWOSLopS/T4lavon96Qu1ACPyr2gaPMb3DsfnR3pN+rSVNwrD8EGjm2vLiX
u5lX4DNszZdqNdAEd7v1UxB1yAOJB1NAU3d5cHw/8syql91vHEDd8WRxBjEgmWuMOk+5V9S52lEC
RjmQw5ihGax5brsUR+ip9cQIqIZcCrB+hcsSuyLndoPm7thOU71XW6dUj/snpzNqwnnjFUF5lA+/
jwNH2162k5HUlbNSRBjcpK5JpcwOC97E2riFNWC49tW3/g+al4gPoGiDw+dYoBuwHH2r/xWcVNR/
SStDqdPA6ejYGb+ySr1EcB5SFqLPKUZc407J3Gx1I2TcLE7144of4ijg5PIJ9AIFOV21gi/ONWEI
smezSanVkSGbgH7zci0Oe7oO8oZWIqNjVHayRBT6kTi4aYUU5kqdG9QtoEkuQXs0bEy0T9emzfJJ
wSvDWg1HUGT/eGRRxh4pmJ/ws+szBCM/DADWf7uFAodigCyJpehLJK2G8Q+KtlL5Up4mjOdIkzXV
jcuwvWEcJ16x8UK4F5PlAjoDKlst+Umepuz6pbK4UWGFNNLu8tYXRpnE+pdakvAf2zz7S9+B4HWw
95Cwz95HYCSWRZOCiWLT4KwL1A0oEPKk2S1VLvWll7bo7KU+4EbqGLG1lkyjR/AEoGoOqj6cal6B
HW1pGZs4Ju7CkYKKdmil4b0XUMeI3kwh3ZBTbNd64GjJ0p9yM2OFFjoPgp4QHQE7qenYZ5aueEg6
QsCnSAPS4BBq8zXoCcCIpY7Pb54H48nwATTFjNzR8+FzTE0nX5+SKwvIzKl/l+0E8AN6VYKuyrj+
KHjkWu5fEX+2S3BXbANH6YN2vyTYnZ617i1mwmxkEUsjnvEqnXuAvkACfJkBGkUzc9xH7VJHvMw4
CURsOO8nHIIRqcEsfiY5ouB1YauAAWK/EA4QE0SeRXtiCSaHrvTRNSYyXw/cDJjiJDCaTRTZ5p4M
elmMTdh80oDp5bEiD3Wem3E/Qqc+LadsWAwoHutxqvIZYISOU9JQ1wI1GdRiuE2YBJRQAp9YMdQW
DnQpk7ZjuBCQh/SkDBLFZKPHNGVRPQ+ZONYnIZZ3sE/NWT+N/OOeFy5n7j0b6pvG9PMcTrLOEyip
4X51aeHLesMEK1rJBNyxYxLy+qGGvZeEfNHBzGZwZZRWFpK0IJllIR7JsZ9X1gbXbMUAle03eFvG
Yoid0Tzs7IKnp9c/A0ly5/jyaF9Hg2/wdFD+xQJW2VO3beXDy4qEUbs0C6ngJjQhvftNgRvr4w0T
k+5Od5CDQHAGJJQcd1J8FWHx7TgXsS1a0vtAJoP/WyzjHuPKasbPFaaZtrX+NS5azpccyJYI6eX8
sQfb+Ph0EXnHzYi4c5ul6hJUiupWKYicPG6CSM8iDVnWsWobsYzGBoRxgdfp21tR1dW5JC3UZXqW
lsHZrYbS5nAL13l7QobgS2bI3BgXo2D7a0fOxFvnYtn4iuQNmifW7Fdhkfm2xlxQ1EwcdsrDiMHH
eI8kTJqiaXRmb9sg89XDz6CwW9G8WhrqF7nGqrxPt8SjACxTmh10J7M18Zai44PEWxvgH0p8Y3m4
8pXY4G26jqpQmdN1KkkAv3NWfBwfgh4Wyt/mlDVXVcWRDp0Zsz62IVHaIL7kPibnWgsn6jzFdfNk
wZObXKInl3UqtRcAx+9WsA0582rh2ZCa8ZrnwMq1oszN5wfjGHPzfkEXJXbygm78HnDN3vUxt0db
B6aveYJJmbGD3WTEBj/0cNgsjDQUedRscVJMklwoc2aJdZ1TK6vQWoUOcjsijUXgirGbNgMl3iUT
sBngGytbEIN4CD0o+7Y69Glpd1spAXWD/G4bvjGTkwM77RmJLB1wJieW8+y6x0+OjpeEC1XG+FSO
gmi5Awq2RS9jIA2j0BKCoKU2rZ6NtyMvkbvHcdnf2V1a1Kh08PE6T57mF8QWK4az/YYIgDaqpeBM
AWGfWoUMpMvk+dmn732Us1cFSD+3Ze+CPopsrbJkSKLN5MuqJZ61NitbrVO0tEB6CXb5QKUsrmlF
jC0wRpRqe+SoFcm9+PfTJyHbCGiAc9mu85kp+eGPUgHEEwF0iuqDcY6ATOunab9d7xBKQtgmLhT/
dSqZ9SYPnwZq3tonjqF18Kz+697l+Ta7Vz1DlGgjHLySb63yreeq9e9TnreC7LXLcQzyb0K0hIJp
0FQa9dyBbD5M2M3ypxy2ve96GTftHRZkmKnDTus2d1TUvQ/6tbCyUG0oyfQAy8AEJzjVczge0QD6
kVBAA3Oev1+e6VtGgSatk/+NYvazWMe1/aIWkBLsWXsLRZ4BrJUJDGsXhIlrzcNarTRoITvxhshL
ujSnjcJ8pwSf1uBWllSLicUPOaHfyE9w09cN32fhGkUf+tNtTIKxtp6SnWPsHTPMWbOJY/0rmKuz
Ic4AVs9oamQsb2DITUBsCQGXkFYQexZQf8S7JGqBcjFlvyz95+T93JyIQEcrR00NnAtvh5Kiy0+s
3TcrLWt4RTu4ou1BrkN/NrJ/DNMVAIXVuZ0Z4rTUPnDmXjH+5EKIq1SR2vZSRJmzn6MulfXcKYvo
1Ptgh6kjlqLOvoVBvs+pjJqtAB6a8jtxa08F1fUBQ2Rzy4TFahzelLPRLPLMgaf8SkhArrGh4Uie
Of+EQTjv9TmN7ZE69WVFUOnHxGS6sp6+6tEOzEGnwQH3I5z4B1lpPBtFkotrDNnsfXRQv5bXTqKm
d4QIkmVVct4wvJhruDPKF7JhXfXvEYOdMvN3fseEMkgyaavFQm6BP6JuicJHXVGd/735YWhx5r6s
BuqHoQf8OlrvUmA0LVSB3zw6YhqNcct+RQ4t5hB/IMOVBBLK0t+nHW0f15HLk+uFhNpW6AGj2qmU
KPWX88S7eZwzCJ8ez5vcdd5js2VlJvl1a9KR5ooj5k6n1slh7Nm7B260CJJcuR3tU3XlDbGJ/mMa
Fp4h9wCg5Yh9RzcSJaUh/5lKCMxF5MZEgBBrRInaPMkjMMVtnmteczTfxjeZa12znuLpSPh/VPXi
bDtUTESiZA1CMPFFzvPWWnm/8ZsgEfScU15fO2kpwRcaXDcLrbrxfTX+hr56ynpwtf2goe7FABk/
+yAVwPo0Vo2J+XfBc6WZWyVldQ05Dr4U6jLGYEzeGPjxalhjBPU5mSorlN1OfBcjCGxaAs40bWk4
JTXbrSs1KD4Uc7+7klOnBBWvXozIqs7aeo7EYP+nnPGOb+cs9uIrOGKYq+YDAld6+R4KLg8xhREj
t28xuFnEdmfrh2+YxXz8zbpT8l8R8bo5iDjQ+rxaG8M9bdNWb4QIZxibiskpIv/4UWdLoX1r4D6w
SKGNDh4fUeBrDtVXNxnCDI5PjSak82Xj/pm7SdGDs/u9Pn0HegYuYXQZaNHoFtScC4WbDuZu3gEA
YKXD73M4nSXnKOZHFh2cEP0+TeJMBSvYd74faFShcQZMaYld+O4hUjKAF5/AZPB+0zsm8gFbMXJP
AvZT9JdFUdLzvcR3Mg4VPTq/w5BYM5sBQ6YULdzeq0Tk6/AnCIXOR18345AyBy3yj14p1FwVsz3W
n3GcdoxJtuZSjf5vc94k2AHdGzJn2SaFkfmjKc+m4BbAy5ZnKTbYGsrx3Erw8fopP19keF6EliFr
K3n/YtlbulyglgEkr4/vXxIz1C+uuc/I5LczCw+jRzq2TDFRBRboEuDMjJlGsnsZ6iI5ysK8AU3T
y41WJHf1SCg3WCSJXR5I1iSDv51CDkp5Vkun4mbar9HaFAQp/9ohr6AhxMF6SScm8VfTf7A6iu2c
Ij09biqL0Y9VazTK9LPqBTMVCDpUrjBupxtmoyCdD8RcqcUKNtbhP8vxOMQfl8NyRFwxyChvrFz7
1eUwAgfYoXqkU9NwGhOnYemuWJxbjTQPDItoIkNI8UfmOl2adL2DPdPRL4WrF8EVHIqZLIllhx2Z
4YPPAiGqnRY2h2TwBq0rG2X0ogzxsATJSnLWhzNdlEWYUk+gIKim1QJUMfCGdfRkEdnenfIuFVsC
uhpX7UWl42Pt8+51NLYi75s3CRzfwucvHkskc7SPkY0vvBo54ON9Me8kjL2tmjpnonwOJ2VTAxfn
fTPRkKv4+BuyskyBJfM/O+BeCl39bVKjqo4GL6AZxJrXT49Zp/vPYWTnVl9Mw3+rFNmnhTtRy/he
4zgCkJ7L6NWwaVluYandg8xosAmcIa/zW/2aDSbKvoXhcF3mhjJWFGaKWcdAyxp8gZ1popMpJszi
ziWgcCiAQ+rwPu3Klzmbu0vGV2wFgtB0lPuoTFGNR3hb3DIpSgs3iL42YaADNvWPtVtR6Ub9VBk5
JJo59ebvGdibMR3dLQAIMlLjxnhN0xkJLFuIEP8rnqpwpMQFdqPIhsUpdmscRrb4Qu9ECNYBFPJK
BjxRLyEAEd0IQdjP5mbNUg8gA5wTk87+nCErWRKMxod/oOcd7K0WXroL9wwlCH++p+h8nSQUGxZV
a345sR0FP5LOceBROeBQBzQ6NAmBTPjyqttft+5mrXZKIHiOQMg/V6iNLBt5PCfhZyd3Im5WKh+/
eWh5VsxehzlDxKcoR+hPumf1AZAYbrH9FelPfPVafIdIrGdLqtI+MAI76VIasErypusdKz3fYVx9
L+ctwQjSaAgzTdzSwMgWPxEOwScJwbe7T11Ii02sw24tIfJX+wg1z7gUwN4O0XKYA89Omg37K6Ye
JxFKvgECdv4r7pINAfB0tBH2WgBG65rjkvBBG4WgaaFZJ6EnNdKR6PLrXt8XIr2O5yqjx98MLi30
cVz013tOIbPz6245t1REUcXF4C1sfzimpYXjPXibwateqtg/25bTOBNAKNMf0c8vWJETAXQOVGRF
V5X/d95bdQr79PUBjN+3md1EuiKeuup6vn7mUGvTBQ99v+l+qjNBJ57qXqGNPsgLe6qR7M1c4Htz
gLX0dZFyRbSQ8HdsO2+utUYddQLPAkOVwotteDfxTc+ttmj0R3OBwRkaLUgRcE/sEq0WaGpE8mm0
KccsQLwaCaH5GiGWGNXsqkN5orcHpiZBGFa3Q9dH7KzY3c00TyyVsGFFWancHTJ9NXbb9J00boOB
qgktfCGd6b5ROut8goxt2817et6cOZNHx14ZsjLAxRD4lsgUJgLNbKmigmEVF05+aJyOueIqXIOp
093r2YoWgAzRA24PUCUBM3ZYA1q4+1p4Esg2hxIrjdrnaOCj18rB5wufKyJNOouGtoJNeUhmNLwT
dcPpwUvwhJTfhSq7hIARNxUn6WOVRwIy7iiUd2fcpCeoh6NwBtnhhjGy+oi30xLePeYkFJ2EDLR/
aicm75VRPo38lPSaSHHwpvUQKh3Acng+ashLZMdIXNbUfF5lSarAgtmnRwDyNVFEglJ9HuObaqDF
4993sRo5EsBpJuHY0vsi/JPcJ8077ht9fXFaLoKTfTxGhe/hBQIU2bGzsnuv8kiOhE0ECUGveU8n
I7wGoNdUDcV8gUBWmMa/LpmU3cKoHNYwkWSMxmfdtSGEAsE6ofSYO3ec4Bv2OAKv7sWPPdKiNJM6
iPie/+Lpy7rcSXeYIBZxCMr20ggs1tWB+GInfOhaKwyjC6VCvUIXAQr+ySwfk3KJGxK/h8nBFXHv
byQ0cI406gqcmmaZt2shKZLKRaHK73yJixW7Entj9OzQLMTOvtV9RsNqGmDPNsUjNEj0/kiSvvgS
qXUVmp2AcF6+u2TYnorlPMsEuPjY8//xnyqPFx+f0HZCJRXN0d15mS5WrhHfnKg5QmBRj4QQuapn
Y1eE9hnJMkr+uq2wLoj+8JaENedyBsHLKtEioaCfy+I3xr5RBX8C0UbL8b25fXrXguaZ77Ku/kSz
kpY2AVZrQumUMo0rB6+nSGJkALl7tBO/uUMWoxLK4xiP6Oiuoms1t9Mx83pn2SVNjR/yZbuW4Ya8
ZZdo6zAvXaiU6IWGgqaAGgCQtCNv9YsI/a6H9r+TQrYhcZktOAK9f2tXaFaDsEQ6VYiorUKBo4wl
uyfkb+tugfPkEm+I73a+7tFlTQKM7eBsxiupQTYRIbnFChMbJi639Gpy0kPxL7r2s/eLrNaJnBVY
tlL4NZE0nn4g3Bgs+7JqT1Bpb4wZr3QoFPX1lG4GkbSpnw4VOHYtBhjFwA+fAF7Xj/5WclDnob1N
clb7CTpr4PjB2/JN39/Wl1t4Lc1E8W8ELV+iv805/BkZ7OGLxuVle5ojkC0Gvjup8oDQ83ygA2OS
2335Bu43O1idcI1odLPNDLxnjLsjQLhydZbaGgc0tkvDql9AE/Pqg+k3rgTy5FSZdlmDqGH4uf3n
OgYFc3Y+nSi0+HNkDAsFqcDWm/2QsyA7gpBl9iuRuLriUnRJ35prMuBnCzjcqun1THEXHIO4qMOJ
cq4ZTFeILYfEwYTfy69Fw+O0EdTh8O5H9EBcFX4Zp/eFXrDG3xxkSlrYdVhNEs7m7Ra+02ImYTaP
WjRQQTfR7crFMXOuYdfQvV0g5hpOTnqU7IgmoDnNgRuexWHuJaUeMYbM3xpilM8LS6hsYbzAhhRJ
GDoFyT9mYpKStPFNf3kaFJO3eSF0P2yH8Vc+Oligk7Z81AnLmVNHhN2TO/yOKZrYmY5KDFi2o5DF
QeN6nnZoxgxBqu9YfL3BeiGMNRdTH59g+HR1Ub4mZqL3Si8HGySZiwmUroqC5ZAE7JZNIt+Ev2/x
GH7Dq+C6/tNUfEN4GHuEGlZkwB8dRnju91T4Lgq62lsRSKctCMSeJhZSRLDCPLm29IdPR2nQ+SeB
C0vv49TjviwR/oKpHhcPLuC9KatrWLjfADDYQK1d2lB9ksHo8FBPt5q+BYSKYnOT9e8ClQw2QhvV
gfFnNJTqCzJBX/XWy8cPpccv6apKAUI70+mpX06gLBL9B3osibViUVsJJ9BdE9iY+J6GUKhk9S+3
M5VHY8TfK15aufS6pCJTD9x1KqtYmBT/3pizeJK/z/Vf/nTaTr1hYTGaVqegHJsYvKDi/Jl++qVr
xRmmxYn2zkYw+vRc5eUiP6dbMfe8kwDE0Tz2pz01RxlxkPxtSeK0RgKGUmNc510Tqwf7Zf9X6Pkl
3G/WbfGCSmLzbcqh8b81KUHOIBnqRTjaF5Q30/3HEY8CISBiBUBQgshjk1/RsvUuZq9Z+isN2ogx
hXm8lMrDQWAKtoHfE4f5502tJoqIUartzzTw/DpZDGL5FooEa3AzWgcqMfI/WUOPL0NyTtnFXzI8
OvZbHgu6so8W8Go6sxS6UqB5dTsz+nSoktRsOCMk9ERq9xK54wTdPzIAu4lofWbMwy76SypbqVfp
Ij4kzOX+XRM1VuueECIFiqMhzwuxA8j/AlFs1zG9STfxYUNobgeZdSucTtwaSFXhA3EcTccE8RYW
HhzSR9XV+84gJX5S8mtQyDB9gc+ypkjMIzaXMnkegviW6F52ReImCFgioTYxrFEJtBGh8G6OkRYw
A6h4Snv3CQyM8wVomI/K0bjDYEiBZ+/3h9UwWswieym5uqL3PFjwOlPvi9qFhb1FHgB0ejkmEtsw
mWgnqVkvOGvMn46tdy2GX2rU/9VaFBWxbX4P7GWxCOjeHun7NLN+Ojkr6LClZE5RKq5L2c2uRx/R
vEHQ2Xh+jASo8V6eELIWyOH/yvd1QaAnuerzo8wm0ftqkW+M5o/JvLBoCoytHsPuufeUtr6yewxb
UAZBq7hVKY5I8pkjOvteCENJB2huEMQjJvOAdjzqUcJ+8dp+AqwQZPkmPvu5VO9IG2jCPfkvTNNu
HiXUhGjIG98NVhEyr7U+Cukpnuwnalci4cLMQ6/ku3R2dxasOtapju6CZIbBG5D9Exeor1NrBBUn
ljkwiFqSeKK/A8n3mmDLXm/N8r1ZpvzwpKBLek4k4AJ4bHC3LROLSFFjlzSldWwO1xTyL4nJmZw0
hYO8DBDbwmSb3cp5mJ1ApJVgugqo6VlHO+YjV6DBE5dJ4bilqqwCLT7R4KDPSNKJqrWZXHQGRta7
pFOVkbWGHSm8uXpxO4qgbt/IiuZue+Jwnpohmw62ITB/5bW9wP4sM3x+3omglf5TvlEA21s+mshK
HbGgJQGmvMuyrIP1lIDclbQqIpixBIXaiYDllIo6oHnCOnUlYGQv5dQY/tE7o4uL2gLWnB8CHfnt
3c5AQhM2A40+6n2rU9u6uKTkvAgeXHFrd3POWpP5CMqxsd+wUqhV8rMupGjaxpFAAPVZxfg1u8Bj
8ewL5ULkmW9cguyYxIyImPvRhaNuXnD1N6yo5oxoapwcwNjLOAInUHxJxVrelCXWF9WrAPDmf0j3
DDqfG4Am+Q4jGZWrCgsEHYvzVT2vhaC642LvzTeLRaO5UGiuWnwMxs/Ec0GRDvtb/2vzskwNdNad
0P8XttiWQ3U4BHFQ6NaptXKMWc1/KXwuNJW5p10FjwThr3SimDylhh9hQNDomeF4FxZl07k/z8dh
kW6y3M2K3/X2RXsL5cdW2qkB/ViTbEUg4DZDYF0y2JeyxYVpO3p/uTWMtRFe3omUdzna8nSr/buf
gWGp3ZCtqbCD2uZQxlyb9g7kY2g+Y81cu2BKLlKRniy93XkfoOP+19QjdFnG93lLv64JBrzmiUGj
gb7nmYHa2CJa3NNovTBELXJ+Iz4wIoaTHoahuga6qTxn7HV2Wgg6ykRCFFeV+6fWjU2A2qe1azQA
RMC/+3OUfuVTyTLKjlZwv4jNpvMa177tiS6G9maVlRoA7xUTVYLRc3cmCem06BA8njpAmOLYh/9Y
0nqcCrFs0mY7DWhuZKbctKSdMitkvrNoEm5R4zewhqCrLnswM3T5W38JWV8l85k/SSNbaCQpOrnn
lAioUaxaB6Xjlkb940deLV3eA2uLHoEwSqRXpF4QYNg2DfmUK1KNNJAjkMn3aEYAuw313CvRcKqq
tXTwPy3NRx3qKaAaMN2e9gT54G14NRMApiSPsGMbF5JZXB1JlWPB2IByVU7o5Q0G6rvXLlOBBZ+3
ACr4U7byV1kZarJT44MYM2DsgF+yIPXCCVqZNmciPH5xBBPSY4adXvUFYUK+hMusa4fVzf2mjo5H
+JlXts4kxbyxBl4sUXmn1bFQHirmX8UawkNta0xNUIU+jTGsp6WhsSoJvpNrBKx1AhysCSUOq1R4
RsYQOzAn8eacmGw3L7hlol/R04WerLBZbD5OnggreMq0iVLvGoRs0YA+BJkqYsmf3WwQoirD4V4X
btO7jKPx98KJi1YC0ZuZ7XVEUtqCz8i+9Hw0BIEbJBURnS3VhPujlv9y2dphAOrFqrKPZFOefr6/
u2Hswy2+hFjby+BLtywBFQVX8AC+xVYv1IQXEPZ5N3CnsIbwT5AiaEqk3N/m/KgjSBKe2AyjXe9h
+jXsCkaj/Hse6maG2KLkz0emkoC3hg8qKlklYVouVIavAeiIBFEHzE7afcl0OUQ90OvvXFgMZeF/
uLpWayGc+/qbwJB5T8O922p585Y+qKAlQuQdqW2E6Q2fvHNBUhysRnjwil7zvdDogWMR8lIvqAMK
Amitxn8wZHvN5b9zN1NopeR1kPv6UfJ9sEK0xnwr5gCN9s34BtGTU229lQ+Ax5x/ZZiuBQQax9qY
TgQcqrDJQlLxEWnPW3wElVOOAsXdg/NnMBYx3Yho6bgbaEmAC8dBk2TMwE6ULR332j7T7pBqXft9
tG82CnJqBDDKnVVUq37RLZGg82bPQd9hTaSFbhI8J35OOTBq6p1+Td35BFtCybecreuQ76g2djeB
DQ3kWbRAbsCydGY46SRziU6oYiWzU7ZrLlpttETIsFQFvf8gc5k7PrHp4W19LQf2KRAQjvBmTiem
lCaPnB0no65Dr180NJkQijNwEt8JgjDfh/QNEuD0cRIdYLIAnE6+Zpmcv0mLWOGS0qm1yMazNlKc
BjdU/df9GAx6c5YXLqv6GmUmrlFCwK3b4/+yo7cCLLmezI5k9Wqfki8hHqMle9NCdFfiz9Tq9j2R
97KW2aQiWnm5VtyyqTcWTcSvOT7UZQsnxo2wDKGA/fLuUYNVNjWLNnz4RAGQspCd9IM0vCR+BVwi
b34oNix+15TilTJmlEN6n65imvsNiMatbh/4+QcfiK1u4CewxlmVbJVY1vo6hn3Xg1CS6fYLXbOK
CiKOF92sBFwEKoU9xS782AonRtx+VBzpDkE5TSFp6zgDCeoBXOSRo8Yu157L/vnE3u78inHVBYlO
ZE3yoZQc4jiMrcLRY9gD9wbNRhy8BSYafR+jN86KRYzwWsawN2/fBXaJg1P9Xd0bZXQcubHTkNd3
y0K/qP+MZZ4K9LvibHkJrdaCCQXB44umsl6pCiLNdEbqlsGMG3bYiF/HA46yAS7lkm/4Cm1Ge9Hy
FVYVd92lVwbOKDhabLvjPdh8mbz79cmQwv1OX1SLV9coGd7cyJGvsG87QexdGHsgOhgSZw5fRGzN
q8dQ2hwI9U6/3v9lx/b2dgevHmnoi/ga7HS0KKoT0AUc6fXovzXuOhrfTHA0VDEYtb52mhWl5VF0
9Kl08HCXDYvoE3tEM7sArxKysJEYpbAXKHtrLpr3RyYLCHToCO34W5FiZ6AhuFhJb5+jNBrkcSvr
XM6vz1MQerwQJbhXFBI5LXa4I5BPsjZOoO3/ITmuFYjAmZLjHidRvWM23JD7frVec2Jjas63vdrd
VZ81Qhk+P0nl4F+pP/qDI6MT+JptwItwrUb2jL865Dg4XFw3ulZWtu5woqzvx+JdeVU2ihJGYK6P
DZqTlzg6/LmfFsOx9HSVkwwZCXdxLtTGKmM5+DZm+RTkwAsBXhR92L8CPOdfvbB1Q588S8mxWnyY
97VMk1rUVslEsCj6hUdgWhX+LqT/G832YyCOww5Z0x0pRJQMh9GRs8qsTm2eqhkU8vSoWwiRxgjF
e5j66yREu8b1VA4LPCSPGMKdh8IAxpLNS589r4PCLJtYBgnrhQ3lQ08u06Szs3e+2SvpZ4sHjuMz
dJiees+/MCQtNoxEGlzVvxq+ZXMKCPilNowdcaRBhKz4GsWkHSkRaEuxBa6k4oICFTVmRAddI1/5
uZb1aUsKLjT0qxutXONZcyia25tQ2Vq75YTxo5Wdh3ZNF2Bp4zrdMy9dR6SmHqdUUKO3euQXCuig
8VY3o3RVvWB7doavvsCTieuN1W/SmAoDhGf5JMzUkSD7/egtNSOSTJ47L2bGHjcx0eiwtx6PkxQS
0A/WpSLHNYV6dVUoxU1VCqK2mjyu64Oxiv61YF0sbUamcvQ9b5jANbCCRfb6Gn4svoPhYX0qfYD2
d5UQnDyuuMqengidoFF69ND8t6hedmMjwiuotDCj6eOkdbbXEZXBs49uFP58fwcm9iWdszxqdU55
id3lnH/cCdmRWnCDkeyAYyWjZd6VlLILOXsKRz6Uryjcg0xFMN5soZhN0V71EPTTiW3o/E8BVMtN
4XOAiQZAXMl2mYEDPG1sXMm4la3EbHpnXG5xQQgkI2S7YekfiVW4EBEOJI2wBt/jrCkgJ4l5pKEx
PYpSarOCDw0+Q/hLrz+A0CGh2CK04MhOKoeY/9tHRPmDOJrosPPJVNsTWi42oQnhVa37GwZbtR8z
HbN3kqC6UkznxgOGFMudpE2+/Pzm/dSJINzzuwAvLQi8IfTZb/LUGknaBA+g6Q2czZFL9zXwBojf
8orqvmaszCphpPkOPwxP0O/pvvn+lkG7u/JrzfI7dxsVRzxNhkcsvfI2KGR/ra/hTBfkWFbGv6Kw
quautGgfVoRrSZfuLiVVE+8u9QQmeDEuvN2Xrsud8yJN2W04004NIfQ9C3lmVdlPhd8KlbvRGijk
z9PjhGDZ+XFINU3wpAOGX3kIHeOyVLguxdtwkRllSHmrVVgKNAK2acgvb04KRcxH8IYNyCk6eL3h
elRH2s9U3AJSrlxOnpcVzIV5T3QlKsB2/akl3qyt7rLXAtvC4+QnHSbFom+o/MT4TUJ/O339XQhi
p8dI2CkYoq9/b0MOULGOSnMWwyjz1maY3KqPWlkQH+f+cus39SU+/CoKuAcchvfndhqYorR50aTW
mrrSlgQRNH1dNM1q/NU4JkjRgXZc8pK5fbaVBfNOv4rGiC+8ehUhrBaocM7rp8JiEgNZD+WL6ADd
H1wmjQkBqqJ51XTwlOGPk+Afqo/mN5nTCaXUnRKejkjDZ1H5QkHEuUkTC9nePVjSKwRLn4hc0ycX
SP+INtz8axcM5R7dxyRwz6nPU4P0240wcBTvBrlMOrCXgZec7r0NdOPMqV33ky8uN6INHds9uFsS
ry+FkvWQD89DB4GfOEnBXFJnSXS4oDPrQLOOMVyv2wSFgIikGl2T9Amlld9qrGe7gsf13svNXB/Z
vH20CWS8uL8u4I8Jpc50SkAXqKPFfnalI8I8feNBt2+fAurSkqJxw2WudIgZiKNV0gVEuEhWbzDS
ZCxa2xV/KxAkESo/Mt9nYD9Uqmk78cFqO7LwBAWJZWyAdM5Ez9vXcJ7hzGCD5cyER4F4N1cMVrrP
gdyuLInRFbh6I2tyR59tv9zvEOjSb2rr93t7w2HZ24jPk7CJ9iPEjToFwSfjHTF2f6v1lqvrxF0Q
e0ZBCs3AV3Pqc2O3a0ibdMmH8KHgDbhUQ99cCtThVwvo/jbn7edHWfi2u+bpE8UsCdZ3J+JlARt0
cgtv76VXCP5+sNIE/+USMTVXFye1hObHRjH3NIJTbQNbDvg7IFGYtI9/3wu/REoE2jvAIySAhRCv
eMiJk98h/sofUnEctVgxDOhv5B9cx4u0yUqTuM18Kml7KDP5e6AnthYR5pTD3FLaU0pr2CnlAtpo
7vgaV2zGhbgKT58Mxy4ccYU0hu8Ns5hR8JUFsrhR/ZuPTDAQkkE2AKgZqVj91Dc0Uj2wNZc1Rovx
300zmI4u7FypSi/NQe0Zm9AZ+EtQ00TlaQGd9hIlqVf2JGZ43+xY4Pec27KzxvJAw1CSfMsKxa4o
7B9NbESkGAmlOaCZjp+CJrmgitP/NCyBxZ9Ii0XjTnsSEk/noaNkPO70eoW43NuTLg8XaxPEg0dA
g28XoLw6752CFq2lrnZ7t61GHbgs4JcjbjfI309F+gJjnh062ZcBQfmGHDjzGPYzqBRp0SYIwIOe
WY3gLDdGESBgICZHJt8Kj1EMBF+x1+v57+ZbMlZ+41ROF52Lz8Osw/17xsqmwmJMzH50ZH/oo1Hc
Qcmwv9UzWGWBd5KChSuTBvtHJ+lIvlk/zclelRYYOzlinCoQPRhTOu1XrP04q2kzmtOq7w8yzLZI
e8Nn5fiNw9MnTEgHMXA8TSdHmtnHOLWRW1c26OjVU1oRelgkKQlJfqkr2cuxcoEl0TtKUvSyGy7E
ixtm0+hZaUKVfGmwkm+ohy246JYK2FAQBM4NYoukXU405BEzDSbR1GB+yS5XKUCnNy1yfu/mwdqK
2IyN/ORnGsIX/tAjYEAa4temfgCh7lGlY4SAtuNYzmKYQbLsa0bWBBD5IsSsP7jBSABurHIjBs9o
o5FRQiUXaDDFUs9rLYmu6aeUwOHAe8a0WH1LjPj/8mAqxNOyAAeDmHyc6Gm8A3qmolOKJEPUhFcJ
+/wq0SNrBPEE0DfJx0J6m+zHrNon1xFfP24ontQtPGLAIeLomkwhToJwRV/7DILw9uGTPpCf3pzB
LPoqBhA/elaQrFbp0QhQiu+0bYeUgDqugXqWsNangEPFabTdzmduW74K6PpiI1j8HdwfGHJHZdhn
hynycBo/SxebEmYgaiF7UTWVKlCdKrz7fZL0POZTO+4CVUDVspRvStPw3+ZvyDc1UKmpCrs4mAsL
I1xDS4EPke+yFJ4PDKlNj2Qrhx4//JEyt2lXs91FGriIXuao1ypxWWpvA/NqF+hWtvxej+LBFMDK
fIW9FKh3E6FAYFzMtZFKF1tRSxWjgJGKAOXTelyK19JYRFiKbQQX9zz/7J4tLuVcFzwXDSZB5DiU
nEJWvDDgTF6nIBw/7rR5KwgkNaSbHcotQHsE+SVf2wT32BvtkDwT9UoCdZTb3yyWcT+n8BRW+X3J
opCKXoPDktMTcwr0HGESv5IGKc1Eq0lu1THM1XBmBVozl4693YzXBhCkyzM1o1oSIQYL+TNZ6N2t
wNUPGYUbeT0CHxX3XvDRdDPjp/OG3FjD31+3TeR0UDtkZzAuGCfYC2qq7VRXCcaMS61QAl7YFiZ3
J7dpb/g4BqC45feAfBWoulj2Y+NnygQyJ+UTRkjHq4HP4jCyhWUxm71m9D0xpaKW2SZanSLZwUFc
cQXvKwWJE6PMM5nYSaQtttQ+TQcNa902ZbBW/fXksIdtORp+bYKfCTgoSBgodvJQ1zWF64/VJp5i
wEA6U0WdO5A1OGJALtVy8bFD7pnUx/peLWyqmTgXAsxcVIdOd9VBKqMJDWyL3H+4tsHdBZcueqLB
ZeiauRUkBWKbN7lBDa7lDB4xn7V+Dh4y7UVu2oQUgI+1JtKoJq1HFlMe/HMd4YDuovME5I6c7F1Q
eK9KcOFV94aegoQePKT8OWjYB4Hsbn00iD8tr/AAinmm0MZEA7eyO2RFa0NfvvzToz3ez8n5p6ZC
FFWDuxa70uPgy5Zgh/+INI5fKokk4Nqi1aq2YbbY4xMuZx2psz226Sv3BCsgG6aIQF+oJIBey4QB
l3zt03ASjlcyWQI+pkPhqGEe/dxf8Yadb/ZDjRElt4SnX8k7TA4XJJjpT+8FWoql5n6v8BA3wzUX
gIWDih82Hj7JfStfsYqpl8bcFXl6ok9S3AJx2aQVAnlswb0FYA9+0P7IRyh2QHuNjGw72E1g0kKI
TrJacPADKjBPMogxIyJpcaWB1IEvNlMAuRTzekqbGJvzlh5xQ3LyoPaIJqUvXY/H4+ViTPcOWBwh
IBXd5oLXGSsTyFVtlvgzGV/D641b9LGaQJfJwGmRZBE9C2RZkjTNphNWw+qmXftp0E3bYKwl5bXF
T3O5cRbAgzu0vEHC3VCEmwtu7aivNAqJ/nZPZEiDWPv6JvGZevld2kOda1F3BKAkbbJZFdNBL4FR
OuluWQknq/cLaEYScVwrhuNh2HRMsRaBbHOmq1wkzAkphKSG0taUYV6g/kknVbspJNtgGayuXqYu
MR9ZfEqsgrnB8iC6Z28ATCpNzc+hU794gdKfVewQjZ4iZZA3cew0Lz0hHcdeiIPWYEkPWkT2KJsQ
h9go2lWkYhIIDukQWDSI4VJQRnSxQTHDDZ7aK2OoEAgLqLdIYZGTpu1V1/SZba78Se3yPtSGFyk3
TejhGuASUMK4kuGfssDkueDgHc0k3Wn6iCfoke+SHuMvHRDTm15cXXF2HVrpafCT8bacVuccaQpa
q7ApYuA4gJq08zEzTn7cvGi3wVGcSevHX1ZCi2bCdrKsKSxEU1AQEruNATx1zvp7aowyb63e4Xm4
y7obff/zCdgl1i0z11nDCVOcqLXOxfUDB32h3PfnA35VaQJAa6GryAWrCfiDzTpWSCnzRyUr2N/4
0QIOOqDY5Z51pr8uKj5L9o6Vi8sJ1BzpxQ1xJnyHO76wIetQ9OfCuvOMKssPHBEU+JP+UReDdM/5
2SDp3+madEgwOrBzh6ZUSEjYksn1RBDuY5TadvUcgoDd6Na0RPOvmSMDWMGjhP2SYJBf+wN3+U8q
ZMuXW6ffBReOlAuQMaG/tLGQx8+qE6eoXnYeDK22xqrXmK6XznAWKSIq9LGJYbKKXuVHMu+UKKmM
cWtCDWUN6hqytuqt4m1l31jhdh568fmfw7oVr6PKLi3MNdby8Bwy+dkaNNdona4oOQy0yYPozPU6
nl7bvwnql7aAJwbIlTDw/2WvbbC+2QgD4gWRy3SReO7GXrPJ7GWmtRKU9hPfBSsSZO3bWI8X/o8X
3kX5J4prFTD+C05ooAVvH1H075AlMkB/BPXIF+rn4AOR3GLpIemdmEW+rsMp8tbML/bNz+Ql/UDg
mPcJMEZlQnkI9AzSBuqWcTSKKAEorByoKUsVoRzETnGGeblxCt8Je7ONK2qsvHGaW2lrKe4pBTYF
OpSH0uLZNldecgvoC+iMza7oCsAVv5MC+6F95TKMj0iUdeDXTbnZUdv0zId8vJ88JLAE3DiXxrRD
T5eiHveSR2cipwDBPFi7W3QzGXgvYjrV5fs2eJlAV8EKu6c9YuM35SgW3Fg15kaLkW0MN5kRO/ZA
UGGD7NOXd2EmfjXH2jLPQrIdTXNC95amC9IHWuE9wGFwXsQxLTZ49v5Gt+4/++n5eIRKTQECUEaI
5nOB0VYw5OMyvuDbSocUs+J8fcNGlPrpvGY9R7Xlkwt9/wSGweN+aAH24ZN/Z8upBsyH6ssBGHmg
npKFnHoo0mf5Llx3cs7h2zQIlUE0x/ihj5zKXRQrwPbsNnOHm5S+1MEnyixUTKwcvUYm5N8dIZul
ie040iFEaDXlRIchbSwDjI6KK9Y35JG8x0LjgBK+DZ/wVOIajw4ixgxV2CKRpOgdFymwnQKHG4LX
ugSJf2Fm3AlQm5VsCj95xSm10fn0SWke9MwvHSw+8xxFlFeHHEgaWkm1NMragEkaTjGUrp3wbo5s
lVOttj7csBFizSKnVigxh8IeO/KIWGVf69Oyp4lhDvoh6knavYQQL4yh3NORRaFjJox91QzVaIZ1
2rP1i/GAj1vurwXZDdLfVEE8UwTPtJH1++WIP65TfZ7Z0oqEqNVyftau8QgObnGCStRW2iYkMQTY
YUI+0kqJU+L1iRh+sCAnTc7J0sumRiuXvdh5YnvHyRVoxo/J65bFoXtfgfYG3zHJTK+NWoQ2Kw3K
IrFKMGGIVx5EUif+aJnKLlbE7uQetXANgnlZ537OGgPrpJUnxCQYfAeThKhWQLs70Q3V3uIjcXlq
VjK4KxQkJUSYOzNvw6hVnO8IhqgE4gfH2fkAZ+x6mAUXS4zwCtyocmiDko9uauEF7OgnjCPCCGEn
DbMNNKIsBv25eJwNqFnHaLXQ0a/nm+vPhOCJIR7u+NOCrB2WELTceXziwGomM+2zUTCLWnc/+pHf
wIP0tC0RahNkhHQKmojTmS9pM9v+m8EoWimSkVSGV5SEzJFc0RGF5sd/HCijwdeGzAnWbxLHCMmN
9nudrUEZ6vMcw06AtlAkp8QSaxqo9epOcDEqlnyb7G0M9n5RGNdZmEvwde2rsZmvJ+5noOeP/xfz
m4wsGMW3yOsIzCdWnI0NJSEwu6ssbOaeICqGLU2zJlRO6jseDVpSbzZRtRQZC0TUk79M2KSTj7uE
JpMnZQA6ELFVE87zSHkUo2LEoVhW3BcsRmUvjogYH5WjSyhOV3C2CCSlKK73zIE2IisgL6Z5jniu
gqSyhNqwNSZMLvjkgmx4p8cCTS9kTRhQhKWsCEVwc327NNIEsOHmnN+PrWmIJ780zM6aa1dnT2db
KLeDG/H2QLHJNCNQDEHY3LClLt2IX+YZ3N9Yq7EuIxTt6zMNAbzp3BWB/NJxxtvV1qy8T1l1ONML
4eCnx0K+Zf6gvEe5iodzp2L9UOYpRAdGIukxpkG4vOFNUUcsukeyRLe3NJgf58QrZHT/vli5HMZR
n/AZ1aJbDkpGwfJtioMTStwVmHOVUXF+bvUVaj0SgvRF7CLRr5adBXzn3OLJlCkW+8dj+mVH5UcM
6Ho7QCXVqjmnISrFZ4VXvVGzT4YZAQoTSFZlML3kNbcFv/SEuU5BT24sSXAJ+8eXd/UfdUo8hTR9
j9iSGp9/kH4RP38PX7kg+L0iNGaQXDtxcoRqUoNUMqzMAQq9sALc/wj0xWEWU4+RLTyLWLr2Dq9N
XKuV4fk8jNIG6lN4jrleIvrW54nlSIbHBsjAkqCROUwwrXIdAib1s3Bo9ZvGMU4RMzNZE8q1S1im
IFc6H9BjSEbixHXdg5kv2IsddJEEwmRJEDtW7Udb1i+bZ/Vwwb5HTB7N7wQwwrYab+693QVk81vA
RYu1UYqHaubHKd6d6xMWiDd0/DkROeLoka9F8w191q1//8VOoQbjQg/hTKgIwPs4zU5/l/OjdeoE
CwQtxy0GvjZoy3KPQRfh5Zfte9BjFmdLTpAl4CE5u7iZ7XMiZUZDe3gAUIaKXiAiWtthhSxY6WEh
DDYMuhESVd7rMj4rb8sG2WuVAQqmLTP8N4s46boPK8ks/BP7e5y3QGh57IPpNxA66VAO9Qjoh+BA
BfD6LHMpF7BZ8yCdiwJ2YdFNNScRWnkGbkunvuyrWno7f2m0976kJKJsTXACqRcCFTj9QEVAGcuz
fA960YeyeOOWtTP7CpeLb9Glp538zhUJMbcWUva3E5Y0Kb4c/YbtK2PWaRjt9RDFIwXcRI4t00gD
11IhPvQYSKIPdq4ykqqKtdADFM/y9R7A2STtVK05NeCX7Iwh0nCeYDyhAD1U/dBmXUypC800BaQ7
olU95iVPd1AJRJkCULn/5M2+XMSRRNWUe83ucKBWAkiIe94ojacww4fazNQPDA4Rk0nB9Kq64jKq
TTnWbQOhjYRaxE2BNequ9yQqOUoOIOUr+GfZ0TvuKJanJYUJIpdorQLohXhAbBJWuRAOABkahm1c
Vv4ehD23HNyfRI7OzEWReE/4PJwADfwxvg+x93sirRODOreFq389QlY9Olya25yTDpPOJr05/3h0
/jFVcsx9F88EDIjiFyev77i9MBidsaZA/7p6apxsDq/Z1FocTBeRmpwYaecButKI9+fE1S7nQtHl
pcrVR57I5424eVbRjYrr1ZKfID5+KL88ayRbqVpHGofHlk/w5jQl3Y8ksd1mF9G7wZUajKHk0DLV
rcwBsOzDZfUri1XgzdTMccY9OYoC383NUTIS8RXLwbi2YuOP4ZxCWGfXEMf2Imc2y6fjEF3cFAuz
RmKQH8RbCudDkRvy7EltpiVrjE7Zt7Qbq/HFdouy/dEGlg8H08HdM5BH5OQ2tidbv9W8tc3kqrxE
TVX1LUedbYBIpv1TXxnNaRr917HgOnaAh/LYPBgBQgM73/fam/pq+ZrXkJ7u9jhq7Ok+Vh7ajLhc
IgsX2EHe83h8tS/yHt5hCGsV2XksFcpcgL5b0VLbzBvU2U1jrqF9uCXXZEPMpaaYGjqArkroVxgP
UbfZbKpcHqjIni7rKWOymEGgPwCL8s7Cr91UNL1XafbYUaxesZyGEnsv7lLMhPdC5Lsh4SRhPZeK
+QdPkvIZroH+U6ajMgY5t2/18P/Ei5CX9hbbP/DRxsKqXG2xjPbntVIMbT1lnQBcf6AObYxXbv90
MB6bj1o6ZnoMj4yudZqITHIRX6UECTqxrAdGatEknpff/fyFF5IwYdH01VDUEadf1zEdPuP5jwIP
K5BBBU3zNhlaHY8rwWkR0YLY0PIKcTpXN7qlqz9ifrK5UwEmopA4S4RmWd49lwd+eQfdsUSjcIvX
g/1K5CYXCKU3I2OQw6osmLzj/9fD9FEAuYUR6FfJFJ++ZIGMh8HsJU4CAEeOt/7umt7wl+jS6dgj
5/+8nSNpEjQWf+84owFaE0FQPmMWXTCSfQ/4/9lhqBGnKBpul7fUx7D9jQbww99jueWRnV5cXc0A
TVdb8C3YauJ+dY4k+xi4Wzvk8ZOvrPGh8Pufc3hu0yc9ECn4eMGca6RDk1j+eyvaFZyZvN38N+gH
OAs3Zf3ZyFVLr/VPsmOdnPrmbgAE6U6lPnTb460RHj73YMNkO5etXI0iOiD6eWS5p8UDDIHofnJY
trU4KBQJTU3upAI3Q8vpvuIF4/I8KrZBWKTB/4/tKLA49mNBDvjTLeX/NgPtZKc7b5Tj/lBf5+L4
N69MaEc+Q38vjmKZ20/IN4U283m6I/o+NZAfP4erImX8ANQz9yKH9EDNxTRtPRpbEM4J3+Rw0axr
MqX5t5nwU5Ad7EiwvJpcD1emH+6t300Uk12iuu5wGYMJ8CeQkrkjrkJgzcpwLRqwLDu9FeTp9Ol6
8ZWUAeYZhHQWBH70gwp943hpyC6iK9lZg1mDil7e/s+qiM7ZiLXsn3qlQh1HYdsnD6ZFSKtm8RBK
2GI39DlEmPD5sFHhet+gf3s3EXTh6kyPKMtn8nlvlK5fLUvF0HTm0tsUGwN6h4uNij39DRv5D9Cj
5QKAhHBrLfgaUhLSEFy3+BU0kqWvBekbUgzfrrczrphabnYaaInvyze32DyQ3NCyzXaDnqyvjek9
xKdz1Z6fYVq79L4E9aGM6eO9FM2JKlahzPltTXf19RXy6TpsCsnMWQxBJHSiO8F46F/7aCW8TFmA
X9xXYJGzi7NmMfEihzBR6H+QEAaHKx5zkDhyOi43a01hPN76g03rewKo828at5EgcHGYoHeVD+PG
6l9CtFaCiFhg5UKqitdTFheBQBflqDp2vDiVUhsMJBVx+PEWpAxmh3rQLiGv1PO9LcyV6gXzmb4s
/Qoba2pLSVfUY+/1UKMwFfnAaR5o+OgTyI5Izn7ckHdQo9XPFdLLStaxGtwyC3E9JgMkFlVXE3e3
gbTCm66ayHR7juG2/ec2MqO21xptMhfCAiSDqZAlRLA1q7slypZAzfp6DPJvoOw6dnhz570N0uaA
EAgGfAOJFC4PyoR9thRSLDZ4dab8055he332FKaukhC24jse+i0opfuS7PGMiY8mpRg8XFxBDdfS
sNqUMqgFo0el+/og0EeZ6LlRsLr24bwvnd6nf8LeM9+3MnOp1YL2r4XnPaISGlQuQBYUmDfp5kXs
3JhHL9RIPN4efmE5Xxj18ylXRBvyV+riQT3x1dYdRBVqQMGI8bOgKHQZylCEz8Z6CUnVsq2oZYoB
zuZVR4+bgKTcMhp6J/ho/cq8TL1A26ydXE5x5MF67gV3MSvMOCGmgu7akvHOfIGl12nATeTvzjZf
U2PTZ/9b/5curLAu3EjR/Cq53vngmS1ARBp/1Rmrbsi3oT1q4lLO4e8X1xH/yWwLupSPtsaI1se5
TscHU4atiQODJiKbGfsM7d/POBIsaJM9lkJVFOz5QBRvPp5FWHJLeIEwYFrqxo1c79hb4gGfPHNT
gnkYq3UL43Dn1WeIMsWnjlwpybZyT59Ib64mr4FeAhoBkKj1I56wsCcpRjVwxfCWZNKC0fLJvF2L
cajEpohEefx2FB0MvMhqAYshNPvm82Xg07QQZ9owS6zaS3toUuQCnfdTOCeSxGkVRwImYEoMTn38
y+N5EwPo6DUc8w+MpgLhvCZT7zJGdCJC2zHCVb/b0JTvBYY6573L3JdjZbo64oBlHYeZJ8p3302c
3cqs/gbtYomy4r0XFLq0yenkKn+nZxl22fZXqD82WXeJ5JV0S81MM23HSldn7YlLxYZbhdEDSx8o
lTKeytikqTmIYAbLeD8uQh52sq8ArPLKCGO6s7xLDrfuhwOvB+MsJ6YUutOu1cZXkA/FcIoThwE/
28LOgxAIQ4zk87AX36xwPbOGjE9XkN2ul7ezXNFHYvMJq1S25K8l34J+QZ/52tKL6j+Ez6cdcxj9
6ejCOtad9EU1xqUz1W8GuRfl6ATxweoYSkFN2kY+jQhOTUO8oyBVIVR8TU14895WMiXRNgfx0EOb
yY5+/9A99a2181W9+aabHYEcQPCa1n8kynZcrOvYZg+1gZrBmVK7LFEfsFZNtq+Bs+DDH7E77FG1
aQcvremjhfPXqCCJY2CjqTvjiSMnmoNw+HI7B2DL5FZLAgZhOgt96zSoBpd/cbyKKt/UhFw5H4Fr
eA7JY43rWeLBtNI0nBd69sbfCsbdhA6bZg26aX1K2UR2fmu5IZL9fsKvK3KmRRyzY35/WwOCffAF
nCRhKi6chx/6+mw4a6g9KCAU5P9gT96duMhWR4+KlgnhUatzfCkWNhznfp5SKbnkV09H4HOJyx/o
+X3xCuCXVSQxOYbvIb4dE3HObk4fmPMvlPedgbuH5MRXAbeOu0ptH+RKGL6ccQkLC1tR6ZELg8lc
4M6VELW2EZ1ilv/Ha0MpwjxGyY4/XwEtzmaLHyTqx1aNaw9Ufx1r6U/NrYeLBhzfdmvm6zCNoEGC
F/xphBTy3UCk9MKagFn3aVliOmEsB9pYjj/YLr6FTqY6A/npW0EJUvMRaLkQ7pUf7irB1m8EozU9
G6ZUcOJX66XoBl1hdKDIh+hdp5vG757iEkR/wVG1zXO99k8EuYm5fNyvwLHQlYPGsV32dJRZK90q
AMClA1Th37//MZ7yQMcJfUwE+14p5ZDpp5i3DpiSixHAICBcdCam4hhJt5e1/cFkbaVFfPLxZkH5
NUArULKx2SHnNq2hnnOaFIbgpblP/N5ppsuuEskEny+teSvrynzHg/iV3+B7cnYBAitis293onaI
sBUxBJRGU4HVQq8d1mh1fOtFTW7k/QQ7vBTrEEGeIKMhek1Md+4XeRLAm6QljHfOpCGrfJtp8R7F
dqJjK+eAic83UA2atfs46tmIKDkXcdGJTLtJetbTyES1ysV6QZHr6zSBEsq2cJ2zw8nwQS9vllmr
pDTyB3ooIb2ScB/2ewV5eaGTghbw7oQv28aNyRun7WCY43ENnzad0v9tONEBS89Omo4HDLDnt6Jc
b1iA6AGIUosqYC0SAnb9tXYhXq84DzZrCRNUs7+SmlwMdEfS7dAP44U4XqkVZTKASRgkbuVdR29E
5MLq0x1vLFl5rxOmO9qeKYWVh0bH7HJZnvtS7Agdw1hTCWLG2dh9mIFMDAA6ORq3hMM6XhDuo2bx
lZMRpKpRAowy2tUbJbH5P/ljv6CsSa9ycJmIR2NpgBlK3Snmk4XO8bjxgAinbyI+OfdVqwbLrddJ
rQ0FirS1uxq8Xny6WR9xDMeSQ9A+Na86bs0ZcFT/baghBHzn2vMs+VzIgrgq369dk/ZGO9P+ZP1r
OX2jTp0ya31ko2Ss1MoH4D+oFEQSqRTsn+pNn9tZ4dAK9V6jJmtyl55UaMbFPbSvT0c51yxNuiqN
DfsN+5lFzVhovy7FNCc/vjl6xX6gR/ADthJDaUbJ8X8yZn3DY3qpFxG9sUDk6seZfqilgKrCAABb
kAZP5oAcxMlo4sTEfm85XYy4rpHerZWWdpWzwZ0MR6ek9f/38U2BF1VfzsEYWOlW4F/0q3oxFMm9
8WvqnrDvLN9/mF0x++M64VGmvQ+1m2ur1sG//hxh6gnmrtKPhujB6P5UYjcLEWj8mkHirk19Yh39
6vdTLcnxHmzNyUql57lhetKIrF05t2nR0MbokWroeebIB/YyA8AKO/qTvDtLje+JGnCQsRtd1RLF
SDIibtRteK2Y/4piIUUrCMtSw0XWrN6HFbiumhHPGeGCg8tNSZXJ+MgTa4WzbC2Q5845AckzUZOf
TjI3Gw4nHflrYGQx5TR1xNLkvTVWrgsgiRASFPE76I2g/lMjvGjIvwFSDc0xjqj3u1zlULmhkcBV
RSTa4ir3Inh/FL8EK4N5K5S3eD8pjM/u6Lsg8HpUPp/Fl4X8ClQYnVCoU+x8RYC6/Hu93DdXMI6q
mUq+S31FI7EATmrELTRrLabA/Svre2TiluTN6/6sjhomtHEb7F4TUm6SCWmCBMi0LXEKasN3rDAO
MGOsqK9Mnj6uLJdkjfCeB/yF6CE44aKsfOPIXuo68uAU7XvzFjC2Iu0EOHww5NPcF2hCFIei3Kft
BdMMXbp602Y9gJ6sP96KE7AM5ARo5Jqm2Nawv2UEPwmwPmwL7XZlgwZ1Nse1gsgZYDfkf6knV3iI
rP8zrez29cUkOq1PU+IjQURYzsIb3xhKlYZ8Bxwc57LeZRePiIW5UDMkl7g2t6QfqSDSHnqgyKWC
Pu1ZHteJ79RPQXetx/uBplJ2gGxsQ4Pnt4o5uvBIzyfcRn3zLYtPy/xKs23qXADMfpgjuNOkyQAg
owGECKzxNLt9G0fOXREdQ4snYigQgY3QGB2rYsiUtyv41e9b0AUN3IKRTr0i2yMKSvv5P1THCmFG
dVATnUppUKy+DeVtunmow2UJ+iKxFcA30735Kt4+XiKAfqbVJbV2DPDeFoIfQ7n0e9bpB01abTXg
yeXigxlMCBKI1L2Nu97x5pTqxMP7XjJjzEjlevKJYboWu9ToLXC9+VYtEu/8MsuQzix5SL6MOQBM
88banfqWeOChF7gjV8oeQCwOIvlMTprm6fW3oSUhN6QQlrruDkf3iolHdCFdcD+DlmKg7uQHtcsu
rGKiwbGpDmX/9GiR6usChNRJFyWkNjhEuhVykDhlVV6BN3motqxfgtOdWS7TjPiSMqvS49zbnQo0
ZzkoMWj7c8PlyT994xML07mIQZuqqfjRtZJLdkRRUiiyTas+deoiuUVwhLHRRkt5OWToOfilmGZg
YSdY4vJ/SM9vw32Q02NBfABYN5XLzGr0yTQ9w4CgpnR3cjUNdOikToQXRi5iDFP3O97eTKJHz1Xe
YLsdKxwYXy9O2H4l7aIdyAFoiVGIbRrV0VwpqK8Z1YWHeuM3vkPsKRLA168y+dabF+dRxLCTCE1j
z0FPvkjWHDvqUliEfzgeWO8IiiJNHoJmLKeeu3YB31Di0XX38+/KoW1ntHhhNQuCI85Ya8XFbTSA
Xejh3yxEsBElFLsUB7R/WG59zH6nhCAmgW9t44w/ilzk/daVF08sWIR8dULjNFeM1EZ3U6UwKgLg
cl+bS06kFwdt/1bHTxu0WTZUG/32nUWEfhvc5d6tYsS368rc9F4cusnsfvyk+KCtBSCsW0aUEMMk
56Ne0tKFiGwJsqdcb7U8DwkNqd07VWj7qpbVXs46bJCBC9SIN6Tu8QvqHjw1LETjEiyNuhJ8GBOl
3FlPJbU5JRD94y/9eh5sgxpf2SzsHyWfCiMkpvxUeGZbC4eXLmI7Lo9FnX/xHhhzEf+emBKxn9pN
yT7aVLvcETBRtuHuUL2V2a4kw8MNT4kSZCuUa3cB2/W/OWl/0YjVN2e5MIeYPOPUDLsexw5NTWFF
FRbL/UWPbIsy++l2EbJ8pO1jU6SNfu04TU9ekYXejSVEUcq1VOFhIxbJ8pcjzAKP4t3/HCeOuVv+
Fm5L1am7S0CDNLn20fwkv7sOqTvyelR6FyYXob/qm94TCTYfh1V5ulwfwufTpe0MZBOdRsK4P8ip
J0cKICV76o4WnD7eF9qNGnfR/1t709XZ8DXRs9z0+BXPMSoGO2O7S8v+1K/dy9RFCjO8u377NzlD
QwzLM/iZFVadCLf4Elan5aZJoXkLFic8cNSHKe6EQPqdP+N5/C3RO8SVMX49oGtd9hPLLWOLgY2S
5X2rZnlu0hXsConFL7P294eeahoWuFtS6qOQCtM8cFZBoPGZAwn49DVDyHSwLJzkXhW8q8wWrVVW
nEQ7cfM2oOvvVJH/0Fh+NwWG4dgZjW5LBF1m7dOeKMDSADSqQQveCrVNHtDVJ5uknnxEHhIaf8O7
qJBs0opvlr5emdfrrISw5yKQtM2qWaybj+Otpu4RQrq+za5VcefuXeVxUYvO8WG72W4YxTsfcgdK
5DB12UtwksPzTJ8CaUmUgJHMZYaD0aC4gAYyh6mgqZDY3VmcJqPMNcAYJ+RrYtmJRSeFJQbQXO7Q
SsO5INUsakUIqNqdmVc3HE3z4wdY+pfv6PnycgF5DcRg6V5xuwSz9TNlUABqhq3ud9N3vU0mQ5YG
0khIoVIygke9B/7dQyC2tf7r4lVbGWI7zj9tUBjipYrX3Kcl4O0w7OdfRG18VqATzRQxjQCxBidY
1Y943P5tb311rmihO2tgrrBw0+TnIh/8KQVx5VVO6GwQ4jPUXr4Z6BprBlO+cnrng4XSkFOEWRuV
Sbnf0r8Y8WyO/66cICtHCaMxiqBYXdqaovqY38LySrue77UigoMCOaGRFHezKVZIOinL1xeA3qk7
u7PVbK/IySIkw1nF36PDMDbV1j4HBxxWbUkHEGtT1F1ys5yJyUoQQXSVCJhlOmfT3FXdP6cwWFDf
v8MR2NE/WzEDpLNFKOqfdn0UQuHO0wCVsb6qyOqAR/shtt4BW/U02bISubfdzOx5VRwkncS3bv2l
WzLUTR+QXUe072oFu/Ms0S8cmV7kneefCKo/R6EAC9/pp33RNe7r5o4mBGHpcGOR1D5DNHv2pEfu
QRS8Z94smLT8gAdzsUc6NYmwPNab8vqUXBxAc6nuhFsGEyb0fBsjBFh+7EDsk9L6W4TaXdTUBBFh
xukqlntU9U9jJh8RQIeVJ/wwoPBTGDgv5+QRNmMzkPNXVwmm8znzlleukKVkLopGhsRKHfGnC8ex
SMc2YSd8SVfA3lE7iewOgAedYIBPPUztDy7CBiVJPsjOPnLU7HiaECjAVvdflGCtbneCo262YdOJ
5JG9QY1W2jsuYJmzMqSLLDMv27mm8DzGxW2m/cYfaXAiArkSTHfW0Lk0YoWJ6NTBpyvLB+s0lx0y
IGGZVBUrFpHRQWPt5glh/8+XmxDQt61feOCw8yNWadEcbTFM2gsxY/LVs+pjsijJKY9cF4pouF3/
JVt4QCmzhkNOV4I+f73efBnJGEHf0Ry279ie6V+AVdclxHeMrbzZxMLzF8vcjpc1yStr4C228t7p
6lLw56eDbBvvL0WSlrCHRlSW5jXuyce1shr5hhdIkJGTEtwDkhnQ4zlmj0xLkH/NO+8VNUalTaOw
pIDARpGLdo3D48WNS9SciWcDP27vZHwlYbESVaM/V5erMxMrrYBVaKgvclvUH+9Lqz7Xj4fv4fYe
7qnTxzJaOWo/QyLf1Gcc1yO3qvCG9JqeJ9VopxArZEJyMcG7rxiDfL4HfPrAcrW3+6hO1QUgztx4
TWnbXUTG66cKR2Lr2j9PXf5HTHxakYymYXsQwGFkYNfn8tDk96IIZEHfLH9JGk/eitgZyYgASPLl
rSlVkNn/B8Fgh4VAr4i+ORwf5Hm/hjcfy9Y4mS6YVPZe5oOY32Ik7LA8tGEeML7JzD/AnulbhNA+
KJUYfooM/ZdXOHFh3q/JT7p+9VZv2QYtn34CAjAzD0tyyHrcj/EFv8WIcJM+UkVq+fTVEGLNEGoc
WaFQMn+DfoW0vjCiQP1gJo0AZxk6Fab4WXvJ0kzlJxi9F7zJ7krGEKmJYoTkm0FRmyVNgg0tM1hG
9VfSe3ZhEZEGf4wUl2n9qbKly5tB5FMnNLM9zSw8izjcZzHWIG9F1rW1PvFNryT7qJdVKKuujw48
wdGR2LWZmka6fbBaetV4RE2ZUxA2vdxgL8BshNlVa+SgQfTal+VEDeJ6n39iam71xSk37MByEH/6
wWpuHDlWnV+pgYU9fPoAQ6PuNYgj8PuVIJ7RiqzMhFN7dEInz0i2v3Q2h1MagWikGj8N+hhPwZs+
nYE3sEwYqBiXPfqN4EV/E5VYweJlFr04IQw7bmaZb4yGU6wBGDDgs61W0Bpbr+QE9ehmTSmaZNmo
SXmcVBZBZmkWxKgywo7JmVdZgJkJCQoIVjV8HmvlDFNMM1HOKrjlMjsBN2CyUHZ9UlvbSkWbxGlk
+71+zQLzTTUeeu8EleSiD0SbWxRzU4zQXax8sUtWVRtlD5t4i1q59JMXqhMwGH7GpY/l7du3d0gR
yr/MtLnA26VUwpdiQDiY7UedNaILq3uZ+4VYIYGud8Z4PV83M641xfFiYYAHNEgKOz/Cl0d+5U1c
odSEmYB6ybXh3xChF9askvoUxVAuTvp4eQuVTZYtKzFuJkp9gnJfURJsaF4VDT4Yd4x82M+26Sce
8bbcRmF44kuKkvlABXBzrMxbn1pHlm4120i8812JcFQrDByb5Z9lVKBF6Hzd2C/Ke+iM7yjCi4yP
+C3RIYYDICbPlqS+WYZvkGoZhj5buhBUvoGkSaLZAY0Uc02ZFm4YwfV3hxJae9kfxtUO/JzZW31N
fnGsAX5gOxchMI6w4VByGlXHtcIf22/NVqbmn7/z34eyoRgIfaFXLYFfxrO1rzPAJS8DfQqbOZ86
6GXQwKDLsXh+YWHp7qfEUFD/0MpV0hohGQFNhM+/oDO7PitHvVUc152GpYC4l8CZZBIR8RLaWhEi
LyhnJfUYnAtAetIEK5CtKO+UWfSEDUX69jraJya7BDjQT2xnPec5npBuZ17ny28vc+H14azvj1H9
4WoZwbLjbYuaZiRD8EXg1qcXp7VwgGAEZ3YSsXzOyEYMwmlVZoIAB881Cf78g+du9eFbmDb0+POz
mgkU08xyvlJzTFA8Vm89IV7Ep16c2qYEegGjfHcslugKSb8AtCPs3FaY1UDeLcekRdWZhg8a5fJi
5GhAkY4L2ZxY41cJAeMZ073t6s3yTs6gy+vg3oFgnNu3jn80+uKTNCy3muHfeSO6/4CqJVJvw/d6
8pfUkgUIWjqBAbeTOlVzOcICZnu4/I6e5Q0lN+QEKhc8gWbaEsjkD3gfGPVmR1KmGPyyXIqHKGYp
j1aoglT96JKapX8k6d5LEEXaDFYSTr5rXzYGsv4RGex4/erwgS51VFrBFLJukeVKvzHkWVL0L3Qt
mTw5qkjafy/2DZuUhCdbS9GFa5RA1HFmfDIaJhL2LkoeO7I899TCHSVrsinoZ3L0MsLDGFMu0t9i
VlnylPeH+aYVTMQHOGVGAr9zlz3B9LqRq1sKQOfNzFS29yGMGOgVL3f4v3HDV/UpTefvk8ZEWweB
BU6VQkNZg2BgpO3zlWKrdZQ8fOCRZItfeakMhZaw8Ygpdjt1RI8Se7k2ma3ssu1iFyAEjZtuOdbs
dq/qJuPoh+K6vjtC8vPGHxh1SD5iLkV48w7tCpc5sRkrb7+/ypv2N4TDhNIcwKsc9OwzNKRr/UYG
rt5E91JwqzoLL+QGALzq3rWkp8EwLBOW0I2joLY2vyGAdId+VbcMELWaVdI44DytFt0A3Nfs7Ivd
zZ9nCnqS1v6C1DsyYANuzxHZsHL/VuCeR+NEPuY3K3QHEqkm38bU+5VVNlFT+vJcWNi+M+DGkj08
mhl1X88fnIRiRJt1mW8paKIqTy9WAv1BnjtwvwopzMfir4Jd3jASG7ha95HqyyVgf2DwKUF52deS
e9NVPFeyoxz8IkCo8oyFpZepGwEIf21OVpqlws1+Mi1XLT7Ls24jqsMnWLWq/GQU/SUwkjRvhRFN
4/mqw4M3yqHyiTbZStMGoPbqubIqLitViQKT5fnzORh61aBhXeaR55k5lIy8qIwdsHWqUkJlECNI
AVUESBMAVNlRmROfbvuXu3XaB8XX0isUALbQKfhVxPZHNW9ukvRM4tF8AdNyakoRibIdetoEeo2b
eWi/OZiUuyKPEhbVZTQGArjjD8Cg1Z0au4Q7eBLE9vC0mT1i1PYZLuzqbokSsaQEmxV6jm+2Dgjr
2xLmHzRqKTLhHuz+RIbfIGnSHBhfpJkrNLpiWvOGvSOjeYP5MkUN045mUuwjsFkFgztx7//X3aK1
Z442ovgDPy63bMuLCCrLnAOLYdThfyLx2KvUgBGHLp6Wtv8UHavMnIWsOF2OdnbLTe6njj7f5lrG
I+BZs/gb5LnRsGzhAUwHiRrSX6bt80S7jOFqJKCB3Vsx9HFtki6CpaNS6MUEBtPZhNxBP+DpuGUe
5ivICqICa9gA7YOcTs2McvOq2yQxSs67XRyodqQKEllZ6rj/frLxLGcmWjSWl5wZAJqm/b/32Qkl
f7vE5dKV8e3C37tjaLzHln+CIIthHy+oK7KSlmhYT62+9VWwfLDU1lDtn1Tv3UYwt22WG2/EfXqa
xHSMAfjEefkAiG4i+yADrUZKTQEcKPbUo9LZ0y4VQGil7OoCz5/DoHQPelHvtGtW9a78ujPhkhCL
XlGBCJpjAMAdtuYXCe5/Psdkt0YZotSgfzTY7hUyGcYiFF1bkY0MvTfRW8W+HpRDfcouX0dkwwAb
8aCBuzT6xoHOB/9K2tskEumuDCQrg1SoTamz8l18R8kxpdG/kwzziB+lYo+y0nudXJdkcSGIirQo
rCWvC1qOsqHSgJeHL/+LVJ/OMgGUzmouhJyr5tCxSv+Fb38jcARbeoswCQxYK5Rxz2eoVXOqLVvj
gFmkamxbJL08emenIVlVTDp5yVa3X0Dco+ZSdV+WTPUqnGPtMQ9jHkV5sxh1Px17rCO1lUIGt264
DxIgLooRlkQztfrBj3fdh+z4CgqA4NZ7SUnjA39q7mLNEUnBCMmMs6Ba29PHZFoIp/p9Xvlui7wF
mruBs/yoMdGUiQ43KjgBygLC65cXmemJAgwq8U4RclP0xZhuZLMK9fJAsOcxWpQaFhrdLS4I7oTp
fVP8pdPrEzo+E+02N8YAR4Xg0ryRPN0VgVenmDyRtEZpL5ZjwKwaNIoG1OQTkPRffTlLMFYs6VEm
H5GqByrm/FZu2JRrUio2IraIvQXuuO+IQmQt6c5I+ZuiIxQN41TKXznj46MZTJyl1AYrNEBhhkk9
g+U1bs1td79RHLg9xcmYKDg/7lsE44JlPArOQE0U+CJU3eDDixcdVlOGXnBbzCnW5+PvFvqGtWo6
aYUJk8A0vhHfpgEvAgP68bxZ2y2kq+mmmiviqGF+QLiWUDvj071ihg0MlgpNxZLorBPLufyz5GLe
qHW4qaW4SbWAgYU7zuboU9euuTMWzlwdpH03AdKRuqeHf93vR4Clk9PG3gKocwjosqvwhIxZWWfw
Tei+7y2Fs3zla8ZncPPN1glO7KIpnhIFlJl3Sg+1isb7XdgG2Uc/23nmiD/ifijLEvRcmtY2RmsU
7lHaxhQlWuTeygiHdqx0faqaRFeW4BQj/TCHALKZ1hpdYgfGO1bvHcNzhzs7amlb1Ky6027q/1Tp
G4jGtLkt/7ib5XJVtaM8KORf8iHnAFMGYAABESR8PnRd9tmFrbCKXgyl/JWLlz5FWP034n8/WlZt
8CYfY4JNPA4bXwBImU0pfL7zSQ3famaVUJPDvNsoD7rBnyGBnqxhVjwamlfvHigXMsRWj8vB6Dds
zphkkU1dyl9DJsKAyauEQCmmKjpGDlRbM2P6JtjACQNGYJYjhXTb2a70Al8N+kA3hbwJDn+c02cP
8a26nIHNG18cEYLhWbw3fQt2dflvZxQk8mILWP8583bCQ07TkyhGMx87MUAKYJMGwe4P/linw8NI
vKGB6IFPqRgGUWFe+BkofAwjflK9KpjA4AtLWYxJm/fWFnuh6eEbc8//DGaG3n8J+1Fz1ghYOM8C
WsIzU9g+nW/E3vfytkZx7G5pZReiiTfjdDfw1y9LCWwKUxtgvBC2BlnF5azAyONN9NdF3lWgGQoF
UxLLfJKkkCfyk7ux4oVtkYtSuVcBS9kNuMztqiCwMm2onqYa5B19ZKd3Oqdc71azW+WyTV/UICo2
bqG/jyt/3n2XdXz6/dKDq8Ahq/l9UFhl6lW6LcQOwjxNNY7yM9R5892BNlX1FjjRCbDQNe3P/ixl
uLD2UlDgSDQNkcQObBh8DBnrMNvLkGArIfxvyx6qrRdCjwgkztStNyXd5sV2cONbtLj0lMJUm9mD
aWJEHN+J0ZE4yGfaAba04KTZeSz7Qo9+4klSVxLsjHvDviQJwZcPHxFmltcmH+uVOImWuk17s6l/
6uMi5dTvms8c7OgZ/m2yaJDKL7//WbcF/DnPNVgS1/R+mO9ljYHzpCUr1sTYEQd1FjczPCdFr7Te
r7CvizNBRxh1LLSfgjuMtmgnwMlnTzcEj4fpMhJyMsvkHMHSQVV2Flrt7VIxKHdXw7Lv/RcGttIf
MwbKEiirOKjCBNpckOJiPIsR8go7iTql2mc/w3KmBygzDd9aq18y0ivQVKrb7pFLc7mzhz+NL8As
iVTvT8xaurxK4fpeTlFIvI3mDubS/TTd084h+fU4twPoIeRfxCJt4nMj+Wjh2i+h4rFi3hroOS7b
+TVM5rlxWx+YlDr5GQS4tFf8BQJrSy16lizuu6jkF4nu9w7qIk9gwo1N04/Ixg6cfHTLobz/7pI8
Ulv1ykikOSPCYXyNTyYscLrvkZzHIhL6UXzFV258AkGvdTGIhibA0kb7iEthlc36yvvqSRX0L0ak
L51mUF8n3KO+71eHt1c/3PkNKykIz3UTW6ri6ATFS5s6hvQ9OG4yYnlE3v23YTdw/pD2k+A98bXs
8pvO2YwzUntEHrPmqeph3w8R34lL8nhvOxcfTTXuSHWnu2v60WFMKNxGQwnxNn2EIRNAtZCydFX4
CEwL7YkA2ojq3D5PPT6Xuo0w1jQT3V5P8LWyvKecTI2ibMw08/FUwI1XLaTtOdbitZd8mX+ntin7
zSIyvkAjStY7lSynCEuUTuKgAm65VApiNto+40JaBD4I7f4plJ3rLpePwx9gwDKBNGtL65g3mRqP
LdgRFftQXmYOZaOXrnAVe+8gOP2/JfwgDXyZ0mSrEnwNpCs4sNylSrcrFc2iqDucXkq1pXBbIrxV
kNSSJbrsSMqB0Xxqx6S9AYEBBXy6M3oa5yHbFqYQoPHJ2ey/vVNhyyD3mui1JpiMYw7v7wBV+5MP
nJ4o1TIWaKsoXitXh2m59ewj8YuHZ9MZre5NjwHhrtVOme1hSpvgpSj02OePiEzjMgdH5oBysU+3
tAfprD1hOj0SwQowbdDHlKypsHBskmgjntO/k7Pc/6L8efPLtfr3fwJC805Oi2ZynsQan7+Bs2Ua
5BwLT+bsyFRYBuYoWnSJwKIaYWDI7J7Kt2sIRETvk/ukSAMgRAV6QanBtq40UaI1SknoF+0GnUrW
6j7BrpZn3YwiyhAPlVPTqYv4Z5RIcUvLTkHuZS0A+S/kIGsmcGq9Ti/GcS3GX8+Hir8CExf8rKhq
7lbYiOPZWCosOvKHU0j+zCamjaxyhfHjUrqhhsudNdaie1TRe60RDedQ8E1atA1OVZxqBbn8Rlz1
IB9Yy4EW0Dt02QlLXADCVEwdVvmHkYe9KWJrwym0B/YU1ORHaKeTQH7LYdjNnHmsDmekzh3PwgTf
OzcmsJETQxiN0oFoHSN7ErhhI/W7MhhJsD9X9h9c33eillN1PuFMoMSdbbLUUvdxmH+Wnm2yepF2
JbsQ7ZNwSBnAH1Y3OoUvO7bjG6e4DNhBmyNsTgRj2iK1FzVnBxZxWywk1vbrUEVkDOwTXWgkYrbz
0HkvUApcD+taf+E8BbJb2grMeaLLLCcWz0z8OlOU8pdJ9eOLxDxKmRu/3Afn6LbZY/9GLoHteGn0
EGIw+AL+IdTr6rSgb/PuLo3XVqDJx8E9liC4wRlgp2p9XMYmEcuwqVxELmHcSavNVhlTEBNFVWuo
kXK5MbgWnhbGWBr1Vq/nvmy5SfY+K+IGcAb3uT4EV5ACw9kGbhnWH7iKbphAi0Lo+UeCpxCLD924
53LQukjtBluOxnu4bGOeQ+KycyEDBzxKTmSIJqRxZCYdYaxXmX82/QDQwguv4ccaRTTI2WJugcrg
RjwMVW9KLEObOX9YNMgInMujUftAY/79rwli/GWmgbhEeZJAuDqDm1OuY1bmycKfZ8TkGTJJUhd1
p5wDNtBMQidcRc6GElGh/L0aCT30WpdtFxEpHlCBs+t2v5aPGLfut7bi2M162fXOs3o8nrKduqHF
QaEtcCg1Bl4BzJkkVoOKwbFNRIZjWqTFQWyGUAhqHgxPuNlZtiGT8Qo/sjNQWWy3mbDeonkrcjEj
v7fElIQgA9mreh/AFCPwQ3RgSkvBpiJZAim8o2Vaqf0OvVQuKqb8GX6UiSX1V+8bn4cJCDI56+BL
IQYfBVe3JbkJE34M/42diNM2asaAz3eb0kfEBIQSs3i7sKoqyuOFxJoUkocleRJreSHrv73EJucJ
5pZzrjwttrq1D/Dg+llO8XxDhOP/jj2iyd2eaV7Oj1Fbq0QgcA7Eyoe6KlzjOVZV2ttFtKFtBgPl
NXmW4jI2Vfz33ZXKOYRldGb10Kar1UjbErt5Erf3fmzAwxgahdI1wFBB3r7LC3h1Q/9ADGN1BNPp
c2v20hvsizNDcsAJ4/wcataRjK7L+EezElWhkfbqmlnkp5Ma+JcJFDOIDEN8qytJEOaAEsHiC1A9
VduZTNtzPZNbX5Djm+/GhA1mI7/VF2TItQSiGUrGBW0bOJTBZEHGSMFlBBIBMR6vOHSel+cTqt3A
dd7l0fICdI8h21MJeMG4flF0FFzQHnDsdF7xMlP0QJeHqHjSxDc6TDtIQryIMlR1kGwSObAZz0bM
64WzZUDQg9g3iEQ6ZUCm0jJ8iI1igO5AEMPv/LSQh1B5SdXe9pMkzGGmV8sPEiVlRJ0k85it1sCd
F3RqCdSQQibN6YL/PSNy8v2Q4WlSpLI8RHTBx7X+ohXXNLDpXfd76Ohwoba+5k3cZRCQMD0Dm8U9
yaaXqnagRMF6jIDLR/VUcH24jlAWNXS3cNpDzfUHVJ9NDly8AxEloQN0DCP63keLKemhEaa05gA3
1YMvRdG94maagszMLMdl0qqK0wAA1lIwH5peR1HLLfsst2FPHSZIwtFfkRDkf/qrg42vYQTMASsb
AQOHQEgBcJ5WHZinti7ulp0M7nVgHOGkzaPf0EdZcdW3l1szsXh0aS58XBc/56tyZwrL3j1Ze+hL
Bpf0q+pSiCW407vUlLERvRXFlhVQOMAVucDTezxkhrWDRZcF8QomHr91JjvAQTzCKVaH3tO67aLr
m8gFBVEPJqqnnGOlZUUmEzlDQA8dlbk7o5f8E0IRAjH36LQaKll2HWQorRCRNpGHM58XanrRnV7X
YfygW2ULRS/bBrpw+eALO6EWjRO9fHkDP0B9XF2KCv82bPj54h/LeliuTRYSLxF4QOTIVyFOmKVi
miIKIFss40tO9ed/+wIP8VmYGkkNEcrQOLI2w9zzb8YYPIHMQ3keG0gzfxc8X4IOhTg8WduaRAyP
q80KQkzcPXWLGFnbTUMzPJm5dyIjoF+hh2HQHtcJw27UXYDCeQBFNx90t7l2YiWK7gLbbmQaAOlj
UWtufbcuFpLsSyhbeOyM1bRKxetaUjFdy3/lhtvn5ju5AwkZC0wg5+Qo8l73Q7eUrEJh57WYdGiI
3afVadHKl5d1oqfIx9vQROmpfJD8TpDVXc4DLpe6oDZjBN4x3vCkONecDWKRCQvvx5yLm56+jKlr
UlzF8jlee6x85Ld60x7l1gdg1LUzLjBBZJCAc3+6dg78GfRDktBNYs4Y8JKvWqeQgA5tvr6wsSLo
M/kcRzi6ic5EtDe4tE5vxt7jieWVwWtPxJF95rKRMEwU9b5vj3WTM0dqWjxPdzWQtMkvo0zBvWIZ
iPdncIe/9nir8si/9tc05orQzm+RUAb0lKqSParv8RBZSAa1n8R50/ulQp0VR3qDCj3iypp2Pap4
Sr/7Ub8s/aLGvHBOue1AYGnU7lUNrDq/9KMaLAZYDvwB3jN1HMPeuelzbtShq0XJSBU307bBcju9
5S+Eld45mj88o2RQJ8OXSHYLcdrVK3KVSa8eBu8E5wGLKlntIqIxTOf8rOkB5e/o+qR5O6vaVYom
Usd8SPXvFSGQDqmWgL2qzjIWIjsA7eo9dPuBbO9PyVHI09mB5DM7mXyqOCkVuv/+cgk1O9VKfFPz
RF5J0DHd8SwI0qBWuoZhXtirKoOLyypvbRGAFFL7t8pCtYsSyE+bn65nGixqwXQzQ+1zY3JW+bKa
yiicSgDF8xVAFT6SK3+PNyCY/7ik/2vg6T7uROjKhFX6ZMABr/lMBkb+8B1ag2wqFbSYHa14B4FU
f3O1f6VnHYuAqwlBF16UiTTMu8QCS1NtBBHrkXP3SYw64IvpPUFjwubXwOMK2ioAzZw0QtErN1oX
tmbNwACPVfphEFiDxRxG8WA3PpI1nAXMBmfYGMa8iFI2wGmBO3Y2ywIKAUW/fjmsRf7ajaITcHgH
HuhBtQMtpYSFudL9+BIuYd/o+nR5R7nsDEcwrjl+D8s5GTCdxsbYXeqlG45QZnQk4Xsz0ukKMm4B
vLvrAg9XbyfE9lQjzQSULd+0r0V1MJyNOzX3uwZZGm2OyPIKwxufUaL9EF2tbIZWUnQCbceX7oQ2
oG876lW43bCQnCYUGfgpQgChs1jxGJxHXC4N2YUt2A0bxrWBsau/H844eB6pXhRLIvXZ5kffFZl8
OfByfDzhw+zHYQ1Ws7jLCR6hj1Jp8aMGEJcLDWCvZWxoPCj1KefiHGlktj/A4oA/OFCc5pnXNYVx
Cj7h3EOHgdL6MlTL3/9kquefp2P4s576b/xyNuWGV9fqdo0XTq6z8tYYyxq/vm0inapIVIWWQ25f
pTnt8RiGLWwfAbCoU9ddoGhKw47KVYKdL75Jv0KbU7J1n0k4e66E+5G1CZd40TyrSxyucjjYCTIW
VeDeJga9iaCRpquILTJpMXLuOUjhaW0AWZrtfPG6+V+hI7RhBF1obPP/aG7tWJz9VjyXg+z2mdpI
PEav7BcthcNsqBFXabKGr248VUHhLHfR/RmI/8b/hRlOmeHN0xnT/W2sz4arSiSIxAXWpr3bTPPG
skcEsppHYQLSJtsZITgDmPn54Ahq6nrUPiuyCWxrFj9Fak/L+kFBF5Rex9ylO9Jaeb+7Z82433yx
isJXAJQFuv7Y8NKioKt8EsyLj8NYOwuuelQnfJGUeHietvyloRd7s2rHdeU8npgiw6pCcnZKzJSx
KNKIXiZSIA9c9JEMwqEN1SNNmWbbMsz7FwKAPsXLOF0Bm95bk3OhDO10TFH+vg6yScC2aVkxsrTS
WCZOV1plq5sV7SQoIpj9mXYY1NyKjBS60g3kwShumye1zdY5HKi5zJ4CbjynaoSPDA9oVZBd3TsI
H4rLCqquh6lHpU6Ka76m8j0tR+C1S6eemHbshcMSWNOUsdxvmjJ9TDMmmQqqpJTKK6Es1MW8XDmY
ejnSlouJKcFwbGtU4hrlQ6e2iHSyTda711Cm23HOv2mmKQ+ekjjEMTMl8ADZYyQf9vu3/54X88eq
XYBaj3rNuDHalcyH1rdcOZacoL4CfgPhGHC+viWQmrUvu5mKoUi5K/LI9WMIdSkv1SzAmEIvy8An
6ukaA8JnMAxr77DyjgKaIL1Ia+fEI7pDy19YaScwFXwBUJ8a5RXeT0m6CznCY4XwSgCcAB5u+zih
HOeonfZcwjy+q0K77sIwcxC6Pz7DvcVW6T6Lb05LuosDKddgshqkJR40ptLQC7tgqJ54n4HEA6tZ
WibDAxINSAd6k1rG3b+d71cXJ4XoaYMZuOdoSWfsXjGrPgIU6x/NepfNFW4N9BhjSbyVGPGP54CS
LSXj4QQBpr9QwlbzbcA7/Xjj8djekAFhcvCSxIC6TkZDYz933xS+PztWjtA2w5OTLMrzHnIn7ray
TecpAvTU0uxT4QzQqBKDwd0+Qc+2JE8mvAfubUwMAQr1AMtmbhLMn/Zzhb5i8fiXTRS40LUMlrQH
05/4ZG4GEy4GhiEkFiJytChssPevJGud4ynLgPfBJI+rl+uwuj4dIN5beptnMpJuwxKk8vEfWSE3
56fqgDc7YdGgKEulC/LapNVCl5Bgg6Iku1UoukvcfA86zW5JKgyTVC5AYN4KImToWesl2vVnlLB0
uvoDW7tfFBGqkityq4ZEaBYRw/d6o79QDf3PjSJ+O0F4UAm7vHNEv38fBdGAuGY4lpXx234z0e2H
mxKloCKFXA8/QBEblPtUaR+AugsmeJSsRz5j7AdkCKVkDj6Vlgyxlm7fZuoZ4/qR9Nx6nZl0Elxn
P9NEmrE/qshUdu0tFpXl8t9l8KhBlG6m/1wCQ0a9EtULrhRtOAF9c91G432+ykabYExJVvelrpcl
veykXbl+VCOL1uTo84B8TbQ+z9qgIU7PIQzEzVsV6EQagb4rdjQFLkoul87eftUphpwHXjxLAchg
B7hfoCfUW99iZPzTl8i23SL48adQkNI9yiWegZnkRtK2qQwLDcN8CoGFIonU2a4+7yJV94oww4Nr
d1D9rjn2HuIHTSdfclwNEqKCMm6dbqHxi6SYDC9pAzXCXpuCY6XHSE4EwEWVGhs83GosB603bicI
rC+Zi59s7FfOb3MymtzQW0HENDubTktdPxirRlVunIwm8KvT/hWj4UDC7G7+hbutm6n+mtu6+KmN
ygIaRscNjYaaKyeoUmCa0biSdiuzcDsW4orLHSBCaDCYtLM1MYXH5o7C6bxod0lOHwz4pcy1S+Sa
r2dQ8spP2OXc+52KQAGGmhXAZorhHto1OJh9bT2JIt8LBanh+h3OxZYigFK/+T5irtG9Mo4YEg1T
7Kc2bRaM7KLG03WJ2lEzsg5L7RcbSKen2I1lRXaifwbeI7AlCNg0Ifv1941TT782jFsvPzkoP2Ps
u51sXpXLNIvmILvtgB0sByOfSfhj47FrUlt+dOJ6d0iyIqYKTkVqejLlYLp6YeJL2YTpC9JOeULW
xTia01WaUPCkVuOG5kjLqgoiO8/zUL9l7cmhx5NGRIA0fgUNUoH1hALiz8d70mcXo1i/KLKeWzn7
GjV9GtG2YUc9Oilww6HamFe64MGzl+j9/FTfAlYL8UK+lowjBPqo7GCIbe/VYSpmp63KkhhgYfJa
P4Jc9KZqdJZ+kHq5UdNSnw02g2CYgmMBc9oPyN/O6x0a+Sy5m2axxIeffCSpQ6G7mxpYknMW9B+y
k+MsdSMPT2eu0pm9aKLl7CKkUVZs6ITLmAf3CKIuuMS0+5Yxzv03Sqy4WADG3Nw8lG5ct+xTH/1i
MWNhfvSWqzvT8+ogqQgcWvH88bsbB2nYcsks0/ZSQ1AkIJCGtYoLYXq38pIcP8jxB1z4PlmD1Hsp
0oP5G/2ycI2v0ndYKUUwFkiY7p1/91FBlo2U9u1QC30AIPu4bcxQIErlintquamWMcCr9dne8A97
OjX+EVzxdnqsmmG+tJcpkZEIUfnf9mkErf5b5UDTnWgfu2fiSYhPgsGJHybQKnSadNBTq8fTIxgi
58hQceCE41oXcbFgw2PwCj2NMJGNfeeHtOhwfQhAtmzK9zSYOPuM0ynerB/gjQiEHuyhE9FRSaSN
/Kg4F34qKzHjOXXpjW5+23WxcYz9DiQfVboWRZTQdPEHTDvzSVrimrWjSn0+KTp4/WtB4fkiWwmS
AVWJtfPzT5P8TUiUPo6zg4saou1TNCv3O3BbVoYfHolRujjIOh74WEDizkb71sagV27o/yeyBT/6
DQt1lVSpLUxTgOPrVvEjpc1TgEPft7PdasJkH5hmB23qHisKcTvcZu8IPZBia8z/5TLKQVEyRU2l
iL81u+BObIfSiuf0tjDeMBnp5GJantor8PWq8Bgi8ODkoF3CXiOJAmpfcC9xAFBFzU3WEpvPHZtH
dbOO2u4tha7zCkOcIMYw+8qGaezdLPJ0wlrO93ETJwc4Srp3Qey9yeANCvYDKc9Cb+rPjy0JWybW
POSNls2RHMzMxxaqoDHGRILL4/mJFvKzQHbhZadnqSps2uURchMSFGW06Z6MLGZsGBz5CC/9DNLg
NOvAkQrAd7RSpuT1CmOdfv8sSFTrGRwgwz+/1gR2sAokXWBQKhtiui7IeSdRR2iNLM8X/CY+6V9s
F67gXtTwjlyPTPkiuyUZfHN9La8fdAbSHqNlpIQM3pXeG2RJx/GEvqJ10oRqyFODuQA5IAj3bhAU
29Uk41fwO2j7mkJZaPj/+8fBs3tNc3inqfvQt9O3q0Z9gbJakoFJ/a6TSAPSdVDv2h63P3lgaiO9
Al+xytfRzCTJja0SbJmtiUS98L65G/GoV6Mdaf6MiQ6uT1J9S65qNsZtFfl1m+QTxQW5atk6H1v+
JfopfJDfSXOXv5lmnGZGc4K/FXWzc51HmIijSnDrzil8BN1mSIt3tOdJLAoPWaDx1USM7h/I8WVI
2rQaTPxXaBkLNShTN+dbURnJ0jR6ISRwqMUhplG+qJWNnavTw7Si7cLb0IZ0o9cONxYt4sAu2adk
Bb0Nb/ltBC6g0HWsoq2mtQAoQtns22FRerejKipye6eRHEubhQobWhCd3EWy90ZTgapAGOuYUB0S
hQ+8xAvrQRyH+nf3zBxxWQWOhrGIZ5egJjkT1LwJ32nzUMzKsfRfeR3RUuEemHfCtSx9Ex6FNIR7
2nX+lYj8KhKjmqO6ha3rek2y2huhCrph3t5bI3tgdUj7jPWb52Rpp49J2XqEdYi5B3HqJmhL/v0+
sp0V/B2wEuu2F09BzG4EuUvt0yu63vToeloxMt1mdq+rd7mxQk4ZZLZhwd7UThHBDF5QPwBa6xAS
H+3UBVyVuwEtQMRmCOufJTrEtl8sL6tJ0MYao9ZwtxiZjSEpGi17TKXJlXVyqx6GZIv36U0YxxHY
EF2u/hmcuEf5IwIG/DP/Xhuyx2ItnBMu61GRFyofPCURFQ3K3iq/F3Htq2HOPMnWNWTMITGFEkcF
hOguwhIG8wrTrK4S/Dsw79xmRCZot45QzLHdd9vCTtkllLiRgz54PMyvPWdn1e6f7eBaz+nUmaMN
ePvfyszKLugZgKad/mvdGAzbgWPLjgPZpFiz/gF+5VRbRjssN0VUi/Fmg+kYZPH01ztAg26jh1GZ
VVpjMuuLDHiRlHe7uXhQfaEjLv7df/BhJyq22KhN6SkO+VJFmbqDpEHIwZ9Uyxghbf++xnl2LsbH
hRpsrWPoLUE4rfrOcK/Qpsls8PL/auLKJ/xcoQWiik4xnmqqT5HCeWW4WNdGSD/7EiQLySQZjqSU
JAzHZtHyRyaYrKSBVS3Wj5uPZQAovcKP6/Ab8crPCJHKPl5HqRvtWz1I41YDKtidmQ8Mka4ZLCyO
ljoyi0ydd64/18ZiNeJ8Lm7aMx6NDisIWaZY35mdx/CBFB7R7zg9aatOcuAIL0OBEGUKOcRsgw6Y
Jxt1AhT1qc8xoMN3p8PW+yLCWro3KnbwVH9O+yxsGMo4Av4JY4+MucYtIKxh8ZHNgIsRL9xLfHY5
gYwaWK6U1Lc1hpU6kpSvKQYagaLaCzRfD9xQ6xKRTTgWJbiuiqFFGN8f5tVpMe9vECj+2Q2ZEnRi
bVpn8ryD4vE2uSSqd0LJRRoqyqbBH/kfTBNRvJuOyqBgGWwjU4BIsCXCYBMOjWmLKQlK3D4Urvyw
9lrPIK87wQLNAx3f3/UJn26YVQDmayguMFXJCAd+SnZyaJ5O7kNqE7EOXptQ/F2ARqQNi6Tn5KUA
6FeIwYsF3WyQvhh7/c941E30zliDqOc7zQbz69WRLuLzFBLtF2O2V60PfLrQl1gbeNGXFe+//W9d
DG+AwJTpO9hiApNCAGE9B3WD3+YgxDMVJK9rZ3fFIVG4kSyG6Veu2LEZZk+hmD0fNnAjgl31xtZg
w4SYRdoEbZkLk0zp38krClQOwYx1mI8Z7IuKbEhP6fJSe3ehdfRaEqC/nm/6GvQR1oLCl2MMlNbU
wofsm8wg2Yp+uz+wKeCkGyUwZnlEjls6yQ03a1G6b/w8rP0DUx540+nZ4T0InxjpzaQzX5vum00j
5Zo+UQhfI33aFLiVyJgKpLM6YAFUwDcZ9u0qJCH1jGrPcjQxQgCuiKMraEaZE8Q0QOc+d0Nwh/zo
hngp4893vxkECvGnXi8zeDYsOUK1urGdyUBWqA2VBTneHxS1utiO3iJAKix84bZ8aCV31c+5TgkT
GqVrFcejh8Er0ZQtYoKvuBPn+BTJ22t7laZRDtHpTdBbZcDJsv20j1dl7Jg7iEE6YtcMrK3wPl/g
zo7aQq/DlEzJIFdZzJEaT62aGnKyODe6jsdJd+oX1/ShAn11pWM9i9iKnUtpbCMOF/18yEO4WB+h
yHMaJaXUDUrOu2dqPTeesotWkaeYVQhBNCPcNOrm68tSzQhpDGmUo6ae2pDLHDAKjgkWNPQrwtxk
ZpdxI6LAZZYTDp9CSRJ8ZKQOWHl9wTlrZVgZZwBFFIyg/5A0fB9cUujRcSLxR2vU4YCf9P47w5qZ
ibHq7c+N/wwXrLgHrj0Jj2U9HaDIPwnTR2oB0uT31VPy3B1dElfhZZGaqKVZssx0hgz+oAuy67hl
WfMcykU8uqvVOW3CecW8hmtNJKgebnjBynx9DZKUAYc6YP2yLNi/gKSBhSEpUEcmd1hQL3nW5UfY
x4NE5Ijj9Q/wdS8CnX53n2KIuoQERDhktHAsNm3trY4TVb5NLPNAxVfQFJKoGc4TvgE8+GpV6P0B
PAmuwOzT/U3eRI13mp6xFFjFh1ZZd3t3XGHW+qPUXNNhHLGBzh0PDevLUcT00m717WB3saBTCqmE
NEsTDH5oKzFzECgOhkIm0Fpg8aNmdPn3nP6TxiGTejyDlghtnIxV6SXSG/bQDjiSbNh1gTkQUyCX
fFfcDtHc1I37xezHglTcy08z6TqG8CmymM0U6IgTs13Vf+hcoi4nWI7wEEMYWX0qfYz/L7fvOxFv
ce9q6HMs2C2NVW2RRG90kkdpHjvwjOWyzI5BcgCDL5nLCIwCx0x+1a4xbz3d0gceGZy+lICFZQfA
dGwRfN8aBPLv2ATjwd84KGFj54959zMwirKb+qCsSPy5419BmY5T3cW0ijMUNhSQzRonibkpAfHP
QJHc6HnpjgnZWhQf/g/I56CqOzSrXjEaGMmbuIoU3brU1HY+xK9Szx/HbmY6KQOVpRg9ufvOCw+3
6GL32hvWka1P5u4HceH53ohmWqastslQM6Hg7r1/JQgyWJFF269jMuG7nyp/ziAfZ1Q7xfUWpky0
GZlytxZE67/6f480oszQa6FTqHFIimpsNourbMJByTsQ1SUFxEuEMcv465Q8ruAmUevnQ4MmAJeK
IuZ38nbNRsEZZ7MWsoMm6XhXguJZOkRVGK6QBICZclT1+U4cUcLSV/+Nq4kZey3N56pGZGExluP4
TCamRMR428LFB0dN+yRmxruwumLHi7MwoHOt9oAuZV6yfvvcn3js/2fudTn5NQQtd82XOQT3vDFz
mCvGFv/H0or8z37BMUWETtWukcsyHViBerEXm0oVVPLJ/4qC7xK+i8UIeTI8Evb+TKGPhbuhckKB
9w+JVvd5rqVGtpRPJFk9MUKpTDA3WoZpY9u9XQPB99ckyHqDKWvGMnd7JDXu7w+E1Ks/SDO7GzkN
l2e6U1eCWftBGZMyL09iG+41MMIXo+9tsubOz6NFwRFVJCZSWNcI3dYLYx4YbYM506awp2TLraFU
VVwVcq9bKfazi90j4pf/CPIDda8uHHk8Nxk2qmlDNOdBpQHHAPwcOAzKuGLkUFgBg6Jr13UVNbE3
1Df/H1E+DZanEj5UzK0HZznLbGh3RAlL6PylbIotRJrpbkktXvTUb7belKJBLkDgFqvYyKWYCYOo
KFT7n3W0KBX0rMWcs+8uJn7z6t2ImLeDW+wE16AJgTBnni/x7nmqSw5Ot8SoFn30wVMUXQW1VrHJ
EW6+R6HgOLyZsTbhRDglg4KH4yaj6HReJ8RsP7/6Lslmwt224FN5EdADryFs5djLjyr0a7+sGW12
gPSCblBgcFBGeyMX7u5KxQss/KdKjuoykToVt9UoK2cswKap6tDutYtsdIWrSwZO4oyxnq2mKJEX
aDyKoSW7VMxwX3JWHRb6INCx/wr5Uu6ks2jNawaPAVn8RTniKQW8Q0cYQNQRVg5no3xFp8RxPnJV
r7/y6SIOtS7XnB0bYNbE3u9JS0Csz7QCD9SulYe0Rn39IvRmPxtIUBld6qnB9911lFUWZtx5dIc5
KfZsVTNRZv12AHBllFPucg1DDZZvaaLHDW9jHTTLI0b/h0IZW54KMc0eMy1aDvCABFW4WioxMNtE
1SsLBMCBGdhT0bimacmFgRuZhS3QsjxbhQBKe/EyEH2nsdsH9XLhBmhDcc2yHW5gUICjhIKmjaye
TyGUi1OrIzdch1sJ4J8mv6rQ/gii1kBAQWFv4W5M+EjphOm7kRM4qwdES48pd7yErd4VdVKgsKhp
ye7b2UnhvJeFCLQZxRrTRJsXC3EVtuONXpiJF3bjDb0UOz9x2byVnIrpSTXIc8rA3M+fujpOeE0C
D5gpGCAhpZZ4L/dDxaHLX68vg62BamYAPWMNZMU7vW980HllAD7tohCpgUEp168jseGxEuIiyLgT
AAmSV+gAHGwTkD5h5aCymerq7THFuCM1G2YIWiDdpE9i+AH7FgLScn5sHwmcWQY2A0DLeQsAjhVK
vRdIG3PUltpD1Ynzw8ZgEDNJS+HTsKrfyoBuneGGAtxdcGYVCdub8SNremRev/Fl652wR4f7jLtc
1YDeRD1ZMFCd6d8OVjeCgCxathMuoLp+NaDsrIVDK4bFjRi7NE0U+aI25QkakYtpfIPDmLoDgBKk
szlrD2aGwuXCoOKibAvIto+2a/nqjdR1hBmYDPsX6LyE8PTgGF0BI1liZQ0hNX/NUTlcsGfTehaC
zHsvii3jHPoiJsjI0Wzaa3X6e0R9dE8NDGyG5SgiSmaN0EBedYdSShEcf0Wfy6iejDbwLy1nY2vO
8KB/UxBpujJBk8VhAuljnl/jPtTHX4tVjFXsQ8vsf6mYXzj2wkncvMD3G56P0k3O6WrjXencOLag
LOlUAgwWyUux00ezzXWhitdbpg8bk/uI2pNsL7XVtZlqG2NiNUlKghLMxfPQ9mcp1yQrx6Kbu9bn
+5D/IsCZg7FsDYdMpSng5v2QM+s3GooV+8LsYtlR+AuWxNA4C0LX5jy0/V0nyU7pjc3xenBAPRqQ
qnYSOvts/RlDI1Hw7en9fBTn9XWBdZ0LoytWMfgMaBkMbPZxWVBMyq1QmZYmRfyzT9MROuMg28mX
1VIIJf+DpPcuJAml3DLy4ns+/s+0XT/J9umT3rxnSYY3Z4qrEraMvW6SjfnQZrA9zfPH4zD2K3kr
Z+HbiwFJU9CMIeAb5UYcnq4xM6em+1zPHN8Et+WDhtKze2YRIv4UIP7oJbLLyFJJzAdY0XuRLbSx
IxTcZx+dYJZ616OLUyCn1yjW+nyQJfgvl8OipLIBqYAXVlssPrWx7XedDj/m5xzhKwdUB2uadXKY
Ed8ib24BZ4nSEwTe7MvSfWKs529QYDEJt5G48RTF9wYPLoBtQo1egoPiTCqHp9C6cV+0UdykGDoR
XYYK3+MQpAeP1sVWCdIz50pW+/rR/CmjhxEE/ECTgwHellF/054xg5QghBhmBNjdXGq6ZNU/+TWx
tjDQ3tiwwcMaLpSnwakzzPrG0/M+XbuRmd9InzMpHypFgurbu4gJYtd+jmd2mLDDwyqZGPJdyEBA
zLbmKVNPjLWmpaDRABJcR6ltBkTjzl5MTERU2dfMVgHtyb8Q0S7/a1FJo3D1KZxmIFWoSo7LgxkF
IOcIDQQXF/SUF6gv6vGk/omiQo0xB8xq5v1u/0i6b9HTtIDdSslahL6O+jk9WGZp2ws+JBddc9xx
gX1ybpL6vFluw8e0nSfKaoxn6QdRqQ0IWyMu0bM+enI0KGOfBi44dTfFFSxeZPZ7bYE+0U83Zo6z
STDZqzcUPy8j/g9z1gaoY8dr25Azvg7ZicGH5TmAiqn71hlY0EaMoZRI+UFw74c7JEzWxNkLWOz/
/+xQp3m8NHEy0MZ2Utw1ErNH2x/qAfnptPDei/h6tc2hOxvM8kHt3RWeYdL57kYyH93fbRD8szer
DFdTQn4m0U5m63vsh/Owxg2mQALFPK5WY4A0USh/IfPUuFqhyMwwDQwZBC8DtJc3+BJqGRnYKq0O
oBeF5oXaGrw8XghMA7RzQrOZe+KheO//QYdJ71rs6ZWgml+OgM4umS52FvsUJY0Jp9CKXtsjY3JF
AhE+koZGCTZvocCiqiOhgweljrzWGdBdsrDBjkhyUKaHeqHP2GFqxY/rzIQkz7txp2JkH5rNEU8B
SpcFBI9GZtwLDfsz2mLG2EXM9hRkNGZD5pqXa1qG76JFuMvCx7Pc/A0Xju6knuQX3Rbu3Hscmxas
vNxFD1a53juO+8hTmRXmMQ9Y1mWnSnMJMyXD6Fvoot4b0CVDJEo+vktMdL1ZeA6o5VDzoEctPhDS
8lb9gdp6liU9jWwi4nLwmyoFRrE92AnohCQm8tm8oDnt6XauSCwHsoHARmncMmOLlgWtDXUTB3Ou
OfXhHw+mGbNFQt03jtrrpr37lGxnaY+Cnh0E4uiVvJkpjR7KpOG6onIUGJNdy7LKlhhWZN1Jqm8/
E8Q1jayUzu2LdVQmsfR6wTrLsvwoAPrEnJPSigXvP6qbk+DUVyIOIhXJzHtKcBhMBbq/7VUuMwqs
pnmRjb9sDRiWNyRu3D62BglwmljvVqRvX+40/G7UWjfLJwAUX59faHToG5mos8pB1WAxL2EIJOWN
cZEH6uf1rrCr7HvjuLT68LXXE1wZWK1HO39iptm5ThDyj/o3rX18z0KllEGDewLvDMPKPSXGELuH
wHn5IAn1lBXvNHPPrtHh0SEY918Vr6RRdGhfmLGjQFP5kERZeb63HZnn7c1mrtgKSFQ2wqP6I6UY
n8a9apSoEvn1IXWFj+7TtZdier90kKJ7ynnfZJY+TDsXgR+9c3qHGAsyM5now66D2AyvzBI9/vXW
IRnt8VYdq6W4geyXbUzaufmXHJUZJ2urOdOA+FjnhiM/08Q3TuYiGiX1NEJCaed+5yh85Hqqp/+k
OCmE2YwOi0PpCMZAQWKZwIDAd6yMIRzdF1Spqp7vnrpHWE+AsyAl3rnJEkDjfI95lNXziQV04nOY
HR4E2rsZmPEG0QdkXxZBZOpgdqtRcL3NVjiWBlfePJKV6narAiWXcn6fswa+DuIpsEtdcVG035Au
ghZF5Q/WdpM3m42egAGRZxpxuzj6c8liBbUqXGWBDMG8uz0tSxdr1yMtIQTyG2sJLRkrm1CzZq8K
tlTPrPjTRaSGxFsGyrLNoX+HKpRTawrQN8JMvzjGyQUB9Yvp5ltOOIJXvT1US0Q40R6UVbu52XRS
33LdgbT3isUi8McugMC/EnP4KvLgOPCVkgVT/eyAqc7D1OLKLv7cqsL2wS7sIzJPtQKZ7KEhCI70
DA1g4kVDCjGY2v30q/GtYwBIpC3fmtYtNpnBjivG0AWvmd2P5SrVSpmmWBhxPfGyRFhNx81B14VU
FzeGHDQFxvmWfcgCJzWxIJEHTHGCbjiMu53Ol8IN+oVe/uQf14229vSzX54qEoS4f3Q1dyDD4euC
pmv1VJON9s2J6szjJE6UNYqB8t9+sEGHGIrDTPw5CT5/xy7r3Sk+D1VGgkXdTtTxDwkEEQD9RrjS
6Xx1q7W0+qcqnVjximhbfynm6QRlwYQ5PxpA/cbsKUEdMDqpQkgzdp49cWMNhnYGyFxPgXSXBK4c
SQpqUVONArmqceiQ6xz9v1jJwolmprpzNsW2VdVdu2BJKBnATRnVA3scyrHmumy1zO6BUSLqt5Gu
r4ap82SPU/a/J16YIDJRTW4yyue/Z79S2Bw4A1Yb6VhouHFiK3RlSohfM8qI7e7/X6cOewe08Mko
hsYyrXqKqGKaZ6iZcXexcNgtYxN5fnwzgetXrVIIan6KTh8wFqRjSut6bHRPzVq7revhc51FfScV
rotPVLwChpUFB5tsiHUJnmfCNsksNq2JLswA0/d3AyNjnI4eJI61n/tAAup+Jm+YMXQL0NFpknVj
NhdatnbA0lyOLqN6FflRyPvXZNdueVM0L07h2+m4VQ58LjSmIp6HoL5RKeCJI+UK8bsc7g/0E7/V
+Sa3svuqBox0sBtZMnx3jHOfz87niTn2pR1/bSH6mK4/IErWmOSbv2NE771DQpr9Ua9Wg9cwUfyw
GI8UwExJNsSBHVdx67MWphz5gwa/W/tWGiU2Rlt0dbiDkI8GRKY7Cus0nlLlLwu76MFMAOiAp2CQ
GHFyUzmODHgKBjFJ1UhQBhfquvSwZ3jmmizkHiDFNa2oOJkMp0pUwMospLer17rfSOCZhXWzBKug
J+EL7hX4vO68Gy6AdcAchoGhbjyMdzEGPgHEWYMA3txovtN3vxWyAS7sbZK8LtameVCPHZjc8LNc
yoImqE4kwaIZB7D66y0dYqvQrH8VbD3kxvvHuD8GrwzaRiQciNuDUR4xGcNzoh1W4qsiX9x2LFjp
IZv4wU76xr4++6Ef8oZQJ1+O/izF/i69cJe11r4u9iqJYNM9hQbcVZqEDAESPJTCEckXwENDEHu/
VDUeDv+0ugIW3K7qDeAioworS9kH3ipdv/leI2+oPqeIA/3vp2p9LunCuEcPuSXu4GvKHGd/bXTM
QX1v/T9TaoLFH/97MXrCjP+qUyrF4aUvHqbEWdXFtZ7sXBe9lEra0U9xdNMCDPmGQeZHfOieaPQl
wjHQambj3Sp2TJZvyKFlxjAqPb2r043d7hK1+srbfrJbr+cZnjW7r6ciNUUcdPSyL1eLniJ/2WTp
PtXxnNO+AGaP9AaOjQezPw3/mtsulIAeMefEwaT+ERj+ppdvXFuH/DzkxMcEC0iSlaOQ1oVQQ40T
rCKcrx+cGbhLreVZhnPWTs5qeFNhmq7//xXfxnGpYsUPOdFGce+7oerKG/bpXIBhKbklIl701xF6
2Pr+iN7o+ZUs6KYnpHCZLCQ4jp5RT2PNxMo7iCI/fUdyuJh8BLPLXCriQtlDo5cL0n9lzMtud12I
4/xKLS0yAWeUwsEoEpuwhq5eIyZSnaFN3FytivZeLt0hu4s7HxKEvunx9KVwqDE+VGTVPmfAyEub
xB++3ow/+5CsKHQrqTAjlQoMCINCWRCEL16gu6YDXZxKziM4IQ9tcYrkfhntyzerXCWReXH9jgfb
pGKaFGaqUvXvZgDp5yPwbZmjdQMyR7w7Ml+TEuvlpKYJENn75JAAy1qJshwNixTULeJhgx+eDJuR
CsxbJSPzywmOyxnA1NSe1Ro+Kg6VzDL9FF9rSJAxNUM3xHM/5312CeU24aDnMg7rxlY/cA0kci+S
8ixqG6swRctamRVgqDM43Hgc2sz1aSrQnz2sCiTXrVKbtEWIJmRz9RJ1/b+QyZnWKX0FV82JbeKf
2RcZYlXGMlAjKAf0eiFv88O6J5GY5hrWPWosx7pSJfUvewc0uaVR9tjXOPRa6ACHOZj62A6xTeTY
kJRmQWc/fN0YBuOFfDFFVqMqxpbeXO3+OFyRQeEAJO5gYxQAN3X9hcyXQsEOhsUtUfdlJ8iteQ/t
5mZJOnj9+ekJcRlj0w+I/rgUCB3iSy5CR8QVrigrde+IpGgHCjTkLgnlytJ47bVPdWRKKDn5Gg6P
A3ThdY9TzPmYFz9BbnbF3YK7sS1BfG4x3+YS2OyhqZ59CIyJYf92KpzVPrho9VoaduZKX/VxBQVQ
GpOR27LalOza2b6Fgza/vE4Xq7+W40mllxUZQqlO0gyF+qwT+lqOQrFNADx7Fy4WxjR6coWEDgIC
oFclb+B4KE2pM4B3eQkPwxYeGs39DC+j1bfqKRNQB0wxDjElbzaKd+pLdASaGalQ+TE0nH9Xg/Ka
clCV1ZUAJasHopHEIHquqwYw0qwfXShBSp26BmW6NGOzu4OGZ6oCFsRfQc52WwSLNBOnXQWdJXVA
nJ3f4UZjUjTNL+60LKkcL/0/TWq0BcXK3JBlZMmSfApEcumLN1sSEfV+42J6EJxdHGNw58Pw68oy
+pPF5LfsSAobO9feQj5/ymXoOEMgBT0idBeAX0mL8pF2+t/+5UuQ5/tHdBCVv2vYxAjeuTm3b6Gk
kmM6x0JWpRGCKiBmIcvrF5v6kDsJFBtdI9N+DPk029GwdLiUoQmaB+nnkFt5EVhX7MdrFz11JSh6
LDbaEmRMH/P9dp4ctFRZ4W8l4VbkP3O8f0UnTgKAYCSeEKCeyGa3JSK4Gtln2kJaKYsuO5dS9DOS
rY9midHhptRhpyNPLsv5rNqcRFI4Ml0WP0HUttYCPmfnIbXLLx/rwyngH8e6mydssSOyQlB8/sCN
tYMhS4xfmhame/HE9KOK6KA9CAFhZhSlHePHJ8+JDHWzteMJLDzqkXtQJ8VALdyj3y8ybfW4RNs2
cUjeh8SJQSYKAwdrQBfeE6lWQz9fZeI3L1mtYtjabxcDh9jtHB8dA7k7bT4EeX0FIMz0p/rVejeC
Tl8E7fZKhv/Q9RsLvn9G7Vc35QLl1jXssRxyOG13y89mGhv9pN/kJQJUthVC7UWmwvEYoIJjal3t
SNm5+BDh6LG3TTLO4ktzKrHJIfsl1EgGjVievlZmIwNCJSP7G9P9pQ+1YifROYv3ymc7np3OScf5
rHkKnP2ebDOi83xAG55kYg0qDrvKj+GXSKtPoGqqkiRpWmCIKnO7954YCEJB+PASlJMzq7dFRzfB
uuVnsNUVvDbpeabIR/BxPOG8XSGFQnhA4Xt0sTOOvXpKXBTpY1itJofG3ND8p0+9zV1nZHLwW7GA
gZPMVN4KOcKF+1jL0jm9pIKh3PElDAu1JYyzkFD9JsfIqQW02HAyUYwRL5/fmAgU35SKFoq6BBDM
5LILb0zm0zHgygfORnKgY2AaQ0HbaO1AxIYlVL0QxmSHP1t3MKhraKk6M9isiTuCuT0g7oB7eNo3
LHwviB0XKNLp6Y4Sq4apRpDxvXeLaoN7O/lEnV4SFuj5wKm5YshjXexGn6EybZPILhqwlXMFsVxi
i+42GB/joOGnpbyplczkTjpszw/qwO/QNHRE9R+87c9bGkSZ18e6UDktHL9DTd/riJM8qF5VEDBM
hHA2iV2Zz1ZANm9zmBSGfioRdY9oPKP0qRHW0u5SZCLz0KaNX2p8w3tf4lmsXB9tji4CPH1TFNdt
TitQwjPrmfAX+QjqtiV6WR6LnY3ILmUn91bne9msHXEKZxJvlNx2UwKEWqDJNCTBdI8d2KTEX4ET
rn6/3PUSR/qzPFaUaHQTPL/qy3HRJRVooiRmKa6Rcu/Ar3IB2vchmdXMfrLOhfWV4hCwJj351bpV
yvhm5x5ttwXuorHXQGeZiJLVPjIMHMo8DP3KCP5tTS8R3hSPV0spPhIshCKVxIqELBZ2VApbdf7p
fe+5pWLOz8tZyaFS6jOBQDPmuEalTEHgkmqHqWf7t5/0zdgEhEMQYObV2BVBT2ZfdZ4LjFqPKh9f
blcWdXt99CHn/bf1ABJdyOVrJ9n1OEC4C06r24bdgG+cKQSgx0szadfHahrgenvvqeZ0graNmP8h
eJpGXwK9OIONdHFA70z+ZjUSH0/WiGnEgYdHHIfq036QkaF/1ibj9ccidPDwFUE+TQt0hxcDNRdv
3RUI+/Lyho+zTabR0MXzjMjeCWBNfC8z89p0NugYaXhMhVjrdLsI/hecIatIq6G8mL6G/hjFufO6
gEr8g992qo3jGeYIpCQ7IBlO/NVNqr2+a4/K3gz77VWgZ5CEfT9n2V0M0BhgCSZrVOOVU/pLKcLa
5uhdYf88hpsd4nzO2Bvj22l58yQszPaW7SnhytLjbApeWnwgv/0mbGi1CKsv14Sn7fikg23IsfNT
hKKg8Y9yLcRLLQd3QPJLtSnSogmR8KazVm6YFufRRLyuyYe+Qv8QeC5buq7udM/2ZAjVSdITy+Wc
c4aFuLJtaY0g6fjgYuIp39yuXf5vGaCQV6NR5bCspmOyFgPIL3eLtV84heQd1r7CvjByf+xOGTAz
TRDmP9rLj4cACayXwK9jqzP5ReigrByO0r02l1J0lLPwuBaeBvj31xXq61dRvutgEzX+tve+HZE7
Gn61Yb8ZdQULVaDw0SovjwVBor7JwkCGA0RJ2O5c2uj3viNo53r8K7fO8Ff3Dp+kcUdvWQq1Fpot
wQzvlOHDFXKHMVKReZ2r6VF3k0adlntajNFEYSmJat6cRc0mKLm3ElvvOpS0ktGq7TkifSWe914p
9F6b5bX9fPopgtwGuZTRQlGsaPcDvtabPduZ6YVvpUsuSzirpvVCRIGLk8HRE9sRU7bCEWIZc7Yj
IPMlxIIrOYUV6gAobsYj3uEJdMjoaDMNJ+VTwgzINcKxAvssCIm13bPLCMfpwDzZGAqNPQlMSGyl
5Jc89gbpum84AiduvIlCs4/5Jq0952ErE8yODES23w47O8ngqQLN6ter3L8zBorqSZYKdR0PULML
LgK85471e8iFQtY9hx/3qTiOI0coV3+L3gbD67S138uQzINO/XHGFJFvJeoKO3yxDa2wgj0Q8OtS
HX+SQf1xPC1WC6FTikCGRbxqM9dXwl8Fq8whK/UNbuCaAvCDBmBnh2q2xRbwzjWG7otZXvnUMLwG
wEoaolQ3Q/cU5WCIb/eu0gxXfdj8lu02Rti9w9VxiIRJVEBZmfany+7Wi2BrWHcay4+VgMmCTBPs
KqlPtMEzAgZQdD0w01AO3k7huoCOqpAMrGglNe/BTk8llyW4jOuDJFR9+5dAa2tQhwf1EUtt0ZoJ
Jwwea1o9i9B/4Wfxl1VJhtNEdtqdRx600mZnHdQv1CQgsCcFVfCUAsI2vTKWL9dMOmjtE1RYPaW/
vLy64aQ8ZHns0jPRZs9Gl8n/e6xyCKRO3yrWTCi2i2QH+6ELtocc4UYjBuDXkIFyH2zQJxCn0afV
RuV/HXTWopotMjErI1Q7U7R/YTkmLFbwS2skB0Lpkqfzf2hC6E+7z5jR0gmRuwSenb4pkPSeVKZ7
YmvJKJdMFYLillLYEU8jy01az5ziiV1EpAjkepD5xmFMHZUrEaNbHSy2nS1qZQvMhhZeqrKrrY24
mJyUJ63VkCRt5GzIcP0qgai127f+IwK99ZfHpOyWwQJjeviVcYQGy8/+gOh+qC6S3WCOHgxNQReJ
V5XQ0eKeZcp1G3HUGOvGy4ZlB52A1PcDu4FXMbG5Fgw7o1JH1NxAp2sJHLRSK15usWAhcy1OEpur
unqPvLsWi9Yy7CE/lYMnWAfNdIq4rBW+eqltqFZut9e6RNl+ZwmBhc9FmnXnKINFLCkZVUCGn1qx
MfLrSpjgTI+ybzTrKbRICWzadNj+jp4YZIgQiAL9TVaFB7cuhRif0QJzX0BHSXWP42GiJLn8qrY9
JYWpNIfdzrWxO8by1QqnM5IRBPkxETex2JqwunjNKlckhtaX5K0C3F39sDirftnkNGvtd64rQfXU
MMcZTkAZfMIOejmxQgmAAoujw6bzQGie2bhMvjiKnWqkxGBeIzigmlCKiNJ1ScZLaCLOenJQEIOr
cgwz6782FFBYZZrdDcLqfvfNdeJblaTcvFeN03tzm4AwHkwbluPmE/JemmYvlIDoR7sqGlIIgwcX
5MOr9+K6jfDp7nrqaNL99sx4yip1mz5JbBHk4EBOmH2+etAgYXnJjCUeV36/39osEk5sU9DST3Ir
Fwjr2EzIS5VWSr55cobph9ltiY3dCZ41OKiDn8uteI2wT685cDmF9LmBYiSI0DwliWuedpsZ8tqC
Ej6izOUwi2hpnF4omJUDHmYBQu5lXAc2V/PjyYo/9eWW6c0c6bi1KPvnfE0t7pEeam+g0bMPYjtq
yT0nWhWwz6acqOmnFe7KMAEjmCtyXJnbyne7p8MqjRsJFXgu5Mli2+ds24lJ6ZutYFHithnJhlmU
RBQCsd33j3udIGGDpDKPvs8iQxIETV1DaRVbvmQrB2YiHDAjehKY7nXqXquyd9rVmlkOSPeyYhT7
hesU8DLTx53q0KKF1C09YhVoq9BAvD6IdB8gWqH0JY+DR+lsgLKWF8gtVeV+7LenZrDcjFhLEOds
tDmaiERaA0pTqWwALhR47IDGWZcKPZzA4xOUtIQlhGrDv6OGcHvYmGzWdLIEe/sXeaf7LFopy93r
/0uJqt5LLP2yX+1P9gQSTqLkTz1aUJ/FXHAk6CgeG9sx08cpGyD8uZhR5NNjAxwkwDK0FBELVaX3
J0mabcQiBeDafwMpDA5zEGlup8ER4Vk0P628ZagBf6Rn5F5XZJ0rho7e6IllMd5LwPRY3YJfbYJx
za8sTPnHxfxgQl2uLAygNuNMwsnIRNkBH/dxIav2ak2OvWk5sCjEDlCtAa7eCQiY36GsYcf6DHfs
Oojuyy34RE5iImQp1JCe5HvWYSo3Q0/NhDhrDHb+ml+voUBFau2t5UlxoNBWmi3r/zqm0fZ6+pNQ
YG8p+38Ey1xn5kKMTLVRKsEjbK7VmHyXa5GU1HBXXdOavcNq/l+K0ro1xGZ+TrFsNaxexBlid59p
Qx2kGg4Wl51Uil3Bev8VEuvX9RJf1zFTsidDDdH7S0cJlBf8SNl51n5bIPWrjrw6tw6McjI6UaYD
VPB+R8+L5rxMrZxqXf98ZIqrvn10kj4CaDwmpj6B/2ZqpPb3coOfehfZdSs6YGN0MI7N1/Dbldwd
5PYxcDYX0OYZhxidArKjujzecsjx7brIGiWJSG3vyC+S9CL7e6QvevcrFBM4YUzbLxARKFdGR6Wo
psLLFstZIRnjQwiC1GoT1tCfETYsypdaGWd7gVnay/vn2/A1BrzLuRMDWBrQbxRSI8DgJOJ26Dvo
v1QyCk9teU3zdnKuIvxQTN33nE3442p5Xu7umzcxN8t3JEMPXb0qiUWCCqp7zkchn6VxgkztOFOI
bpd7MqpIiLatBmYQtwUfQNmy88Jg5dJ8nU+GZebaUDRzwuqyruXfAsK16oy5iJTHVlonxkwgKlxO
q75kW30M6WLbYRJkrH/mm/qhZ1HPFo03X1rF9/DplJWk1vYBusTHkIDE+jFJh6m5+PKmOu3Ep69F
a2VQyIVPv/DP7phnpY1HkCLarfCN/VpjJwW8tpk+80FMVqO/dRd9dfBGmqRTCBPLabX54fgU+sCc
FxLvVykad7THJ5ThFqayEZLuUeqZY+Q9UvwT3p4LPbBBtT9uaFe21Hc5p8Ll7HIVuirc7kah42VX
1VNzLqLwJWNkHQK+GNcLxgpbra3wb62rLZSHxfVMmgn7Mtuw9JrachwoCiTa17Sg46VorxsM0wAW
upcr/qjHd2E99UBGMmfKyBph3goTozD/H9U+fbbO3d0L7G73Osa74PSpCmqUE5VVfh1hk0aVa1Gg
8vLWkyhu3D5uzZyFo3c/6UKxWZ6WSW894jSmywevI1hNcmZCb4vCMFgsw2HIydQjklHQr3cgJJk9
x4Qj19cWk4X3yklCmsK+x0n2lym+RVPdyOhoHeAX9OIPxE/ng57UdatbWmGGS324WIgwV8jj4nK4
/wZdMAUFiSTgr2D+mh9+YcGJCgwX6PKFDYF9VMXCtxNFhb3vKv2RTeIrjD9XNSc5kA+hn4pC4MVt
sugfwGP1rYAaVS71K42WIr0Yc3nMuyk+dB1GNJZL9XHrMXLO+x8Tgipa8BDshHMvOBVZv/zvkjMj
T5eXUyWz7VZI5mHcVIwTm5mdniF+2idhnZvQS40E11D/eeQBIXJC9bg4HLdorDflWwMta85K5WfV
xwWD7r6LQgCAtex5ggXMjfZyhneuf91LO9SdATUitdIcMy8ruiuuIazEuN1hK5Bq2wEQ2RytQa1O
dwLT4443Lm9iWpVlg8+44ngkmx/gtpd1sOch8mVuT41YduAswrVo98R1NjxlQ4vh0QQOXoWZDwld
BwmYYg5uOodp7zsv7YvOHyvElNiwrBYZ5ex767F3Hjtmbqo3j4uZpGZsMJEzCngs6ty+gHLsrOZp
miw4F4gxrHF7KthYRB73aGTC8eEJE5VsIhLM/UM2yfNRtJ+8dckXW/Y7jm1q4FnOwJUd+B9mX8Mk
2l3oYojbVkJLKFRdQXLhDw/dOvGSPziXNg7J5l8Mre4NS98kBE2KRI64HZvXgtr4cLJ4bZsfOw5z
VUDdRpJtdVDGs4/hAmQdcGV3h7fyT7aeRmfdanL3TfudmqCsdO8DT+D01mMDne5+3ClXyMh1eFKN
1OhXzMrov/xLEdT8w27VuqYFyo6CPz3eZZ/WeiZ3UHYaW2ciB3lRWfEpvXK/SkBnUoUU8Pd6lTNX
+0hEmjKpqhlWfdzrW6bPzS50ZygF/TSPzSpU3g2Va7AuFD2KlpB/Hozo5YBuygoeoPZBKgjaaPu1
3q3wWi8LcQh7BL/Yx9hPqx/pqaKmtFtc9kIXd/lKe4stwjkXYZaeDMeOihlnotCxkBaNFgZ4HVaY
P7OpNxNPTxL4i0+aZsGm+gEvb6ApgNxFRwcQguVqVXBScE5qsBBHfUXgRjfhos587Q9Fh5d6gXn5
H2fkTh86GIdGIPxHLuDIDNMnxN/TZbMzjJg7zOuZ7nHpNqCAo8ykAI1BerVNsO71/XQNe98dXpcC
O2YQ/Tut3bM9rZ4tS2TKzrquoLYrIxR39mV73nOm+0QiqJpWniWEjO22gFd4EUbaDIgAPvaGOjWS
gAbrBph+rQm7qMWVbgiHfLBNZu4IJgV8DBzYA8xvGUUATcYxQw6mAuXYFPeTqTEl73fWu3dSE2uD
jdbnyM8BDNdbqeX4f87TUvQZYx8/RF79jgnSZ6yPLNvh55jfhlfavvZlH9VVmQlexxNMPX+VfWuU
RPXXzd2P+2s72LrPao6QEiiw2cVBTR3wtEyWZPnQupNTz74W8MnNpQqi0InLBn0ee3ZQWWJ0qbmd
LHGEiizSP1T9aOtdg5MeuYlHMp84znf/raIoHcf2nA23ipUPpeLLsTZgey4OWDOQO7cOrj/aqSjT
h9RTbM95oyD7sxhOq+cgqb83Z69Dgsla6Wr5NOHkGObOzhEtR7uwgnhRNfU9Rqj5L0O6QV+OEWu1
JgUbpGf40qB03sJMnfjjP9qdITYX9u6O3x05lxq7uFVdQvJiigKoRmasCbyz3V/oen0pGUy+rWJn
W4jr8VYmsC6yapYQIEAetDR0M0bleJy0PiDiRuHzxMsZLLhG0uAGPUhbiLrE5EJbM7CZcwuIlSrc
k+4wAbLKzuPy5q3aKl75hp1dMUVf8xibavXzH6r8UMcUUwBlHYI9QudOKjL17AOy7Z3q9d68FeY0
6puET9pz0ACPblDuIM4cwMgOHBb8x/8rJ9l2ShvCVBh2S7fHXTulIG5FbpXY9x4A1urmIbtH3dPW
ILdbVMuntgGJKNZ3ya81fcdyTAY7toWBCXqTjeHKCqXFsR4GZt8/31sJ02GFxN6Wf8ARK+em/LGD
T4ZXWlJqk+l6r55L336djj8SpPEHhQQFf8Cd2oOeivWd00cBbgbW8vHePLWml+n3lIeh/KgdEt5M
E+3lWO1CUymzzhgGY7Bj9RM6EC1IeuxuGg6XflXFm7WPd4MGq4e18VCtKpjE9jFaav8+QAMFrwOn
shadqLyst1wbrLIrYYyBwt6FT04xMBjtzaOKUZ4qa8JwrPcBnd36kcPBLraEiMWTUboEUqiSTkEA
ASxkBJWix+kIm5XtextVsSrXLyTk0zMs9mloMzab0oI/K6LZIRf3hu6ThKq0wx27SAoXL1hHosqO
ylCFj9RYaFEl/CE/xKYw6fLTiWpbq9zbsFEKTbxGbQMLWf7FU9HJWVBEXSv+sI7TpebCsdgN+QT2
tPr5y0ODLNXJg6zTlaPE+/I43nTmgFC4gE4lHm32Xd2pGEv6idk5VtjHdaEfPpA+BvOe9g4uHQmK
TZPCbSqQQ37igijDtKzKvCfyFl0k7z6Z8Ud95GlvnIM60YDrnPkObUD/4gq4hERTZ6Ys08IaCwaO
Z/PvtradJPTXx41GADo0+rStxMabdBmg6DZ3s3OLwVd7sNYqoAbXzAykeb7pHKkusqidHOPF9YOq
mY4z1vs17lWVykV+xF6GSKwhgsVStnhQVGgKGFrNT+GroO+wNGku0SYuoARHUZqDWpl48SyIg6vJ
qMQxY1Vdkc5Ophg31gYUGxihbUWJhDClay0mfEzSRJQsdb0DrKYosV+1yqZd29eNW7tQ2CGNZFIT
sOzogZ/3CNnG+6aF8e6zoOxFxNdoEDe0z9tTFfAgk+CWE7xCUQjo2h9tQ6rRAyEMJzGrLnTTCpu3
36HZhsyfD69Hu4tIOsO+y+EbUn+eFebpSidm3SFCUBIQTwhScavAyVGTYDgyj6bD18JON8s8FFNN
IV346sMv7iWBJBjlVMFAhxPYZygobf9/YLHt9T19bU+Td9I2BP7qhgcuda8A4HoNsk6AbCYpYncg
xz5N+Aa2xOax1ui0/ZUlO7zHHonPbBV/RZ4KTUKiBq2m2gWfh7+WsjTFdY+5tCi6GiVmjfTpes6G
8hVEGesMvkDnaW7nykwoEz+CLJenygvqk5R6TsIun+wUJBzqCrRW10OdgfIgRtX6rS5SexyCREOi
mAu2GRO+adUX8oh1nR34SxMFi8MipM1pBP+MBwAXmcvuw5ymZ+w8hcxiZBr3fGFp7tU8S69GNZP4
P1Y526xeRbRuxTfka+uz+mR9vPv9Ji9AVpYtdcTCZpLeFaVMvn96jKS3f+f22gFj8RcebFWmlKxe
01DSMePLvGhwVK1WiSR6atkJ4f2Qkvo2AZrs9UkpTGYT3PZaXLq0XQ4AuASVwtubzMSWuZGcfrG0
VUrBArk03sMO/zwdyZi9G6IRWCMkSXCXh8JlKDW4N9ni4DPBtn2iqrJpSCJpX8u10Tlf8hiGbzn6
AyCMqoniHs/jZGcWDnxW8EVAfWEVwKPZNDAYuyzRYuNCknXmHdLpJtWKGjwoRMot4o+JmrSyczGo
l05J64vkYfYQytwWk8rZHg/TKENk3ThOHdsh4CZfw4mBKfjGZGYctaGWPajQLrpOgmQpIishyY5k
Ny405UiIRDiJfxgM3TpM+F8oZAhqHCl/OxcZVYTRlbYWxqHgBDXGDDgr2m7mwPa3lN+TcL/pBgi9
KlIIBcY13QJ5oSvlgqV0N84wpqldcub1jVN4F11i8P2E8c7IbOTaMMjPPplQ6xjdqcmDt4zckmoC
umJ2dVmVTDKNL8KhKvVO9CL6lZIZPRpzsCnH7+2tWl3/NBZL7QN4UyLkEZo0GFqj5NPFxY/RjAKa
0nXYYZFlgGemF03CLbzzHrUGwi2YpZxurVNIevsiiEnTOvXnUDPANCMY41i62yjnTYC3nM+IIrWJ
VPjzVhAeFsBSpIyOBiRzCLDRZlaFyIgo1tjdoyNGc2QuNFIRTVqwNPv3wt+0lN5mh+QXhICNpLSg
mYSFmV/Nn5+MSV5tvRXkA+SwyBKcBVnh8vpFOMS1n5k7vY0a0YAQC7o4QFssNEUtImIeTGRuJDze
+0DWq4+3tAdIL4WVxLC1uQer6SnM2MBSuomKyoonuwaZhhQKbcNOkgNHbEmH2SzkBRl2jhpFcfZA
Q6pmjp21tyUpNyLAP3Re494r2QRcZazscRSd0ezpUVMZJbPZ0gtHMdgNer0Kr4jbyb6hm847ioAp
XfTjRuXwuW0GiI0w7LDvy/66LUTy8ViE0XXtIPtWxDEEr1j9x8pIwjxv/ZyrylHXfox9/Nf4iseX
a+lpiD3fu1EvYy1+0Ihlh0KyPdVwqxn1cL5kPqSS8WxWtgJ2jFKBRcTBsaO22J7tJvqvWCabHQgj
Xr8UXB1NIGc32Dh0lMN/yARLddeIpt9dexNGGDKX7vjU92d9EirFH8edSq5K6URNSyJCpsvY1HJH
S0MuKdGnHnVEn2prHqV32uJADYrNlG/u7//cyYyCcyC2QfVVEA0sl4y+Lm81n+EDCoidudvPkoR/
6LeceFVe9BZVMCmlnhON7fSZMenPsRIY2VJkMXgTXHIG/KenCn9Yfpg1yWpCi0myMNiDfslU/9Ps
2OtJ0qEtO4K1A/GRN6QPT7zsds2Jf+RHR6iWrtbCJ40GKTMuTRN+gtxLJMODpd7/RkS43B1hCBNx
wm3AZlq1aNiJnIz4mq+wJDEEwowIscBF5XznDctbJBkFTbumQTXkN2f+xRG9J3eG5yx/zXwWYNKi
f/l2r+g1rLnyRq9/MJB0vHTYUF3Qxb22T0pE07NxCfK1us2xWTWBt11VqJ9lb4YOWEAtzz/0K+qF
4P+sqUaDMh3s+lq2lar46/ZjOXZ28c7AXrQp1n/RY+C4Fw1BbCr+8e6OhSadyGGZE42hypsMrF4a
TrdYU46xoHs42q008ayNsO+0wPBXIY8RWAUsCCxztqHTcc2am8fQFzeEhLldNcI6qjVoyzEEN6lC
IueC4M+0YEOA0SkNDFjNCdSgLDHKPAOs1Rt+5UnjRPscH4u59zf931MOCDADm2iqPZVm5IRPuGpW
FjlDbXRk0UpcTiYcG7EDToxozk0u/EDa6e1rErZeRH3NoD+1pt1vhkbKWt5uowYRJblutVa97TVA
bsBhTlS9hnSIlQbhk6BD+g8Z0SbET6/RhvEhGon+VekAB7yYjE9rxu/VTjpvouC94tbSTla4LQIS
GlM9wIDAkvtBloXO75I68so5InBIgTjKWTKzt/LfLLrcjUNF+OEVpX2Q2gw50x3nmiNsOVKCfs0d
P3vz7UDrK36UXQatl80/LEIH4RjTJeFYg7DCv54UlxasNonHYwDaynpPzpjlzm+PpAgYwoMLP+eU
RE6RL8sBXc11fCnv3+WblcD8Tlluz7Ffr1v5je9pniffo1WxLDiUu7WDZAJimu0f09UvFY8cdM4f
26+ma/DcazuLcfMG0YJ+rNWNx2iLwdLC2IzPMr7UNanwfhJpcPLjwrouAXX1QM7RpyqAYBl7NqnH
1/lPtnJDIVdPOsylOGBGL+U3ZB4TN5e+PGE4f7Wfu5vlRdjjX5ECHxdioA80BFd1Dcl+8ZTZ1gkT
8ngn+786o9Q9HdH03J6DGk8SFd0P/9gOwAX017R+/fgpt8a70EV8yR5UDXi7N1KEe81rSSxDAFXI
TKnmMXtelB2gTm9jEmujc+3pLaXsr1kgorZ74IaBEt9Zap2m5J+FxesphQmw0jbehTLtfu8l1Qxc
JnEPyCgdblLbcZCPWUPsyB33bFQp3W650fgbdUQAz8dIwuvDiEQkY5U0yikwTwR+miCXyC29hT/y
L9s707V+Lco8FOD54V4LTyJzHT6ZoPSdWfNazOHQu14/DR9UMnyskqy6jiHZW8LanU6kdVD7O49e
xNjclhi7vgs5Gdcj51YB8kfcXy+a2M4EmjbiXfGuithyCJC1NwrenGBMTJVojZtr55lumYp2vcXl
VDV7HM728MrWo9o/TU0/+HiIuoDkqAq+1TxBg34e38h2wwyumh2OzWcHqsVqDVgvNl3/6PGneEN7
qkp+xOxgjzJQsGIU+DeakcQdmEDKD0fpbLCeTpmV8BPsZ7r//98/OZQTMOSqCTqaU/+MwlW0qfq9
9hf+leu989iA8Mq2ntypyuionI3QhYrDlmjJiZTNNLUvdrsscu1byF6P11mnrv9Bka795EMPGS0N
xcquGQ/zu50V4lBNTBxGkaOcVfwdpOFrhqCFb23f05LCNo/fKFDz+D/dLqBeuAyd48Qb3VxEIcEJ
5uuFyhZYo12VE/bOSQ/87nURpLzGHSZ+K1FpbIkG6EdtfISDkjtljn9C64zaWURVESDWypne2ijL
s5eOUnKATgJzLUExgLdBo5GNHOu7p7Ao5eMDBT7UYtYg4CNWVnH7oj7zIlBDOJyN1jJyaSBoHnxT
4TSASvJrDCFYrX3bPLUChvdgmjKqZe/ErntR1jwtm8g3M55tJJ38as60WUfqAfsG8Jwy40+lnNmq
mcwp2neiyVgQhctxyLqQ2TkGcucAxl0u+uEffeLMR05eTc6G+0HhnYNHCvMfc/g+GXZ4blLKE1Mb
/V2bYG/e5pY0wa59D06ztPdavLBNaG1VAo+yVMbR+tcEy5UpXHHtzh0RaoMV+gvL4HiU5/PYUlQK
4y3ISQtKw+95tfSONOVcVjx08v8Vy8LQQ25z47AcHPFyxaMuMkADURfdgXVXSjQjf+mWQF5cQybd
Kpc6/Mssu8sDGle8hMlJpQFhNjrlW8TkhEBSgoHNN+J42wm0zcOI1Se5Pvkgsgnnjfy0k5929Yek
p+QL6Ye71+DHqhfSwiK2v7B9WfDpvkD8PnmipZvM2j5QxW+rJt71XXjTc1G5swbMQUzDrmTsJ8t2
c7dXHSP0reN+qgNPecDivUAB7qbZ7b0jMPjzNcRSnxrYA2vW4NO9jxAoV00gQlU+frUumKfFU9nx
B3YTHMuH1ZZYksD8sQP5+HLc+30tR5V55aLpBEtoBwzkF6TOsc3+f6tdbfbA4jdCrWzfu5ZEOJtU
FS8E8j/1EaFroaRmz5A5mYjBtXh6kJO24wJqOiai++E1Jo1YvvsSt8eaPpquXu6YmYI0Dncl9P+O
YeF2XN6RiBqUNW5ywdojDfewCzZhJVMJMYbsRfe8R16XN1EqnRd1C/1z89gtZ9687qiazO91SRVf
g++yHMSLp/QJii06rLwkU3OT6hxhI+85hG4AalygodlpiviIrAegwQUWO0c+uKb8TafJVwjPsSPA
fRnXj0eTpTaGtRQCS+p6DEKROMVb6Zq9s567mIEF42hgGJFuaAimrR1oqywzu0lQD3g7xyPxqoM3
f17+AADeacq0ckVm1yyhTied7tXnHtXuxTiV0tiGC3H3ihMplqLjrsSV3RKA0O6G7grjgdMZ40Sz
/iCfHiPbs9NQavzHthx6YK6NoafcgKN4tl6ZItf3wSi3CHc4xUMdtP+5RWpF4pILqung9RZ/KfK5
JocjlHxx9m24aJHWF7HLKZSNL7rL0s7KUDNhyKSTTCz8VSWQOAIkztszR+D5Por6oNvFsSaEk5JB
/AwTR2/X3BX5vNNxd1+1BeE+fjFPYViJuquQAeRVLK10lLYjouXiLbMFqjrts1674tZywXJd4VQ6
sJSp1SZVnmqdQdTpFxmDYIU9k5hTR4gMtrs7cd2pWsRvD65606SYt4lBSn/54nqKZ305+Lnwgiq9
zEHPtWUvMVk50kFk/RQAt0zNGELl06vD5VGGrpRsGd2ofi+GQeHbNfSJiLT7OraAA16obmu6o4GZ
rDUufAONjWchqUl5NhrWvtHRIU/x0m/CJDz41g3qB+KDpYjEFyNtIGacmpEVbyLL/L97mdoPf1BJ
laDUwPgGpz6VPVLrZcCZCW2xY9qcwAom1dOX2ybxXvkroCfvlVGbXBw3ugOLfHrgrKPMp+UtlV16
kLJ0Nes1blx41xD39enKL9xoG4CrLwGZ0sCdaUblpOn87TfT/zl1NW0mcA0VQ3E3gy73vCwnW5EV
qRwgJRVIs/VNYgTDPfOiIHg7e5VkxdcgbiJ/5Xz5FiXeWcTJN60PwAKFmgVzJPtsQZKPaG9llTaT
hUR1+GwhXqgy+12eraxO4MzPzBBZRdiGGjQWyUH4sWYgpx47rZmbHSXJQf1M3hFl7LT9KZMW0Ap8
m09+77ZR4oEPbv0/y6RsrFWVEXScXvaEswsLnr95RDO2+ydZaWhbnKqlZJNkiGdfaYBSHw0Kz4aQ
LwZNaQCy14nZBEe4KyYf55B2e10uMZWYuaJLlMTqL6poNb54X0W9yW/2k8b8p5MJAItlhTj8vIKL
CZbSDMSHJ3FSTjOtw6hRmEruzV9PrT4fyKewfYtyXxHAh8QdmI93dvRPlLyVhW4YAGu6U2SbrSd0
3/1YCpbcN1vo/1/tmg5W6Rzff3YI1I4XtCD5hFZYyFBE2hVBpB1mU1px5YiHH4c/FQakip7uQ2Xz
h9jM1YT8K1zmz3h2mDROky3DetKsUJZ9uSr89/vn0e5/kNXqZrUDQaIH++00QnPCMRAeMEubVE3Z
Xhd4NH5+jLjZvGWW40BfHtdS5ayrsMBBBVgSRbw8MjqE7hKcVO8lJd12hqjnIbsLtc3PtwvNtnEt
7Dsdr0Yg3fs+Kp3n4ae3vhNa0IedD3ZV0FJUy0yTgJ88d5nnzLcQr9WzNBGrIzu46P0k3414GoY5
wFdGn2JUXmSj8g6YpTNIj7M4fwP9A9Zu5BIIL03x3x53qOQrCJ+LkWiOd+xfdIhIcmzDu1alC+AM
YymtqR0WUZd80UiHmfTvSBL0hCctjJt8/fjlXSV/RJAFTcA4MotoSb05zIVQUFX0M8+a7g/YcxmQ
3m/k66pp15+tIlCeJ1UEDpnod0fkeV7YV/GSAb7oxKfKDhjAQ+9w2Qe6SaouMx+IXqG1NnYeE7CA
ZgQDSGH9PkXcDCQIsAdGKJa+FEHvl/W7n08BrrVnwG6gg7SfKfSPWb8lrk03fK7NA4x+bCGdYOLL
QxuB5OmzlxO8GnAcyYoO/yH8C0eNchD8/bJJNyE12Y2PTXl9ALLn/1vexs+Nf/AAGljE7dtft57B
2MqHlKhieLA6Xh+6wxN7Wgo4QfFMKnZETo5IozYD0wzg3MUdZ6jaweXQ02AwyRnI0MU+13FLQofh
zEc22+yMNXByy+o7OFj7vMSVWjKc6mtY44PSqbPIIzNB9wnaNPVakHD5x9/tKRajGKkNqSTntH34
bx7Vs6PlEr54ogM4ihahl5/WyxnPGjpqLjjMOxWj5vh21sovBqB4gVFZTHbmC318ZWw6t5HAE5qV
uzr0xAA7RyPB0mUr0aWzNG0PkoY+UhNSxiGVydGBFk5WS2sORpzxtMd3MSaPq74Z18n6g03660gv
hHiHFsBYBNFa7nypXo4dmk0DaWzkGNYfkbUH7QnYrTIbk0ucYKpvqN35MnzO/Pk3bHqNVZre5UH6
nggT+P8lRfsBr9+LRS1UR45Ewq/tzFWODtX+rIzIRyFN4/GRO9DKDtFKnJRIpGoN5g4CrisKggQ3
//4tF66s616dvEcxDx1U5JQvnN7njNUKav/9FxS0cO50nrhCWaiCTidowneSq9pdOJp5EmhKPOPP
p5gscwWNB5iBDqW4qUOxYYwBRC2G0CYkZZSEzp5/WaEZ99vfC8rdjcFUcNFBy35LvuKlmxUJYF0u
gy2vdhS3eQ1ZU2u9asHAqwR9NhrjyQzLolXC7BXYN2nmRjc6+w+YOdzYU1xTarLweL6Lf+TeBOjq
ccgpnwvTrB/g6nWpczM+E9L4qQPnl+ZX6HunWyFh4dZAvGSpuaCOEFT29kLqjD5QoX20YM3JfKwr
aMCMJtCsSLPY4Vx1WtwDQy/lYSCoQabgekzBp1sxC7+WrrcGmc8A3b8pZvpL58lkRKEykEnLaclJ
scP8NM3lzURiE1xOXRyYFhF5bAfK8R0cu9owYCokCJ1VtKggqBpoO6iqhhrXcO/5lrU/T0bIXzlZ
OrDHST6i+TIRIP9aE0zgWL/v4zvkkkdV8Le5SCORfqVnFlRpo8xnI7LMmDWsVqc9F+Hy/BshKnx2
ZTSJpwIJF/yxWNzdB1uf80E7pbr6g3r1LnnO2mhIuPARIKclU9BOMqePz8WvfLw4sjy+xfWnMceP
szuyyGxcMaxBqzklyLIQMmN1ziwLefB9y0zL4Fr8Fr31zjQPcI+qgc4FXH7qfg7yz0tnkhAzFIf6
4qoXaUvt5KBVl9/+f5b+eQyqzz5ffllPuMT6dOU3VW/ZYAFmxVLPy79dwrz/bN06kJMtX3M+aBDZ
g7hV93MW68sweBv4iadnZnxc3EZrZSRFOQQOZH332b8o0QuOrMMmJtDEfTTJjJQmtgxUEnpHqU/I
KrCAj8fsRNryrn+CeRkhtN00s4CynA36C0tMBuXd756ZHZGJgTr8UmlckneGRBEKr5aAncKS+RHn
H6pCPdDHt9sedZ3CWqd9zFrs7IkJlD21RxRdm36amAdqbzxkUxzLkfIuZYQdkvirasSgf9v5I0oY
hZj0CaVYLbQyZ0OomcItpFkY9F9Z1M7Jy7UQ8Q2KoH/zvdPcetkBdm+dMuHHfx/hjYi+PIxdbcyb
yOE9Yynwz9UccNT4OCQeewYIDOlHa+aG91jT1u85D1aPxZgFl46WATCBmfFm8hf0qNiKR0wcxbQM
dOICrdtEmVMalJz46t6VfwyBD6nyr0BClvaHtrqqEf7Lk3E+Z2w6Ewt9mBH6OjKtJY/LyS3OAwGx
Y1jLrC4/np3lPLdjGDGfsHIr65N8yTgKK65EtInR02tXkuv1TejjVxlfVj3FT0mivZ8FXkptWgde
z9i/Ff4+3XW8GpIYfm4dIRzcnSIFWXKfeTYIBTASHQ0XtbS0w71O7KN9GnL/456kPoM+MX3Gi+td
Hdf6HSFGv9ICvFqUETKxnTy1I0jZY8MbdxaPLREKJdkTT5mw+VtWkso54nZzWQLoMkJcxcPKwUrd
YAu1HsebwYM7I1ZL/Fi/vRyoC1bf++zN9Un1WH+F57DaE91lKppQghzMsNCzSh2XcbQ+M5sOd6Zd
zSUKfTTvoPkj3yfRHxJbOKS53KKj2moJebYgMXCPjNxJeCiymc2rJhHxidnX6FpnAm43C9NSy/5A
1oyv+HKN9YkFGqZpkhgRiWW2pnbE6IFyJB0zVkz4Ibo2wZJsQExw45H5S/xn1naagNpT+61xmD/m
vUK0bAgS69Vyd3ewcG7clK67aEiH0B6MGQJSr3QqZtpZsW7zpM2kunZ64nChXiHnSmWJSQMEIVW2
ArY2naQetU3b27w340WK4DSQvdfo1Wp5mixQON593wO5bwHum1QDl2B1QOpxbXNM1L0xNAgpaYko
mL45Ya3Eu6L3+yBLuGRazzEWtywegVyt+qJ2jwLCOH/BOoQwGxjbaJvGsr/5M8DDtuV9Rv2l5fc2
98sWJuohsz9HXsBC0hdI15xRE6WagUp7bW78O2OLPlbJz3Wgs8SknK+dR8RI/oujyc+sX9FZ109l
nvQ/4VcLxTCH7GJQJHaQrqQXfRPFnvbJ9qBjmvco2kYsKnyWeiOMk2b3M27tt8w3HAT2N+DD7YNC
hiQOYZ1KFHpS9+/otheWRpm6+NHusWYQ6re3pc0DMrnDecA/AEEHL95mFfytYQMFfa77OYWZ7Zlv
vkg0YrtUIUxZJns3GNmdpX8WCc+YTXF4bADqIq5v5gYvNN/Se1B6odBHOA/A5qQfndo2DhlKo+pN
hjqDP3lJbDjne3ADRxunGAZbKSAFG721rqDSCrP2XeQ1cO8W7MaTp/qj6YGu7yN2YEszy9KBrt4T
ysw9+aDor8ETypL5e8SPybBkSP+mVtQihPm3FGFwWfIB17/EpeYGBsTVz98TgBhJZZp4cD9ybCfW
H2WW9HE6CpOFVWE3TAJnj23ENjk4MekGU1sdOu8K2weXr4VkAQaDxCIFQnN9QLFAqgk/T4ME4Ro6
AwuRGRxVBjFEv1sfoqXfG1q7B6GGcZm46Vkv5HqDTfftxDehJrlr4chDoF8+goozxlHZGvQABffq
SRnnPqGsAc8Ynb1sruUCreI9qS+VXxmFHOSu5KmrGt3fIaxLQNP7DJK8UrFHcBZKrqlPa2LrymMh
YsLRVGOoqiBrGelZo1c2g/SDCOtyflVib0IRXj4w8VwS8fR18Ur5b+Rv6u4+8pDbtEuP/HTNlDMM
a3L9Ii+DuInipQrImjBLeJ0S4jv1da4fqwJBLEeyTmOSmf7XrJoap7mIwk+cxvrehna3FiHATpiG
FDKwchL6yf8Z4c68PL6jcLneknLB3aUP8zJDBEUNJwc0CI0o/79dAycY0hbbmaxMpR4SYQmvg0RQ
5NmWIs7XiWApSvOpUbM6dyU7OUNBXj5tu2zWeDO7aWsqkxQPX5q8Y2hEtsV3FcCzvpamIPSAG+PV
0iDKA2x0mHziILAULr7A8me7iIUAyU4mv8Rpcwt3yzWMui3fqnNW4QNV8e4FiY8vdQg0sCWBOXQo
SSjA7XvsN1HGcO/xLET2CaBmZuj4GrIGkwqSWeIa0s8EGNO4X5Ck4ctUT5qhule8kh7mO50Z8RGR
YvGjdZnL16zgLZlI1rarcITOHsJfeYZcrcURgJTcxuWwdgphST+JoxUB+nrAD9ROY6vkWRCyJopL
nHzj4/KV+VowumRXcgmNbOY6sloruofEM8T9iYP7skMylaUZGZRcnu5KTqjX0fTB9T6f96/ZZckd
FTBh88qB6fUTsAgm9TM6DDDmdWBOcPUWDfgJNCTrIZaW7NEujk9rmj4D/G+IwF68EFHsbEolF+kM
49Zt9T2pZnBvMOLJqOwBhwTOHaEWyXaTiGAatRtOH8y86t8Dr3F0RKkV+IlolZlhV+cXNc6q+K2/
92XAtWlQOu2xQk23Bwl3ElhcglMLhClKoZVGZeGUBC4UX2C8I8MerWihXxXxHtUsHQezBJ/zdJ9I
B+Nc3AiB0V8Np2fiXSwbMlMACMmAC8fI2EC3HisfJyW5/+nk9l9yvWyqW9Eklr0UiZK25gWjZRv4
4GOvllS1lbTvTO0u9isSjnvZmoI6Ewz+NPSD1e/lG8XmRHz8HkoVOkuPoRP3/3/HEI3I+wJudnug
N0ECUU5nCYXmwuU+GhM2ZZdUiYiN9LySXbe7BMwqq2AxNpDFwSgyZoYntcqe6NeC0GDNeoX71TqW
HPDQAIBkobrhvnOsETNLHM7ZtSr+EGt7DKvY3SE7es7/gxqxHhmTYV0pSBw6bko5myyBW1xy1xog
fF9W877uTPg351fc2T1pXs/yzRfxUe6q7DOsAbzjW3EjWvDZvrFvMlLUcmlaXt5bPUxpPfjsaVfj
1Z2CEQL7sijwXJPKi6jzV/I8k+oFMC+uJ/eSvuvShiATxKu+CPyP0vGFQJOGBgQER99fJplH9o74
UtoG9yi386vXr7mDfZRALq3M/ERLk3zgyYqUNaZOSL0T9O/SP+431HAc5Vb5DFJNoSnDS4Y8xstK
uABOSCKRlWtNIONO7L/uhHd3DwshH2lfO2kd5ilukzDDgrGBrOockCAcRC34ZHVlTqxsC4p5DCun
dw/f8sHWXHSd8AxTHgSQ+14pJaDpt/GuKH1+wfIksGKK+Hx4vtuhhp1QbEv7cIfNwJ1LBa78MhE9
jgjQZOcw3lTmZ1mBqww3ZALlD1CgSAMhMk2fCRBiDybWDIGDdtIpg7ktZ7lx0L4hHCBML+Ob0Dr1
LkiQqQ52GX3BzuXPsXoF2KZrzvoWihsNz6RlV+qdL/619d6es+HrFnEmH3GhE8xITIzrBrLKEjKE
kGpX8cIkWNV+cnP7CGIHW/Tp7QsH22kUNqHBNX3wiWVyNZMGljLVDxLYDY7mGto//N+S1Z4qcb21
9BP1mmMsVuA9X1xhtkxLyuCtD+UJOTP/TBa7El/w3itX9VhCRvqYswFD/bZb9OiSVVND0E+o7Js5
CpgvWfQqkNOrYD8N25Wrfa2OKhoIKWRLLotxyNgfHuj+SaXeohCLV+WxIotFuxsny7JX4EpGo5cC
MvkTJVOwWHTjPpmgFxWrWXvpr4WQeegE7JZAqLZSPo4HyZAhxtIyhjId6TUmzhHg1t0B4CSNOb5Z
BBYhMOb1uF0B8xB3949gVPwFyJ+Eni8nNT4UJXMDQDZp537YsZIF4awh1Pnf7g8TVyxeR95WtP8u
eBuvfQtlDWsvMYN2WECkUixflwPasDBYhaS4qi2Y2Djyirk8Y6XnfdrgxbrxS1v0vwXJhmZRQnlX
vLFIfsF4/0+PGYSjNy5J0HFe42/RwKusgvIu0qMAynmXfb+4Yc16JWq7Ta5TFQu5h1Nq+EQMRAo7
0/d/RspW7kggBisp5YkZ6qZiaKhEfc0i3zTWCLDY27S/7f6ZGDejGIBNlETts66RAcJnXdLvPFYX
CltJQH/rULs8FvvhKHzS7tQm8CP5K8WX4sYqxgsG+Z+P6fWtzo414Q6VLLuefQCrLURa0psoBN/u
gBsvdTeKGeDu8sCqjGA1LR/b631k/0BLR9iH9MPnl1k84JIt+inPzgPQRPM221FARwM3qOKLNh42
QDmvEPFw24dqKhyjrRvfLJay/ie4WkKUPvcx03Byv/1O8mRQ05rC2kASsVewLarg7IrK/ERDrC1b
EdUWOv/xm88eEszb8DnpYDSqNZJshs1pFcLdyZKDs6OpiJRx0yJn7nc840+MADrR2VbE8hZWieX6
LdTDezhd55FIX9xqj2j7EOHWXrSK4xZ6KYpVaTryUgiGvPWOD1lNcQGhWpZltw81Pm3Goi/Xw/Zl
x9kFCnhi7AsAbjJBe2US01xakb1CCIKV2ZONDEWnZKR5wgrzWuIazNydIR2/CxCp2KE2MYG3BOoF
yL3xLXK9hUCt8fUMn6Fa1Iftv7a7AR4B/i+yFDpf88xg80bATpD7UePIwhDm60T9C3NOgVZaKicE
0lJvKO+xcC6aMIzE5pJbK5mzvdX6+jOMIrJvRsXzByMAYRcr/3o3ToOhQmPEQJiAVE+emZ0a6phy
GMSnuXXdULqzhNhEW8XGUxnNJW37/Ujy6kXSJcRH5AypdMdrjSZebBQFVoj2LpndKLNzjYVnLvKX
WL1NgXbxr1VNNBNxf6Ohey6N1di+h1S0hkOX5EKXO1J979ZfgsWRQsfKLfcOGW2/G3aAy1VBslaX
PMB522oylir4c31B1g9X400AeXlfIsbwl3f74UShNzP0AafR9S3aFTAkrEPpx6E2LrKx0/kxPEgI
i5Sz8DQCGsJNHJdf/aBNAb4TZhM8Crd+r020GK622NrQe6IQTs/oBLQ+m/a4cddFgjUEyI9HINJG
vCiYZbxdoZVtWp05MKQ40CENd8CVl5uyEUj1lt0rXNbkIaFdZ0MOR3Zxlhu1iDH9EN6VLoKj25WL
xulAgXIEsrY38tjC+rP+rv8v0x3nZIaYdS4zOfNMisQDQSRs3AxkusbxYGk+kFgTLRIzNeSGL54W
zlQLnQFDM2SDfOlRNZD8+p4NSEPPHbbYwHZdBOaUuavMSMsvN2giPOgY0AC1ZkZV0GGExnQnSHTI
wxOmoVg32+8xivnd/HJQdPehWo8IO4/GteWexXhf3sVBqbST26XGpXwianCJEKjEeRE1hK8qq46x
6kYCYizHA0SF1GSe9wRWSFI8ehYmBPNekdG/199VwQSc2+FgbsqG1azDBx5pdktVagUpJUZI1f7D
LrvY5LVz73WhX1kCdKJUJixIP8+VyKTW17MPHyWKz0nKEtZRFLwGcN6QZfVPBQVj+zry88K5Bcg/
RSl7e/Q0n+F8Oyoiisoakt1nUvccHSxo48tcN47silPcdL1/ey5SA1gwn3zI+HMNWn1UjzzPg9eY
JLIB8lnZ+e6h8mLmyk9ikp1O1MrUtkQr92q4hn8kIcudaDlvdjDDiNJncPG/BohuUzgC7RTXJQkW
05IUWQsuw+3e1Ob8a4N7qAE1qKl8Zc5Um8UAAsBf1Z8ekwpKZY7yRCyo4J/VlXLffPh7gySRsjMr
GtkxGmcZomUUlxpvVTNCEUj8inqAJMcR3VOuIhqVmYO/lIrv4ChwIF6rqLrjl7qgQmGYTL0TyP6M
SdcJBEQkAw3cl60bav2VqG0NGtP8Isx6stksg2PIaClz/omuvTV2LqUEg6bLp8NbCix+7vradmGa
EBKNT3nKG/9tRdWWeAxAGzekLenMU7qO/BibaQD8HM5Vj0ikAx4jKmT9HQ5Yt198KQ/ywojiylpD
mUNSo8rzXORpgKdNGLlgxWzgqUX2hji2cRWaVaetdT67iNBEgGWTV8flSulODfup/W8RRdUcBjao
5wBT6t4LOouNdQKHanwv2F3AOeXE6sKISxEzhCKO++gZOwPKEHVgkmsaCYwEeWdfIQ1RG3EpkOhz
+oxdu4Qf4tvLZS6Eqkg3wsiddXewiYxPzKFDm7WJqD1LmY4Dc5iwZDkK/HJXT4a+cHO86K4rdcpG
bd7JR6Gw2geLq19jrEqI42u/XRiJX4cHNTmOglJ2mP355HdcD8cyYTtjNY9LcoH1R+GVr0FcvTgJ
IGKrs7SN5VOlxxzz0HWHV/E6D9jrE3ZThIvMKgR3MfUB3UJRPCg+arvjXoKofSebMWDrtqOjYDt8
nKdcWORTJ5/kSC9L/auxhxkodD4Wor3g5xCTLBh6EgMMWj1KQatfG4qNTIzWId5TQEnXuxeXGE+G
mi/UvVDomtfttG2O91he/RhNLsPBX407tMSLTWYHXQfMR+t5NnMUqBGFYXyZtE16kzotQ9+B3VTs
B6b1pe4ZYmT3CRUzxMIKRBIChVNlhzl1RVSu2hAl7KJeEQuNuLPmPr1tJ7dcNqTHlK291vER1yFS
dCGC/hJOZXxXt5GRvg3NNvclpx2ibMmeOPHNYlE1pIayn8qKGWfjCSbwcTv6nZc33ZoOMDU/Etjy
oNN+0ame2P836WrCjDpL+dkWGE8BT7u4nKIppHccPMV4gv9TfZAzhLYzpFc7GFSJEH/lkpC9RAY1
hurMBBoTwJ+A6cKualDAqXX/lm5YHedw1WMYBhWy9gsu9xeHXcMlO9HfaRzRjXt0x3lmyCUT/8bt
nMETQbSipkpTzkr93FmaInO+QMEvCHEgzIjH/4c3WUQfTL8C98Yb9Vys/GFgmtnmrZue90d8+/DQ
a27EwDE82PI+PGoGfDbRyMS5L7CwMa5FOOi3xZYGbPg2MDfGLMD7Xe6HSJPMSaV3OVCln8tO3fpi
PjKksYHMJrddf/sPVP9mLORRrigG+PVbl5CoaPwOLi/XqwYnognR4cfjyrQwUaUpH7sk1kGIVpqL
/+Wh2RFaxxVCVqoiNKVA9jQo2Do7Bjg2kV2Hqp5530NUVctX78KmtQbW8FSC54rAuWbsytNb7H1i
n3ApKqX1X05dHfhsBVAij/DcQE83C5QqhyZFJ6/Z7AuVxAKwHPahHqburcH7W84UB1nHfHnM6MpT
O2W7f/WP5x6mCIgFumzXoqvpKaCoDZxB/iy0WaxGj6eahzDjubEVrliwxOgnP3s7SZPxj5k0j8mE
hph3Jc+UPBS6/JwhiJu+bYcK6gQE4FosYNkJyJ0bx8ZJgU5muS1V//0hGqty/4F7N+5jGREQzHHs
lRSJCw7WYHnwQKqhoqZgjUjXdZQ0ogNX0/EXjZSmhOM0wZyOf46I8zR8tSl/mc1znq/jk6FeFph9
R5x1gzo2hjyTlNVsuVtQpBgG5rGKUFGIMcBXbzuOZQQRxQNa/0xke+qwy5/uZQ+K3wFrw2kLFtLf
WDULI2lotq2JBhetW/joVW5IxWytWq+iRGgInBwhCpAByRoOKyuJR0KF7ePPGj7KLJm8TEfWQDoj
Wxc0nU7rftmJehPaa2sU8e66A/Q23KvwxNLGRHubbc2UuxT6/y/OMfh5yPVCyyxc7DVs90RIuxqh
R4Op0B1g6T4HTzNjyE5Lb24+6sJEU6Rzax/q71yRCeU370QAo9n3U7IzPcJ+hQO6wR6i0N2tVNg6
CkOkNdoMp+Bz+YiQ23vODwMSuOPSIVelIi5386E9b0sPNcrqQrWYM/7J7WetmJQhp5mE1FFXWljt
c9fIPkIC3g6hCMEtVvmK4kekHfZkkVoy+TIh+M/t1w/SQhB5VpNi/N/8NHW5j3lIwY97gntgUsKi
74YKI0FYBBI4cvgaCtrD5aD2M+m0y+7B3vKsR0lNAwspOsHoUM5nv+BQ6QmTo0EAaA423UsD2rcI
AGbCnkRQdRKWVKYzqXgfltWpdXi76I0yD7lQ42H3YY+cfCMj6WbKL8C0MNAKeGyY3glgB6pzQJPr
b86FEShbWcVP4LHst5A0qWZEh5UxxpnxQM3D2fp3bOIetZU0pbbelTymD5ygnuL0eE2HgOF1iunP
KQRivz5p8cAWJFDLVa143v2zLqDV1vL0/DAZSMAHJwsSzFUiF1B28upSL+pxLBN/riQgbTeZt1Ar
3OdL3tjIcTNbIQweCRlosdo0dIAwzSYDThXUiNJgSZSTesgRd008g5KIRS2CfrP7QwGbqORcIuc1
isWphhwGzrJHwBrvo9MtKW1aFhikyv5YBnLz9i23KJU3dytrcJDvlYeII+ek2xJ9xZHLxOYqKP+K
R5iuG7tb3KVXsuj2jwSspSbmc3kO8O1AGT2QyZTY6KrarlHGk5/pK1UJg2Jxcg9wYD4rhuWkEFo/
9DMt+H/XQ4KvkrhmmCcS46vAMN3pd2dR0tBcdTjOKi/bPEvHY/6yJjSuiXW1PEXPv0VGEYyfY5bO
h6vgiPVWf7m8pAqmKW/qTsd19OH/TOoqzb9oep5AiUfgrofdLZEXNYMNvB/M6SXO77sX5GhOUvAd
Kotm9L5/dqQZ9KeZ7wenQujYS/FElXJ1MJek91yz9+QslTa5m2dF+f6vg0QCLny17NcFYZM6rpxI
XVjFmhaNWx3IdHZyqpC0A03Ij4cG4hhLleTQJEdRv7ay/mXz2ZT+2rudWAqNHo8YPvD2pYnP3UI8
7IWgFxLtITCLwUCajDt9cSpJ9kC4T5PSW9QU1/+EWUvDLNw/GzEFw5G3Mowcx1cmFApeePC9U62b
yqDWKmSAytZTVHPOJkCHnceR8vu8JmLebD19jUNQuMJVqXLGxkhsfs+0kLtXf05SU0H7Hps3VUu1
YtAvmlAg7vfr6h/jW8s0yIo+WHAP9lNjwMQmSX1lPPJIi6Cuzi5sFwY3U0q+efq2UENXZLTkP276
xJ5UUoGfWoshrGBl2stHrbdj7Bi3DKTEbg1I0W3x2DA18mkrgIB6JjqxIi0wdrF12J3lTIlCDuTs
MwJJTkonysC4GAWLswRqK/m6CFZS9I18ANm8Q+O6dZhwsg44h9FiP+RMH2fUnZ1606xcDY9UNNnr
FAgTq5CL3D33StHfSykpQdbPpnTVX5BoWwK6yLH1hn7aOYEgYwB8u/5rgk1jnVHom+d9gbiq2MZn
CuCkUBQCyhb2zk4M0vSDz9nRs7/UxGwYQ7bQTglSbA2Dzf8JjFz2iFOXmCglh6IOCABvnIZ055I5
vva/QDOxjV5dzchHGRjjXeAMpF0T2IbwQgkoK+ABa3ZeJK4lsD1tr95k14/iLhhsZf9F2G8ixSK7
B1PKbzE5uPy/zbHRSPP9zPadvvZpy86qnIVf123uy7TDq8VlPC7+9CdsenVHVOzI7eCaRP1gAXeN
GwPeeCxU1Q6brMshWlR6/fkorMPW5RgshK6LIwjhCy0Y4Z7gkxdeztjU1VZSAQdXAK86SOPBpeGv
tX6fiw0TykzKq0COLnpkj0ZDiZ1XEW2IZwevWzzXkJPXaGHV4da+oJRAQqYjuvbBCQGPFq6u2/Oj
E6kfKKtdPEewNgxfjwkRbed24Rv5m09NGqfGtXe+LX62ep14KvQA1m0gYcAj0LIptUBkB3e9OWAi
3c9MJKtVypS3L2oNcAX4ZW1WQJQxE2x/LCDZfvSQFh8NCkYa5u4y/lk9rtlZPBUtMKqGyusBTXp5
OevaA6JOPqe5KijqIqBQ5L34RuI98s9J9HzZJrI8aNm8feqgUyBbraNguMUIhkrPvYprYnx1yPrE
osHbNoRk5w9jqB7sJhUNgv4An7Dalv5aHR1i2i5Zl6yOozB76k+p9uFrLHzUhCCb1660nf2oI4W2
lmyFCCJ6C4SGhryMqi4trQcGEkylW878REplaC9zOGtpUB6puXV6Ybfbtl+m05Mzd1j5sVTkZ8+2
b1Dt42y1KhZQ3Z3lt2NEBkTFZTciXV8p+9hgq/CQ3Xq5YFSLdkN8KjA7gdKnQCNTxzttlWjl5h8i
RKI+gvH2XGX2Mrlpfeq1fnsP4GHUoxhgiTGHtKSpuE0i3Ue1E6VX27P32EKuLdt0JoNYw4gAoEgb
6XDgE0wcEG+6V6lq8+p/x3ErzEKj7XCUfnXlw0TrnxqI2y0djU+w9U0j3NdTrUOMpiRh0/HfP6xb
oNdpahHNE39WG5JJ2QOL31KSNIjCgblCxcoLNYonDIIUSwVwLBzpp6qerOlEv1PzFcnmN8iYoWnh
cePi2pxOSdTj1Pww9/BGRFgh5oifPXKU3t+l3ZLKKAqq2Wz2nMMOayqEHuhLtb/Sx/ztWYaSnVxi
wz0VM0CptLEN3udt+/P+vHwbCCgJMZN+2zugSZfo4rTEsoH0TAdQOdCN9mXqmjRWlIN5uxTh2xxq
onTPMQgcA9AX104luC6J5/8ZmaImTweKqFAHxAbtkMu8qZx0Z1STBTx3XbjRN5aysO7mieidUkly
n8Q8RANWmD9gFyIbx/X5UbCnagFqQ6hIztlw3YzUVkzowOYKG2j/nZFei7O8rFze54pT1qh7Pv+O
Q3u3noAqtZtdGh9z6PgW23jMXM0PnZTCSCBT9ym/jv/JKbkysArk5B7kTh3E+1masNP28e5/MlmA
SJPgnX8du4U161w+iq4r0B/tFcxbyN1RmD3ggcAy1RxNOn8DZSEJGMKj7xSNS53be/wIpJAn0bAE
NDj58YbGw/Z1nBN5HE9XYetr8uKDGigOk9dua4gCvgD6MY8wC9fIAlWC3djz9RLBC/kwFyOm1zAN
KwQZaKuPRcRT9vGtUy+pTZQc78TF26bVZeoCXW/CAQZG60c9KucCwPR9JrBamb6LHINNDRq/vYsL
1wTN1co8H0pt2R6MWiBMgy8KS30EQzBXZ4P6zmiMjub/s+0G2cIE1z+Xn6DtMpstzHOKNPwzHCop
VnwHhNBAk/bP+ZfdXOVW2ZHe19HOkaMkfJmADdpNrLgJNeUTpHvgfaQgQomB5pIMzhEwOvRedmXU
BRQNcJXeCWjsTKsP2DeKHyO46TOwdUK4xiNIO+sYglzccZPVPcPKXh2KMalX69pndW5SEOjZnaK7
QjK06Dy31Zdil91YyzRqRivcTjBkFRmDH4vHFmWs964tqmvkD/4eMzNLOMjB3qLwDFKaVCWsoPT9
lB5clPlma3+CeuOY0gXSMtKr/w2r8nqlWHSqXSOT5f1lg6Lp4oDrKPYOq0OXq7ZY3WQgY3LY/cvJ
rrGQsXA1VjGZHuXz3szHPK3qnAnC6UugFHf02uJnjmzMJp1fzutbe4lWqCdz/bjqK6BB8vUB2L56
2pfsJ4WqkVTs9t9guMVivrioxeKmd/skpW80pxnU8l4M+eztyNtPGju0R8FtGj77XBDRDG5yJyc0
0byglmoEp/rMjtBSBFbuU8fgpxDAHiTJKx2FOO6GQl+5Wy7xqbRyOjrHHdTphLbuDJJDVG6rwAI/
xf3RT1DxV86d2XdEaEtAwigRxiuSQ8zunqdCAfMyZA4L8z7E3p0HF3C6JHtBVKj3PYsV+gGH3WgV
k96E+hLtrCzNIk05lCZ0WGVhTOXjyKYboBJ+e0VyTR4f0yR1wSsbLEQ+LCRIURaHGOA7ApetpDfd
xOwdlDc2j9V6BZWtzW6sThVe09x7LzXL2TYLeo8S3bl5pv21ZtuXSYDiLThDZdbajho2+1WB+E81
2q5CDKjGJ89O4SIU6iJMZe29J5aKW5HgrNUFUpBySGdTjbJF2HEMECO9FzB2Gznck+E2BIc5Zp1q
zD0HfqlU8cNiDymgM8UMML6vY7zvc1gWwv5nI0LKLm3pMJvAB/RNSTHW/n0KzaqTRCEq2rTnqpsv
/IW41n8aWbZJfxdAxwtnMcJqltLMBVVhEbym4HeAwOvtGHkj+dcJyBYCwE/TOaYy+bZPz+eFkhjN
gP/RgteLbUSLpOoiSQDpyNlqGwf1FWNAHoXRyRj7Iax0uCtcbReynqPkkl1KDCj1rVbrZ43S+KIF
hEJl36fAFJm6V7nVE2K43Xl9SFDJsoInKVeUgO3n2/4AZCqhHHeIM8fHz8dDByQpYXMlFcrj5eh9
Gg/c6Y4o2n/rNPpzRF2Q3f8wbU3zpavVdw9u4Uy9UookvnDuEoA/lNOsfIQZTBUneONzIsq6MQaE
Ak8LJMW11CAiNbTkiwzda2HLuZv/4NXP249kmJJma2TPH2uSFWhQPLXJyhvQuwrMV3+BEqQ6wjv6
4EBLz80yVFItJZ1m609i6TWEj54WVmIsso/iYIS0NxNh7NdTn/nWGYcZtz8DWVEiKGpTLu4Fn992
xzYltsZdCQDsr7BfbkeQCCYoaobabxN+Qs792uYIwhHnVDCYB3tahCa4FOixXHN1ZKY/OnFYCE5V
j3v8pEh+mM8b7PTYI0yIFQOq9gAxWct/InOJ0Qqz7iodX1W8GVVI3sFTJudqBjifyvzhXe7kf+K7
iY3OhQWa54duIBtM3QM5bnEhSeq6ZemjnovzKSRuVfov62CoPOJ8g/82DfXKCaklBD+rI5dU6nY4
ZeZk32J4Nlh5rDR1aEQv0KM6NNo0CXFXHBQINNpKGbXeUVIurEu5otSA3Fhv5JugPh2Gsh6yhMl+
LHrACxwWSQ8XjXm8c2mHikKkyem9TVnFwBX5BApthhrs5JICHAtzLTZ4jx65f/fBCw6DVzVBfU9t
V3GIOHxghj7VLRIzJoxZzV/sc+H6ZeRQZg7WBELjH28TLF7ZJvQ9R1WBQlkmaWK3CQGXZ9mbdXGu
cqNfzNLBxz7b/7qZZs/xlbmRHZSyLDXW4W/5HdhzKmZUMfnZELqS3lYKb9TsuhTxxkj5SvpLcSYB
/P7+A47L8QG2cS+lbUekWSPjH045zC1Uj3npm5hcwp7+6/SsznDETljHk/e2E68WNTp9pzQ8p9Mp
Op3U1dMH5pdRpBpUOv12lc7qgVWLrPiiC1kFP+EFG9J8fdDPbKq2dRn7BSNw4b1YAgv0iYzfZ2Sc
2zbldWYWmfotfvCD6lKpniH7yuPPZ+Q123bhWz3oD9Er/K0wHO4z3idY/TeUDaYzDSS5HsFru2Au
YVM19U0ihUYw6VKrlLoUJzY4k0nmshd1liCmIMaBJYgEiWttnMu3ZfNtsPDP/3a9wFH1ua732gg0
qPu6XxOoH3E3l772+DGAs5t774cYFrKHSi0U2nSUrACvi05/0aiEEtisRrjtdb0QcRqVi3EHuerU
9eUAZ0PoMxEA5QRjlMIGZGCA7+jYgfxoYGm8HuTsE10RDex2IorRJyul7jKlEPzFCqbovAC2at4p
MbVI9J/QJslZ//JFuma5/pQ2NzgwpP5bpFxcsd7kzv6RJeW7DBfeiOyInXkK60M4lRcwz9Yi9EqU
so/v2e2rKxmsJ0TJRiDtppRGmAQA3CWoZ955tn9VzYFa9YULS3QyZ3q7lXQhm71fhA++xa96CINz
si11gU7UOSBqYkGbPTX7/ltsK9UTr6+ZcURI542T6rEIdjBedq+I82orq3boCkbJhPvXGr7rv0Sz
zAHaNjQk7orSEnXPFm35hBFsMYObA0+wTNSz+G3J48jNrlNqxJ8PJgsOCkByd9BK6PCbmJwBj2Yy
uDgSYkuaJjSc+VHkCUunJCeW1eC43W0+nxxfYQ0la7Nkn/VusczUY2Ph+UECpvU9UVZlp1bWMvuK
ETtxzJez6OupXWHPlH7Ypij7+eQ6AUbE8xwmSkYjUP8HAd5EyQV4gQiPHTZMyAl1HJueW6+2VEwv
OoFUARBEgrD74dGr3bFtX3uyeo0YWto7Q3UEQffSi20v6L9Ie/h/A7rT1rKQHe5cZzk+be71k4rB
WvkmFV71XO4pmdcxVF/tyZXouBWnWUcMrV9ZYQLiGx5VYYsUN7kbGBEMsCmJ2jkk1b12mLnDXV7K
S+neRileEWX3QaY4mdQZN4OzCRVU7X388j4mEiwn6cgoq66mercG3P6Squ1aP5iGybj6fqTwNzle
RBCYfkZ/0S5o+hVveSBZKUpilj3LkT0P+NGbSC+QZkD/V7Kkq/Mn9sByUm/Y9SAM5sEhst2doc9V
SHkrVHEFz0s1pbRDd0WX5TgNjINpLC1E9xUsfVufVfftudmQppSJl0AjmqWm3OSP4paC/DSQwKk5
xj+6gUnyrQM6YH0T+HLsVywpbunkPpwjv3bXjaOFyGw6PWjUoYZUN0+lV97nLJyWPysBkLFG2XKr
TZn9iiUKhqSRzymg3QosZ/dcxrEAsEqoRChNGuRLiPZRWfYmrSghZP3hsawxGKklhdyqw3jzMk2O
HBZFPLKdK2raSp6GqXUH4lx4t7UOg2S1J9HPUptOHXLhydTOC7UETIpRXYP9akfGGbD9VZrn52HR
cRRRkot1jyRlxY0InYqGmuJF5G8H0BsL+3l7iAzBjIY01Rtd01vGes4SwjcW4vO17TaznESmR6Jc
m5h1LmGZsOt6xPEShnxy5VbU9kKscQ1DwvnSLVzPCMU1WATI7chSM0oDVZkOaZtweAMBEgP7CxS3
/yosEywt2FbqD66sG40ZcXMqIYKfLT6ohANhQJD7pAHU6NqDaXshzqUikoSBH/QWKwPr3oGDla8Z
8ZRIX4PlJy6OAi2TwS6AgHsXvAFb9Pq5J0/lbm/YaJ+bQFBXWgVrtNg1m/M3w548pgm+0VL/eYnw
sQkDXcACAEPYvfXNA2FkiHiEcEOHY4x/H7CSWtXCI4N4nCrORnWO5GVXXvtnKxruKItaG+Go6xkR
M1RVBSjfjs9mWzjgc9+w2UrA2ryePgiuNLxc9nKcfSPiDDh4HDOkXJBXtvv0nhhptM0lwqGmDK/9
WIfMbG6RqoVtkeDBg4bIjB0v1SpOEC+T3IvtzjHbsw/us9yOHSnVSF++6do2dGnftqb3j3UEaKqd
b416CV2TT3slFExfNUOkFfxJsbXKjT2C4/f/6/5dZ5XaGbVjdOpgVSIAJI+uVwI61HB1eSy2GykC
cfut866z85Hq/VlGfW1EJN+2OoxgprTxotJslkvlVTBNXJsqH/Y2wSBs7eqb2F8+5emHWNMZqKMU
AilmrFMOCb90Dd7Ib6myza0RWpz3geFOvmG4BM0Qs7uEyyYwEkeHKgQZA8WLsR2ExtF+vsqP/yes
XLbQpmeRaun0ANdpgCtUKyfEu9V3l2x5zZeVcf8W58Im6Bah52t1lNS/6Ak5evcpZthwYd5hly0E
VWKkUVORjfC4adRHxdh19YI6N4lhQP2bd0ocLfyhlSUCegaLhVP3uTWB1K0XzRfIV4EhblNoRAQX
yDiPO/AB6f+B2XYmy4CRqcO42RQetklgG073bp76yxPaF2SOV4yyGuTV3+VWu+7VP+17qrLs0EaI
Yh0qlUYIGTw+jHrrijR/J11f301YWVQhIq47tiBQ/sxQJMZf01PvDUhPr1IfEdTUcLoiPdB9Q11p
3hJlVn3o7tpxDt3nhQioKKHBG7lihNuF5r0IIZtzGUcdoZjSDnud1rkX6GJ8k2+zc6twAJvfl9q6
utUZExFm/usa6Nc52GncXXTErlql9w9xBNULhNopUP8p5e3sRm6TWEbERDfW+z7QYz5/Zd8Xo0zM
5uYk7N8v9fl7yX7gkMJBDn50FaeBdBaSmqUdaMpnETSQHG6tZE/nYyPlkGGiwzURbFqfHpkatJom
6wW35lfmvtY1QryjM7zaUVmQ1cNRiUwfQRbrLGiuXiRtfKBVyxalQpPV8GL6pcFJPpT/P33j4oa4
cXgvGny0g2pemnuAR6tPJNXwZZBMKijjpLF3kpWYUDH+iuptgFhNm7Hovhb5Oe4pTbYnQBIF1FX+
6oHn15mRy8Q2w+T3TwffMf2j0O1DU98dCszZPiYUhS289u9oFq4pDSsEbH31vgYu+K4AKWrNbMkZ
bOZVJkO28/casg7ACSRd0J+oK/biCZbhNbyxbmTz4LLYTV+U+spGop4wJRsJatjWa92Wscfjxxn3
Z1BN52IVvb/oxxkh4GT6kceIWv4Bi3dFmbO33RyemZIRV/KDM2Fxq9qy50G/8ctN7YA1AweQig4x
wT4XHasf2v0vpW9q0VBFcymAfGDbX12XafkQVqD4dPjj9vUJGNnPDtJ2WE/AZhtflbLXEsv95w63
hGtL2YdR33JJgt6+dsbUKsQHX0qPrESj3qOoCtCliuyKVWedR03wswEmhFM/N9bhsGllnzaXYFHR
s670fMBc1jh1+YWNLCZDk9MWDPELzIFqwHNINfEDMQtDKRxBiBkDfwsAwsDu0ECvvs+ud8Af6tGC
3U8FNy6NsThz//ri+Dw/mcMFgM/rEZ6YyC8HeGgzRfr9+GmN0NDpipB2f4aTJH5N4rjmrenUumpe
vif/TxzBJ3yrLB4r4zq/tuqgeN2OvaZUemprxKT4FPQseIfCF43NU5CMYs5wuZk15lJVyDE41Exv
iXR90vQDWsANGYDFnhZIKBVprOc9DpsaYGPqlBmvSl3AL6cBqRbl8w2SOjs2eWR421Pl1JJL0Ei0
9zN7McxXpffUMlL7dDk7HDZ0iAzLPWqxuydA74+IQg2UhqrNBRh4PgxVxn0dn5+k44VmqVhh4VV1
Rcbndr2d9XJlDeS/HCus4+Y0C5xmkf/YOkrjewegfM9RDr1RiT6CU2+PUdfGrA1Fh3QVXRQF+7sW
LI7gNU+jksZVjEWQOJs93FUd1yxdm2bJVf5UqlO7PnyYLn7v4qK6T3aDzDDAsLs9F8yP3ke4UhvK
v8xU0dHNoAor0MwbLlDbVnjMR8u2sHcFbJZNgbVGkx2BuEHoX6rg0BJM4SRITbAuggsD+bq/vn64
vqWLQxdqlzTFrkaTXpaNqFGDoCPbVb/aJHms2PwZ1fzHslKmo2XuZNyNRneWTeWSrNVfFzWtfmOw
59AKeQySZya7a15BfnUgOhp6yUfRnzOnvPXBS+lg4sfIgFZrjc2HKQfdFKJUuh+3GSXODXaGkOLT
0jTKLPC0FCVHHpjjdgpOF0ayZT4dUc5bE7M9bJOsZ/MuvLeul/AJxkyCTTe64HNNmdSmcDgXj5Qu
28/4Ixs1K1pgplQ+mJuiYL2FVgNLEI4K9r/5GGrreccmdjMqCzZyjFo8vWRpohyk91MIqjkZ+sH1
/rDxBRkSIBA4VRy6cGabMVPrSq6fmTODvB7Hs33RD2qJoRLwRmfBlXKtKaaN7CBtYbLSVJjvj0zV
MQheKwWzFMxH9Li4Lv8lIyDxzsPxUd3veKztdDXIVuQ8fw5qwKqUmT/yl/6LeTrQ2+w/d/MLSI2v
xwuRn5eYroXTs/Y5TBH7TrJtd6l0y2bm9eZncCFC/im7jEiVA8sMaQvV5ygiZpA/hxDrvFfQvcZ1
4CHFJThhS67KLkl/lWkMmCEkf6/2epxC1T9vvgkV90cz11mwpuMtb8nhuRKF7Y1ycv9JuFy0BLpK
8RU6i50O2k40NBcUGgvbv3jii0sIclKQoSb94MMDQgQ90h+WFGyf9yljOO7o7EVtlXOBJ+YzT5MP
LH2NpB59meK/r1EHeh4t4EnBc9AjJnKUYNeHorgi0GSgR+v7FZGFC8itxzF62nerpcd7y5af8Fv+
7jU3WNTIRZFfBgu+TdvFYYWAjmi06nB3wSv2H/kWTD+kPoCEtgX9ZZI3SdYF/cjQeX1cBG+azVfJ
BIcRgZB6/rEVhAFgM4ojrNroR2NbUxShsvod1yKvwtLXpC5bSUitemWUJTfTai2FbmQcS6r4NhAC
vlURVJBdAUXm3Qocj3e0AcAd/+5YE1kBemW7+pgYvc9wYMpqsKebYGXGqLyokWTT3V9+WWGdXO6W
1IGHscavvd5YgB/bIfNpTspD9oBbHrgFAZl56IViYyhS9kBp71/OXR/sRLu3R6OAgADzjXiPqna8
K7YtZ0PiUzWoCUuziZ3qrLwtOpFnd1WvElKPaPhPCMOMHpjrS4NpSfJ5gEDoOCqib5yXKLkyX+wP
00l6d+mShoGrE0/RrpzOlEQvAI/7czasWdS5HQmDF2uU7FdE0Asg6iHl4bOkczfW01W/GzCfXSY5
HPk4sYwFBpHcSjmf1s+A/Mf7DX3mzD0ajKEsn1iBVWBF/tuokD6EtyaIBFO0AY4LbSNtvNFeVi05
o3iLpUFPWKbJSZxjcV3C251EPbgpPe9gofT8f8C8QJW5ChuQ4Utqtr1WwoiREBuOrg7RycRGe60q
mqsuwIW0ZQLS29CjUppKDtoNwcMaE5B1UZn9gA6L4/1JHSS7mKhvHes5LWrQ2vftJI4DMm/Qftgl
8SaTYPQJK5oEw2AjocyFhbL5J+BhXMUcUZ9SHqx0BmFcXZaVF36Fe99kj3vDJSJOdIv7R9qrzKe8
XR4KFVO1lPwPDnX3/zB1/LOoc5WBVqagpcormoZXx7sYKW/7aHcIXl+kBBKcvUyLAAuazJTyy9qP
kKYaBegk4WpGkvt+DnCCiwSvWhwWZWwuZHma6t75C2pJedPWhrqi9uDzGjV5TCXx6LHGC31V7jcV
7pjkegOcsDSir4fYv1nhJV/IVO2MOXb9rLYgpPVA74IOVwp2KjXXXtbpfZoVuDh19w3jUnt9K80L
GzkNM1yU6zRuCSGJAc2cTqH9a0XIZ1tgvUVIj23WF5FO1peZZwY6YzKr6bxa9lverUiJB3LvZnNz
ssAtXvQhFGmTqLo0NqGcXd6ug6Yewsg576eiG+t3R8B3KCOHzpBk77j44mCQSJAuASRL+u8Qb51d
5tk4R44EbBKBA+CbCBqKFl/xVWAVfCwhNkAiS3ehrEXeYPvnjoSOwCS4XjjAgGVHRSu+hPH586fj
uop6roaKv5LMoN3qzNRxnns72avKvaV6ev13SJzHEVxorRiL1Pf1KW+nDrLLaOcNhUXKotY7KyRb
vf2J/OMxHlksl1BqgX/vu4fqZzOtbM2ZuC1Bnpr3lUIa3fsuvCFItPfq9FP6JMbx4g+0LQ1v7V8q
j3UNkmocUonpyM/cFZOHdH6F6XZp6cCRIM4C5JerHdbgtqRoxvbM76nDSl1gA4oWElRkYL2qb3Ze
H4m6tMEi73Gvptigbn3VBPtA4/DpIsdY+hJKhmXzaE1MIuY30IDnox2nlyN4LATl5hbqZEbgDMXX
SNiwycNthFpi+BCbUjGmArbTa3KN9oQvCEY61B12WKjLu26cDb3CDf5BmQafgkZ7CykLe79eWaH6
Q3DUs5P8muh2VMTGgiFntn/UWUQUd16fckeUGFkZ95KafrmWQgsGQsC7GIgjP8KjWKT35IBAtMbB
NpobAWHRPZLMQe72S23o5cAlTr20uV9ya+4ntZ8oRgE0gqzzPPnG6eSwJYMg8kx0wKPPga3/nwi9
NU+apJBAFgUCfhxC4GYtRPw+AnaVXRGaJ1mNO1MIBPLsBV2fvID9IfKQKO/uKzCUBLfVzVsSKHU8
ze2KZo8PHxkELUKi4ANdEaGuuIn73BJoX8XFQfPPi+Di2JxQnW7J4ix1zfaKPVjSUpISHnIQtVKR
JbuH5xkaWabpJGYwUfepIjI09kY5Jn2SbCOwCfjuD+5bNJsOngdsFhpm2ehLJ1ia5co05WMySMq3
piBZDozizP4YRcwAqNj67J57Hp5nOHMOT3Xqs+3wd/fovvIcTIP1epuJgkqUa7/KQtuN/8//1sTI
ac85HWrHkENbh3wTBGatolAj7z143Sj9UrQ2lXUlX1aSANmefCpMg29I/HMdW5zAg0OfTptgzyi/
D/Ng1dsrOGsRKzXtFyjetozDYrCq02aa5/Y41CtQ7b6ABcV0oLfK38zyRGHuy28dVCyNAHbz5OW6
A9gBdaQA5ZvPhki174zQPJMsa16pJDMmVsPgvqAke8WvQKiut5bhL/AmQSRJnpOxPUnsff7ojFYG
e8CkGVFfZprsIKADk3JAITSthtfINAg0EeKRq7vuvGOf48gFLXDHe+PqGLYCXnzyals2unv6I8wC
160AUAn4uWDuIk0iAACh1v4JQTkZfchq/AED8GPIAAr10IOUWQ/J2uI0UkXVHo+zVva1wrRAjEpu
OMfo0P5khfeaDhAEHjz+/eILU4f5jzSSJCbLqS3k44gUtg7UTOA+3WQD7qzAYuLvrrx2hICvaoLD
qaNNFXIYssv2AReukiPw9Qu/HA45bQivYgFT+L+xra7HUCEEkHmbIOMLxVnBPlCzHpAGxH40bvnE
vRLpzbDB3Vrj/zNWi0DzpPt69Zatf01z3p9uMyEgBNzDV92xeB3MA4ggeWg9oAUiEZK+SslP81Cq
jPxMoKD2NXsuCu2mg/E3acN2p5hE5cj287Cv/izfBGbcfkYVh0eMH0aOcMf1Pnxk2Sk9yL+wru6D
Fd5qf5gOc1NPQeXlInj/Dm0C270sL+xrr5U0qCFF+fA/YlF22XmesGno/RzrSz62ZJCJjoyuiVdj
DlMOv/5ZmGiUYHgs0pW3nvV1NImU42HgdHOeq/D1xHAzxCI2X8JXBtLJEFD7sIuv+LJzFWPlnReP
mZkwVnVk7F9QaH9i6wjriShCgvKbRt1rK5phLCdpQLppKgyNfkNuOUnU9D/PzU1Ot1UmsFLhoyh7
Wy/spc3iE1vt9gelFovc4bNSlRGoggTOO+mFhB/YjeV/UwtuvxLm+9gCiELUB+RAO6zVTUx3yWkv
F+soGax61MDAa/kJotQrPGeTsAFdYLJ34fnb73Itw48Tooil39zRmqQENViI6JZ/c0jR7hVn6m0Q
Ct9XZaeAEiN8pRQLH+NefdraYZikL87Un1MDcQfb0/XqemiLH2d3ZARHx7KdWsPo5Pxb4xhbLvUY
DRgWKZckvXECUKm1xVuF0FNFCUdpDIGT7WPPdk942jwozP1p1/nhrdW73KJAJg4ztjfsif4QaHJ7
Jjq9s2LWdKstUxG+VlwV5bwtx2Er6SiQhQpQOyi17g1VXuXVM2v/XLI8nFF/3OVai6xXhhKOMe3R
I+Yv0VE/seRR7ZHTSLZb4yAlS9qa2aJjVm3t0vvuuVs/XPhNgne9RXz1mdz3snfo/Ov7k2U/8xJf
ZN4tRN3el2PmRLfso3bR0Tz4af3xSxGpPuqaeGU/7UKDxldc/UPEyF8vrSSYACOiC8f04FFVPWHg
b5BMBbnsr928Ye/lZPKsKamjiSwbJhuUdvOmZ0tKQ3dlw6f/2ucAd6bqy6vpPFYtozCoimHszRM+
jxFDVPS7V3ZWWa3a8sfVx3YY75CRo9bEnLVqVQNHHW1PiwgYyBx75+CXTi8q42gH5ItsJuAT+JVY
4WZH8jw3tyZPehtU0I46IQV/1nMOD0vjr558EujWImvLcY8oh0S8CUAUwJWSJ1hc2P+d1aBCz85k
16Flmr29iuiRQEGA1YziDadu4IIM1Ngmzj9+yz0w/blgesXAH+3+ZN6YUijPca5ik0mAmT7jKfKj
Rvb9o8w2k+KxW1EGTF5wyGW3rSOlZq31RJd6tVGFMc0n3RnLzeisgl5DzDlzcBaaU291QS5/s2fo
hDY1VEfXZOjz/f6Z3hdbDctWDIS10qSwh5rXK841rZFSVVSWJaqhWJ5m0aGBxHTEkSWD37hrqAwF
H/f4hvxqw2tdwdEAayKG/LT3lWQY3fGm9CIh7eWiF0UF2ha5RwTdAum3amfzliYiZ5vShppcvaCG
73fFV+gX3KB8kkoUff/UCx9GNpZw+KAXDJtx6PYIhXN3Wa1JJYGbSz5+LqphG4ad63/eYNhC++KL
YQAMJO7+Q5kTIb++TR6/+TH9qSt0iQPW6E1Gd1z/32NBOvCXEC684Uy8vXa33YSQl5OuWLcvJOx0
T86r3ernREJm16EwxSYR2AaSUyqvoT0c6FcI5c40yYdIkWhaMTwoiP18u4NQNAWcMJIuuNSYjXte
eRXdwXTCn8Ny+4r1SxN4dW9x/H/wr8BHSGjk5jRdycn1EkqmAZGd4XwPZA2zOIFkbjZqDwFeqexc
/JRfXvDkghn6JhA7dMF9MuCU7dqw4hJiD+bd2gW2eBL3NPfkUXmBzlY2mNBPyQaRwxsM3tjQ3Lgq
OhEcdYaRdg0+DseHND+2W3s5zIiRnauff6nn8/29kZpYSp8H7ght5lc+ADLS0X5HjGPE9iI3zPGD
t+M1Qpjre3pRuN2OHf3/k6xPpQIiexTxwuF7okBRhGoKehM0JaHVRnAEbTu0NfMBwgipjZssrmzs
++PXKsn6IR184S5oO7qpDQlc4OiXoaejjRDqMBBCby/eUr2YCX4TIn94A7ZdUkGEKQLgo1ERii/8
ib+DRzFTpsfjjJUoxsKutLaZtrEBWitdle+qd6KF5GxaviMan1+CHEh4kK7jU6Q1F2l0Q1Z/jDpN
2HDB6cDaJyjgMF2GFfT8wP1ZxXsaseH3T46+JnfBnQ+HLJpvgzqIL9qbC0VzjdJ0Yh8E+dV3xz/K
dfxbD3mP5zaS7+mN8ShoAGdjwdzzjqK+h+8ffyKVYujCCCt6p9yworPvk7pUHgZjoh7xlXIntbUV
8pkAkvPCBrjM2g4Rd5UMnioXmk6iILdxjJZfW2C16viphQD6mkqSO85PNCYhtyChn+qpKyJPP8w+
ANOEuOXCExv0TqHMFej9+duq5qBNA0zIerWhHR+1enKO/Ld04Nn9QnPL/X+pldJjCaq6Np6W3Ugb
w3G9A7yO0Ipu0SaIGBV9nP6X+9x30uVMLH98UyXL5hWx1yvHJEmLlLOatqLrOHDbn0wmEyggKL32
JF0I6Bk/6bLbPbLSdOUyC9WSjBjC1peq7Gv6l6PV+oIPvQ6HrRc6fZUlklDGtt7snTVIQQVCBLmd
V7b3ik5U34TI7qxcBPBSQ1pv5O4nyyjMz7pYcjuvBsHfCvfDAdLUdXe8i1RI1ZcFtYKDQKWEA0c6
wPD0EzUbNoWZuAfEDhQuKmvK/Q70LZk+xpSq7En1A7quEGQuEZx8RNoe4KCvCU/sQG4j9QNrCWYX
YtlgRJCsffv94xyTB3QDhbGzqdAAkVi4KBEkQpDb/oSB3/GRw0zoxBvOVKuOmJ5viIdmcn3xoW0i
LHT+wLDduC6FjBUt+DuI0n6VbbfDVa2dvK8Sac3HQwWtNZwXd641UzGkIXRn3krAtFt8GsNYKT0B
qqfKzDrIs5BDDBPTbAw8ejJuCvo8M8I16dXbT8kNaFNJOWnIxkTiLqg86RkXvSaHf1WdM/aRPefQ
60adjl3D6PAga4t0UFzxoIDNh6qNjfvt/uBdAUw2u63PEJRLBZ6AfnOEzCtgInUvuOZTlBvOD1c1
gt/bSAudEv32zs+sIZIJlw9aZTAPIrlJb+/KsDx2XYKUAef9LLWnnycWwfeX+eaydgwPry0BrZ+3
VND75jB8pCjFn1cQkrcLSnc7z7SfZNpzx7EZE9uwPdSmjH5rgjIT3x9V8FsT6zzXq7AH2rGZpNaR
LruhPGux59tfVHQYDELUGVdToWrJUd5CxT6B0I+BVOV2qGXQUBWi12iZcMAvYdnK2ffkidTanCak
nWbL3Z76MH++Of4fOi0iYNHEqXMFiLp9x+18ga7mVUhI5OlfII/tc9RjB1c5UVFRlWXi5EKKXFDf
UFV1yDrhVGwIZhhnHg5vkW9Fod4tznJfreRwqkCXc8iGT4ESi0TltCKy33vj4iVT5GF4Azn5chDX
l2KfHrVTcZOn9N6D+4czsGG2eZrcCuHfvlBzr9ejjRofpjzp60WsFKaxPzrIabahxPVEyu6ATTEP
G/pVCCWEbKmNifFMeL9h2HGptjHTzFQX/Pkw2kcWTDGPHMkynM/P/LPI2xUMVA5BrnfG3Av7Afbx
kqblhO+EJFtjYNfA0hDhqY4tYbGnV87F7elJTkcyCkehTvgfwvea84uy1Cn6twdrPER773g/5gJF
dBDpg0UY32O+dCSvvBwRNbH08J4Z1u1Uv7d8JRt0whxz5SpqCTkJWHJppzyn/14hAvQJj7psnCyI
zbpPP/T1Z/s+uNCKSLA1+TcfUFWFM1JJFZz7xSzn4zjbLXqwbULX9IZ+KmbxFKQc3lINX2Il+kqR
qL2t/kKAoKXc3VLGFbn55Uiteif8/sFGnRvzpWOzNSoTE6N/qp1UuY6ZM+tuXkv3ggf32sUY3/IV
gWgwg8Ihvi2Rr4jClB8+YsnKpGOQmdYGr1XE2Q3Uh+246BQKsGeo9R48WdSlrjCXgdQPGMW3i7W4
4RgFls2lRj3RJOKa2WrW9qB2ilgDy1yt89ff41Hqq18TbOX+DF+x4uAHiyqowJRtTMeMew98JknR
JsVPELGNeL5BBGeT4sJU0phsr5UU5hPHMcasmRheRwwQTpCyhoEZ/+ZItCbYUo2GiF00hnXpcAFE
XD9ASj5I2n63BmqYgJ0TI1QaoMgMMIkWm1qsJs1Pgf6OXhV/SuCdDeLdTOU+qdsrcqyJxSqeozNn
6i9IxcQ5uUgTeb5gA7yktJv2SInvfriQMFLLc0Q19zKc+vd8DQHADJ+FFG4UbjK7Vs13ClPmVsYT
44C5edYMT6uDLFR2PyxB6Z2intmA9q2r3HQNNNLFgA1P4xZBxVdPHt5fKF6ZmZes+8XUm4YTtP0E
16j+KH72xE+KVk6QI9dW/2MBFPUfsdywEWT8c9m3w+d6wV52mqz404LL1Q9TDYexeMqRQKDA5dcM
G0+LdCm+M38z0KBmzLVE44t2jjkhPqZzC1bClMotWFYQ51yJEUVRQuOoTqWgQ4d4xuL2u+XyCeI+
iT4t1/qrCcUnXborzfuF72ocTdEf3bzH3DkgDrK9AaAZCu+3Vsva2lgB06LJP+CGt39Iom1PjEcd
DPMCF9TzHB0CcQJXP4p+t4CSMBRlei1322jyrtzP9QiHXHDYsM5YL4QLrMYgwYDxEED0bBVG1iDc
xkmZixe8q9+0M4+VexfKaI3GGOyJyUkrO2axVwrxBaZOURBMAd4jBFr8ooeoYIbllfpLfxlhvhPy
ZFhkpGgWdcPyqxsGB7/WAb1dyzEpdM1L2Kb4fPI0xcGrrvChWszZAlH5rpMDoE5LlWd4LvN0QU8l
WWIpXbSImXR5RpIcDWM2AinuPGb3EGL58eDggrAQmphk/xHMIt8cXGW/TLgmgDPyH6H2XnfBgyw1
HySVRjZ6GuRY3ikatGf5DIKunSBTraS240mrVlnR324p5jBii3LbrYBwkw0dsDFaGSHAtUU6FQZ/
MT2LFVDLjNMsgggLOGSCgNh5UMMzqGH+LxTnc/ZOoFE8z9rEOyN5Z+8ohvnDstQ4JleEq6Qf12yD
aED1NqQzRB6+HSSxPXaYu0nX8qT1Y9MXpdHyTB4hzoJhveLTBQgAeTaLWb3S9uhkMW85EoaDf9ij
tiDSFykRtZ6Xw0QexwDDay+BEqQoqu5RDl1muxgLoFzC4xgiovKkOwon/jVdP9CXUNrBTlZSYQfe
KXRylu+YQY7YY0ON71OhFPGGhAJ9ofJJDTpJ3KzXs/9Oh8SgSZhKhIvGWxyjFP5E1yQ/wp8dj4zc
mppe117U/0w7AdrhxjZ2YAlX1XTjROaLf0dX3EDhXiKKP0edTk5lT6emEgyHEMfhqmK0qea3jp6R
iQUJKYntR30lC1HtA12OynzI/ofCN3yH1uknKTj+O0GjcuT1dWbmcz3tJxp8ha/ZHysYWt0sWhIh
bPwJGGoQhLRxDchtxmT+NO1p8nNkZMOribhUZQqg96Gq393QttNdjWQjduxYNHXi+e1AmFaOahKb
ny2BOm1T3jQhsLuXuudOrUCyQQVukCifh4+6ieBnp89casmBa+2LGnCfkPrSfg7IeeC5X4BNrgu1
FLdIgXY8oIeUGKMa9m3cpeR+6BOnCfn1SXybq6n7SJqSty09vl//W4G2vapqj98Ukd1RlaeDkF2e
DNmmvakzSzEHMYhbPZrD4Vj48E8bNl/zZuAaoHHY6PiPh3uFhWs6E731YJU6A5vSACAb2FZsaH1X
vsNVY6nBqz9vvjyETaFm8Dtv467t5ImGJLTiu5hInpTfb8UGNW2gxFPyBAIQ9565x2BdhhFC+x2n
nEdShUJpd30j7CZFDzVmRX5n0oPyj7yYE0+s5aDr7eYyixfpZPrV0kR5Z+Al5baXpxf35JXIUBv3
gyw8ekq6zB/4b/eI8pt4PY8ia6PKMCsJg5gEWL5BaGB5V+hUstQSMigLALGhnza8ztCz8itaqQL0
jwQIbHgN8/z0tZwoA58vOZbERiluqpmcBtJrvfQt58t9p/SyOfGVnFUbK17CjDiDXKlarg+5U9Xq
c8tG3ToCZUYYFQmt3eL53H8DarPlwsVzTdwlt+N9GMp3CX9lMNGPcQKvtCUC7s1kPRw+XDPqn7hd
7UWp/G2OURn0MSuQOIN6UEIptLwdGQnrslsucryaAEKEQnpq+Hc0QaD0GAdZapqZD0m8bRxyLwta
YJ/0s3rpyvKkQ8P5pc3yNHwz3SCEZaui/icpokS7bGcme5N/3zRM83XOisGTuYv08nFa2AFoT45N
uZ4pXr+jszZXoJ+P7YqKaJo5dCsws+kIfHiZPUA2UIoNwLCfNTSOGLZ4KziNHt+cbYmwSvL8fwSP
JV8KEjcKYWVMOYXnmUebHfRJdwWQqTS9KBzjzk/3f/LdqhbcjO0Vv7VEeETpuaNSCVe1X5UXq0E/
Hl6Gko9+TOKyMCGnOauPetuMxbhH4NLG1Z2wAtuNm9SNX6RtbavPhda3l82EU+GbIoFzfzBl8ZMj
yALubWWeK7KAyQwXpEvsquVnHnah18mfwSBuM+CH4gZlQR4CWcP0Q5lkn5Gox458PwJIxd7O4VP2
HcIX4HBqzFb2COo73WLlKuwQShElg/ECnyZevY0KHxKlecFT/HpIbCeI4PeHB2GWdk8wxh+la6nD
lmxrurZA/598ZIBbUWFdMPzLQlxPOi0xWdw71K/+JrXZmMPsJ9P/Flb9Suxx2d9TbFfWy9OFH2DW
9H6gnxF4XAjngvAr9Dnj59OHnE4sMJqpimJWv+eNB/+EBeruxxHMxt1/ttu729azaQekz2ZX1x8F
57YVKx+WIKG9TYWE06iA+0O+/fErsEb3zu85hR9w728YMLUViTV3wyov2DVh9vC02w525vhrqTqB
tJiiSmw42sgD6dfZNPB9K/y1Iv4n7HTNR2GzC95QlwKgIkio83CuFnirmq7b1uhw9ojvoZWQm6p/
I1SFEnl1i9tY/E2ATxS9Rg7RZdUzEWKFixW+PjncyZjwlxkX5imbXpaouZgtuD974wJ8VICAStsT
p5Znv8yqMU6Tv0ct79oHw3ojhCu1I++vQsktwqEqeBKoKZTQFb0zEbGRzbQB7u9lxtppkvD934Iu
JTwXX3kuily19KtXK0saZJeQiIkQrkFmWrQycJHya72W9KwJI7umeytPq2qZpmp5Kl9DqljUefR5
yam6KtbmwazA2r0OKrgabmBS5HjwsTQWEqncNXTshdaDGwRdsYtS9/CzV2yVPl81NTohK79i256N
UD1g4I3Lh3RZbdIlodrFAafPugYGEyF1aj9vNtntBBulWUEwZAyoduCtqmK6FZje3MqxjDxKVi5j
pC41m8Ccz8QJFhEwuxgweSelfXwXDCiu+zXgAnGLXOyPjbqGohZDFfHzNfv3oPL4bZLEa5NStcS3
8xY4snSctV3h8P0GxmkcFxcmvYW4KjeFNAmpDqVnCCURkmR+cvBTJ1T0r4qW3l0uQsQxAGLQcyF1
eOfWYBHZKh5G3ZGuKt6L3WNqNmLN0X6syKBL1pZLSyBfU+YY6S55N5wwOE0WdMqCE/1g/UZm9O65
gdZmTc6NkLE+Cjk0N4svQv5pDiW0GyFffixWjr+SwrxJ3zwonHtq2MUlQhFpR9HPmcBur/zLEdFq
i+8MdPtOyosjpHiDWBINtdoxQKl4ZPVouDs6IVUznhk48YfrMqx8GD+723kln2f9ucoEjvaiEv29
raDt6qaXR4WDmaCfokDi9+FvChT0XigdWGNMeJK6YKcaf1DyYYTy6UW5MhDZeUreD6OOqdCbNjG/
fuRguKpZjWTB51nMA/zJsiJmOm9wsrjC0V1L9dYtyB5y5nOl3/AJLk7ENutxp45rCjlyPj39n6YB
qRrxbIFKSMkipmQWwKgOrmzoKtsBT+nQvqz9r9SgeFbqmOCKIa5XJymVQ/0gRZTy1Hg6qTe0ch8J
lB3eNjVvjER8T1FaGJJpPA7pOfKRjE0OdBLvcAIUdNzVGzCSFAQ7h+nZ74td1cjOiMyKXoHew4+O
yakUrprfr8hu7Uuym5q4+MSJD4FxcVUI35QKubbkV/RJVMAmpNyN5CGYmOtkfKrC8rAFjuYETj4W
kIc6beRLsVDGfstq/gAlaR6es5KC2ICxou3iVSzP9ezWUVyuHQlNcIu4hg+5L0ur1pJNmETIcNxE
Dc0F9m7iTeMtgheY2ETx5ejbEVuB3wkoioMlIHfaFBmfa+E1fvPwGc4WXGi3tIVnzOl21CnTDO6g
AEuztoBBElXVykEBANtW5WhzTtnDKhgINSy5GJIGD8WSpMflRMWcqzjYpT9ShgRgVALSR1V0Ja7v
NdbFN/Na+nSoKCMrDZP5aj2v+1dAWosN/8hXfjxML1VajJhh3OSlSbOiLUbkpdyOmGn44U481WkH
BvdQFCDa3eARZ+ENFk02bnIWE4UOcJQAw5Zgt3YHaSC2ekg5oAnc7TIEk9qo51jSn6zFV7QA2cmD
hVfXcdxk46RcTv73FOvx3tZU4+hgKhgDTcVpnwrZeWyyEYOEnyWvrONzOTEaNQdkFAAY9kf7oJXK
EZuWFqy22ePEJgFH+0tmNH8MKaPHDDBQmVZYvVBUvp8HL9f3nRd+/RP+OeG8T87cIQMiz9aP3WF6
TRQV6YabhGdJ3IqoRT8CkKb8ZdFu4gPn8fn6x3K2p9QcWyfDnrv5xqd/i9gGlFG2riHBCMJAPR5g
oLz2OoIELSEeBD6KtSZPARCs/xf2VzHfnbShpmI+Sm6amX5AZIVcoQ/UUxWDrDV7lYiHbk10CYNH
GTjOnTM/lZ4qvm9Gztuqf1RL5AQCjsidGfIDYTdlgBZEx73KYyfCNVwDry7yMePkYFqICw5B5/R1
9MD3dY46UvLw3izEUytnoGLxdPlHMI7CgFJXy7TDFF7wdlJI1ce83/RI9pYz9J23qMIOxWZ5stfs
UtgFpe5ywhoyOq+JGhBG4wR/Zs8//JABknMDBs7LqNalCR0Xd1AFSHAcH0KyDh1TvRBRlrmc0vr4
W7aqqs6MGMmWtmJYiAkNehPLM2LTXaw/bAf4NI9LcimnRx5LYlY/J5hEJENR4uXd0i9YjMLiVgct
UwVq2T57W0SE9GjCHfek13cXTDi3n1RMKQe7oHeU9+LetWQJ94GO0Fbd9yPdtSaTqVVw5OOCsPiX
glEmujwfT42V+M9PKKZ+813UuRUbFWyvBOl+8F60bD77DRKNLvUUe+lrnGxeab+kUhSyiKIkerXq
oc4+ofcHYrXmYxrpAfhYyrBEx3sZ4ekxjGHt0uI3TF5fP7rYZ0UVNn5kT0xheACJzBP3VkdpN9nF
PmZBewvm9rY9bP71mMVXJR/+PGu92TzEZyoySoCxG4Sxj1jSXkz6dFj07C4jWTfPUajeliY/WWzF
TNFnlr9/L5+2SOGX0DDj8E2unhMdC5YXveO2YpSxrC3vgH+QhhxQPL3/rkOG4+V8ddKNFhFqkfYe
y/mFMZGURsRAg83VR3ssqB8EDZa6nBRS0jMXv3+O/lBcQPY7UkwdnEhGWvsHZkc7FKnrrF76Vohq
bzpCwR4srMvK22GEyfpcD6S0TZY3TM/zdEEMy7xaPoK/vcP+KPbCxIOl3VIs15hjBE4ZyJvC5u0T
lWCFhPYG26UINqIcq+fCx/kCCFVJJzKdZ7n3di7R0xSEpZkeaC3IgF8e+1VBfpp3mbDEPM+Epi5O
qvFL7mtozf4AfHzILj0MVlaFiZYFlxmi7XpI0IaqxazEeU1Dpx7DFfEKNtmkYemsCllX4TE7xAvP
1j6ZiHbBzsdyVNpVhTYL2NWnpYpOXfcNlZCp6WfRcIQ/WpitrZrgQbJAR9nYrt7Hx0TVtaxQ5qOS
Vl99kW6RtV9aDPXEGuvMnuN6JS8gJRbnylRHOmgRAXRmnNWv8KaOQQ1y1h8mivgeYshMymR4E5Cr
SjKvGxe4/CnNtnf5dqYdxRTRSTZoC3PdLqKcmUTCYSrLVm2Tudvz+BEaYtgVAHLXMEXNK3Z7LhpE
9pIUZYno+LqPogxZJ713MCMvqRLqyce7obSGPP2LeYNEqPd1Y6021id2YaFDds1bTW2kznlRBpsD
w3F5N9h0FW8xGgBb4e05Y1z2SwSVhJ0kvBBZShzB1VkZZ0+sMC5kqvILfOsEcPTDKW6TJvpVu+ip
ycfiMp0qWcYkJWO++c3PaL/pDFEZhUiQLSwQ9MHMc0xItnc01iLPfycOnU1XRsfYj2DlQOABrVBT
a5HI2J2D9luHyiXQZcWwPR7/xnEbPq2Sx7+rhVtzo+XxAbXSXkwBxM1vwrPVs6cCHWiptbAXXNfE
iMt9cevlf3ko4tTNxPHjqCrQ4ORgR4HqwgK3U9/pl3655/K2nRlJqIKafLTT4bFqB4ZxoM9HrwRj
/GbAaZ/iVzUqelpcuA+6aPwa48BSnMd1SfQXVQiY2ydlnmiPRL45Aoil/Zg/ec3YSab10g3tvOxr
IvzSQ694TV2WEaXd20H603dxfN2RW9F+c8HZm2x6gTSMXOaHw020Ri28TzYZuxbzLxC2jaavQk7/
ybSBFdGg7TUg5nBkNPygGWChOfDTBEDuLPpNkUD6MngNI70HzOAd7qZVlCqfv5p9Jggs/ggSnxnO
HhVY7CnYsLBRad41nL62r76aYU7KZ7TBJLwdhJuBTxbjcqz0TzCp/SSGpeAttL61RR1Ezy5tlymn
mLaiwLN5YEDU0Mw7dI9ki0h8edb70GMkP61iBTIe67YO0ZeDLV5nIEc9gvTQ7oAFOBOzb+IbLbGo
IFbq7ilFav/rAVHozASZvuomCxJHs2acOs1fnMTlW/3De7JYs+lOR474cVWX7rejNGA/Bl5BH/nQ
hOaQAEde7RrJGe5oRF3QrqZkzqvPzZOMFJCVnd/LcBz20UXWzwsBgMJ1xt+g4ncp7TjdU3ZAkMbA
dXykJ6FgdCute0idwbhwsO7yQsqfh1vXcq/KI5RerBNXc1Pce0cb+PignCQWO6PAjxM71+r4b676
DwgMHR7sTkfPAH5UOfCi/prjmkWhz95UXpysPF6oBtcNYgZESAIpk7J5WTlEZpR9AhOoURS+f/+7
0WLVoeidIOtHBJSbit1kPCpRjoCDphsEsvj8fhS9zTXrkI/VbgSsHs8F+Hup5/qyv260SX6zLOzf
r765FAtTXeDIAbn6s77Qh3bJwZXfzwGW2IB62J9167wlgBTCvpsry9jQh0CkKTqkBmADnmLDu7qH
dsKCHndeVjimw0wBsRB+YNzp5XS+HTzSwW7MzGzKoiu040ZPD6j90Axdj8HT35OwX0Q19cmUAylW
GcLpB9yw2uTMnSyDXf3oMHDOxmG/OnYrkdi0JJ48uH1iZbZeZQBpb5vce0VXWis8slY3idD/9uXK
lqAMW57HfxFKxZTLITsXIqnZdtiae9hXciOyCYhW9MMyMPvVAsg2jXpqO8CTypaQkF7qjxS/x31J
3YARlECt6N+cpa1WpnTtcGInAPqY/ldRwLn3WIBMwSEabbfiw0o/YpQI/r8C/gDYwesKu/ej270u
6Eu6NGWnzYJLd6E6KkB7nnjdzYWC+MAVDwxndB20PFUDVRDD/Rtl+AIkAEzgO/20nS0nVjAiQKBk
UT+/4+KFqdjlGb6rxFgvkLNd3TKFPYTMc4UgfZi0G5A89IC5vZDAyGVIRO0Kh7SEpuP+IwM3K3zA
81u08tpS0kRpanXMF2Xhtas3m104MawLu88WZ7152fhQv7A4+yv4MLim3vqJnU98IY5fTfk4hxoj
Kk+8PX8yq8Q38jG+dWSxqFFSdXzGyzMVQpgdu2j02p/VORNU5rghGZ9z+dnlcHl4/ZquY4C+905W
rw61s6P/5+y/iTCisnXJAdxBP13mDMs+keKMHfeRUr15rmKJRUkMg63Og8txRQa/N3Dsm4JSJAWL
CoMLYRJO18URfgBRGWk7ueTkhD9R3GL3t6Err37embOYOFC3H7cZQpfAtlr7z1gVuWkl9cXgRcWt
i2rUp5riYGLudX4mbJtiZN+wVHqfRKmVlKxDXbx1T723BP6gDwztIMUlIvjQWUCfDhJsLmu65sDr
1f1K2kKiMNgnKCYWukYnHwX0jc0nzIXQK6AB0GSlkoAM4CLKz7jCq8mVmhW3YEp6Msx6qMy8VeU+
xVGXombhR5wb4p8iqHSxynutZIxndoQfwiJ/AN22WdUZMziP9PIuIRa8RYHiayip/xiBKyUtrNsw
y5y9GC/V1VrHTRtc4Z8yuihh4IPbaXKOOjctTkzehUX1mVZoH5ATpzJITb+Ii4wGbVLZLKFOolGS
pPwhqvmGEBWh99QmjvdL2LwGTgKw9zs2PEYb+UbUkCsdShKpfSOgdXEvU4RnpTivG6Q6CcueFOy8
gWJfwXjgwNCPQLehBjzZg7KvW/HZ61jvio8HFMXzSJzPq73k7EPXtUftqe4xpb7wuyFr4BsR5YH3
pR4M5/o54GcyXTHloTxLnf2dOSLtQ8Ot412przXlAT7VqdPs1FxbR7gRsTVxuBXw8ot9ldNmnEhC
zDmTkr5+9P8T6MVIV1hFnA7A43TLWU9jjTNkjzojJBDrM+n2FMqwekcX3o0mpP8A/AW1Bn0+plTe
L/6+Gr5IVa6m/mKVKJwqE/OZMffVM5dShYw01GdbVObLg8OkHXFEA0RCUab6ATWIQBjvwJc5wBw9
jiM/y9Ew4m7a/rjQE+CYXLt9FMtwEf6fZn8RW7+u6iSrS3/DVDwpF7zJU8HtguhuUpuyJFvyqi4e
2fv9OTt7gO1Ub6nOvIw3OGQ1umg/S7qYxulDX0E2RAU1uIwZOr5KZKK4wZgeRc8XbGytpK7fkwec
8TNPO2a+3kmKzj8qYaBTDB1M6j7imKDnXx1XeJUqZZ7rVQ9Qe4/s6Mv2ISO/hB4rumPnwSvvnT4Q
EoyBtnw0WPKtlQMrAs32cJVsKi6k3RzpSd2Jt1ZWCraGih+zMDtZsjDr0FRoITugYuo4WNFbysgJ
IIuqW/40zn5PQ/tHcJuq61TdVwTviD12E5WdPZMT43TuRAVxj9favfHZ4Irvd6YzXvbjSexahFxm
ORpFtO0ywdcl3nJCpV1vyTOCqQRa6WFT0u+XxVNI19IRLjgEPjlcFYiXr/gW4/RYvlodSMEt1VvZ
a/Jnhafaor14aTDdtVJm3jMr8xbDPOXq/rPbn7FTfzDvK35AObCfxAJAlx0/L+fKwT13wE/hFHZj
VaUH5CF9gl9ithPir2CiFtCdUXEXKfiiqBA1T7m+y+lTkJy1bda/3w4Hpr90w1w9f2LIIC8MkZWY
uoevb7F6Ii0mjph+65RGN3sN7uVTq0Vzs0Ue3Ejn0p4ZAcxjfAZ4L4XFZekOeMXOCloPMsvgKOvo
9JYcVQDK1g5FpK9j4Jtlv6KfjNrfGmsCl/shHuCCbTAep0beWbgwzLbg/rlnli/LuU6WWdAmOxOp
wyMaDxLoQ0UG0GMyWnP5IP+l/EaQ8hqc4nmvWd+Wg74lKdltPTbMQy1rSy0baj69jQKf2NqNwyM0
dwbShgOL0FbYut0PCAky+hOHdZqbPjIKF/BESqAYnDwoJa/euyn4CMTYtTRNgI7cCIDOmcfLHVFs
ugM77i12l4REziICrbLO+LkamJhrQHwDbrTEj+SwXBnsWOWqUw/RJM+/8bEtKd8XSvkuxsS83XQr
9H0j6qOpl5bz1kBNCQysBYeM/4HMI+Hl/eluKDqRRl/5SXYOPjRZTvGh4AbH8VrIn4d+wuB2bNwU
bziif274jvZvIC8OHMxVkAautb2iKFn4RprkGAcKA9FTROR3om6xIDiebQmzGF4jmIiDgxhGKDvi
1AL33jQaXbfalKj443TH6D5kkH8qXYG3eWzXp86JXAGqvgL+DUpiYqN6Mo6SZmBwiMwnUqoskut9
QDAFBu/OGHlfHwdShPgjqSxGg0PrFxwZlLpztJ7fSqu+IVzUq91mNaa7ZsNfsOVkzW6c7P/a8VRp
IwYMZrnhUFNtY9lZq6FRYThzkvlUs7ziEKe+8+5F5cJOYDe29V4GQ2WEEup5HBK+ZGahd4AXSAgM
OxSqAcpflTqxRjsoOW7ZZTJRcaNZnRRR7F5y/bgsz5qsMOLWdJ/kOPSyk3i5dR5rP4XxoSm/vKVu
mpgTVOBGyaFFpPbnrl4EE3MIEp9ylOA7iKZu9ugShxl6ZaAUOZ23yQgYMNnmHxx+dLZ9BQcKuJWJ
5IVlaZ27Q1uv3Vj8jgh7GFR0HscaJNPXd38JbjgYxjbNAiN1jPvJhV+Pldw/58lGYIWxEwSrsVil
DyUtWUTPueM61wqlpnbZURQjWsGIInupaoj0Ab1RSd4CWWE1idxfb9UTB/YvroBnqZecmuBhFokk
3WwcI7y3K4OjvwjUzx4GSAmcnLCSQ7wGgX+j8+K9oEXTqFKjjII6eR7SFf0yRZ4iwO5dvxSf0ZRy
u5jLqOQQ2tmsFN0PEpzY1+rJ/5O9EN/3k+R0k3ba0GUweqRAZugIyqqs9v69e94XcIv9L8WVi1DH
ANa6reD+obscX3ldALS8Cz32kjQUkg+evqSQ+QuSekCo0GMIRvGv3SWBErBingU6rlQPr16LCHzx
duzX/IM0/COLyKpzHeo8by/MSFHoeoRwT8uZBfWBVHGBe95gLLBPGeU4ff+ac5GjEEONFyUGVQai
7Yn+scRiE4fbjnevY+gvFpm+lUwcKXRyXCk1q/p1DiZVwWx97XbWZlXtSYBOcbR/N2B5kW0IRIQ7
Foh4OblPIjiGUU0Wgr3L9QmFfov1yI5VsUvPyYbJZYcUmNqV9hiU/7dYDTHc2WlBR9JLj2Y4WnYL
OKDUgNVyaMJs3tIh9+yBlshujhy6NimHDnG2PT+zNhO2rWQ6wdYg1K15kHV3Blo83veiGyZqanvR
QgPlxRS2uXxYQ/wVxLf+Apn8IRzWP741EyoYiLVRb8v6IeeFi83XSJY0Slpn1DJYK60Ts79ZapWK
gkaOV64cc2MHS3TE/CfblHQvEGXnz+fVwaS0lsJUn/Z31AmTmdMlgIf670E1G5JIRmBoKnEWIGI/
B1dPtkvSX75q/in7DSkk5GNmLjO6+w360CbHpAfo5dTmK5EDX4gbekmCdjeQEeHvToDVZiynTPDO
WN6VOASNHtXKNwRBPVy1QsUDYs0lNoXB9BL+wPj2Kq9gaS1wbq89X7x6ttPivmjUSY98qMqVZDXW
P3CbNDFKvTMhwYmFhHq2qGddFUWX71QnFhnskQoM4thgjTWNaOVcE1U8NAYvwefFULfxOis1y7i6
DmHxRpnyykGuN68MkF03nF0kpd8ogKqfGkG23s9sHas+p5OQC71UgTgSTx4Hq8RC5+T1wuvSQuEp
hgldT39/r9yoQkeflicIXhN0EB2h8qO2edEMzOu78CmVVqEoxd3kbi6ZUfi3qLXc0Z3AczICHkj5
ghiVfKsPKnHhdJd0jax51iSIaHGzXtPD66DAT3APsWPkJDYMO9fCY6kod5clcKVothOS7XNtl2tp
EiGfxHJGFdHDgg6Dyn9eTke505pP/3xsNXFSjuhntMg7AZSRpNUZnjGZ/vc1xx9cqgJcR6yG14h8
IhJLmvpBemYURy8BY6w1SEpVR117f7sH53Ed8wjLsWm2nJ9HxD80bRVo/d2V4YluwlLTgltf/0Mq
Gs0LfqP1BVoZG8zTSTERJZRxDvU3XM+QzVlxwx4U8xSdwMQbzw+kgMyjzsfFi1sC6wItjg290UGb
GjotSbrX/WC/EFMrDNh6O91n/N7yrVeMi5qj+hZDOlKGs+hNezO3n4INsDcx9u4xflFd2K61pexT
C8iqDq/poUj1IKikgo2cxfR1BHe1ImKOTwBB6M/nhzuIBRm7yEbWg5cIyDPIR9c1ifCx1nD66lPy
GtXcYEBvsQ0EoUblnORjCAxiAg6Yz8Ripnhy1lF7iK0BcCgY82rAZdrGp6Uzo/UL0C5wHip3vkYu
msM1cwZIiz2kk40ePu+Q9cGy0YTyhktj9WcLCtHd6apoW4lXe+r4N7BJL7Vil0iYmQX259KW1VqC
SFezDHFwkd2tlXxOmcCwS/Q8pdVh1iSh3zDAxN7fJRFT1wesETwIA/Cm1jYsz+7yGbhDLkwlC302
bMBvPLV1erkLzs16YKVA0mSeu5hYwkywm2IPP2wmZsoSMmBDIv0Wrp97U6QlA/WZjdNGVzgvbfkI
6Rq7YMdJo+kcVKu+fypZ1KnHHcdTKeNu2idhVZs6MgdMAxzRhdo+h7sl4Db501uK5wuaVekuANam
6GdACsuw8i/8AzETu6UAc+R4vOaggHhzv5IitXsTsg/7+S/yGU+yv66gAsSbJKvlYoMgxiqLK8Sx
Uwaar9hgrsypvFb2PPbCBup5FZiUm+M6M6PFHPVKEDkyfcrF6kUlBSNpYM25LzAkGFSqqJ/Ez4j2
CzEPydoeEaYu5eOEdpyaWXZqlhU0kkHih83+bpcSY98hSDedh4cQX9BiImH598TqZEG9cTxqi6xE
PhgAhEdjJPAQfZeTByh3LnKf50y6Tf4ZiRiIR2VaLF/08zkzsGwcOzu1H+hpOAqanzRKs+OUFA60
HydOD40hGiEVciG/Kk/MQfQutKMjoR3j3m3OWFhoyFoqX2qMMW59ZxvfZw9VNS+9DAyUruSZs7dr
xdsb80ftPskpiQg0rceQv2ZXqVH9H/A+wkWOeHTbAVpuKIIqxrGUytd7Wrh+lDCA6dBh5zZherZc
0O1ZsYvHkEnnTTpXmEkVMbKU9xe5zxoFGoH1egNm5Gk6jSOxeXJakGdfnmVPz3yq5nzdLh8X3KNz
SqsgnH8Ogd0nffkoPbRL7Sj6xIoxClaU5W7TjsiCTFmksumjP196mUpJnv0ofLlcpbljE+8J+Rmd
r/aZVP4VXdhPMtpLk7c3Srs699OAzzseoqi7Blimeq1YZNPNxqQqm7aHej6H3Jv6Kf7Vc6Zz5q9D
mWXCizr1xFwMp1AeFw7MTYbp454ttnqIT1FFAa3ZMsHsfOFjKgnINtGGnoSyFNsD3HBh4v9CQ3As
ftwB1/a5/4d15m2wwuHsZzheylIiK7aWapT923JkixArM8SjhreKkwTJlJH04sBF8sgFAR+J2701
69JAUnWQJb6WCVlbwLo5KBEXncIzv5riTyCDdyz5vesrLF8u68/PN16J2YEPYnKJZg/gVMQD8Ik0
JXTRqpysHf9YGEmgyjuuz2Pz5vbIJZq+T7Y1sy4tAG51V8WRjam3Sopl9hMsNyJvJ/qGsGhHjJp0
GtcHskeOcOndLtMWor/qaXbhZJJCT5nxlqskY5U4XZus0eIJIunDWgtJwgKllM1SsnKjJ8tOY31b
0CnmiWmL9AxYcXmRDcVmPMBNxkVkdcI2bT3IEOGBaR24rxXDD7II8H5P8RS48mfFIpcCghKQNmqx
ShMWbnQzzVxv198NkkH/5gt8GsES6IQeG/KYmkfD1Fcy7SiMX8ncHcxoBGT7MImtdLa9//22REXj
e+AjSm9gZZRChwK3zLrhWQH0aecMX+X4p7ar61gi+OTwvMCNxK7HDnqYBn2snaTk6b0CG9+wkNxa
jaBo9GFjUgnHd6Zdlk/kUnO9BbnjOZCT+N+g2zN2D0Q+mXGrfCFDvfzSnTFqPJonlupfoIj0zIZV
H7uZ62w3y4yH/42YxzHBrqG+SoNPoUoufVhctAC2vrLKL+wLsr9QtV3JivDF7IRgRfKhqFPMF+03
R2okaRyW62WXgvW1nqgz2LL5xe90yEwvU2oBdL7OXp25fbiIiyxZYgWBrGYCnxG4fvvLx65XXgkU
Rdw0tnNrw3KmvJqXBP3W3A3zgZbCK9jMkwV0ELOrTutp2waWJri8cKMJ79kjAZ3JXbt+lmsMRDUN
6F4wSwN1DhqKCja+BcDX5wsptJu8g8O3ucqx9aN/xdj/0ZpzwNE6tSdtee8CnpGSrS7TSbIzGFE4
RxoLT4vbzHXVA7hqgMeAR/pO3BpHWxfGDhcQ/8wBDqXjS62CC0myu+ZYScy19PlgYoBBHhgqW2yJ
qJIO/AK1hZPrAYUTFUmXoUFd7OZ9S5msYQdYB/UQrECszm/3gL81p5qckD9r16R/42nWyng6TM8d
KOCmiERUCQG04yOC3cewtjKidO9c8fTmvm7d6iiHLySWrl6RGDoSBee2LHK+EQ6NwPpyRlfM2mJZ
UemDCh0dT0KtUeENTs7+aJdCgkny8BnfYGcWlJhSoIAVc5HaltIicOa78lfZx+1E77rRWmeU2deW
mU2e6Ej/BYdzUKDbR48L2DNCwE9WVV6hj3tDoHPIxgkKiC0+rVkBZ/VjJXpupmUk6ofIuOaaS+Jq
NXQBPcs7JvF2+aYKhbizjMO1fq55gC2oeHQgyEZXIpKugxqDlM1/7sHQyD2Vg0s6k9P65kmzrUy6
WKNHgncCsSn/scbOSjCFaIWmfDlJssI/cvwuppS2zwvJO0W7P7A5kp5pS40mlxEIPrPD0hNzAAS0
WJlH1NGJ99HwkSKkoQgU7VuF1PODhO2EvrN5a4r+V+wFdMMoISDKwalc8P6NL8VMpS32Hx16dfzK
KePpxOLeQSL5jMpFLepdeb5qUXF4q5SbIoieE2Hp2JqAzLqU9TdU3SI98DuFRb9bBTglqd2JEzGJ
BChHXxSmdIEqD9sNvv7VOPrFg8hUr9jtMFKNotT/0OSFrvuJxhIknoYhjzUHK5OYtE6eKe4Dfn9l
MMHVagu6LZ1qCrnhBH1cLIR3zXzrSKyclAggnjlqb7Sd+FtBH3Yys0CiuDlYAAzHf5rMLkdPfVtu
9Q41B8txjM2C7jPRccELcemCC2UZUQQ0ZH/LGWjgHWiwaUqnrbc6Ha/O/buxUQs79aOD2kjbl0wL
NvjXHZid/4QxxgGxAGJRRsHzltRRDGxJcwurwqbZ9xo6kjaagbRKm+SRYFQ94J7u4Xxzs08eAv6K
/CaDTEDYrHcCdzeEzKHlZ/jBXFvonfG0JSj2t5zQHT3CHQLj56AiR6RNQ7M/IdFsmCm66DhF35fb
RhlPFyyg4fziphwJ/fCnixYJQYKtbQpjc/E2hksREipvp3GMFvrpWtdaA5QcWulahM861ZRBlx75
Cr/+TgFpjmR3vTdk7rl7QoZmOvYJ3d7Os8DFD7ffIkjAouiika0FZjhH2GUi9o2ubz4Sl+b/Gov6
E1CwE5NvctFjwO1wFPy571si26BXlWfUsHBxVYMBAmW+9zVKnCGChTH3pdliky0JGfXu/en+wMXs
cNng3ytHmXwPCvUO4oWgJuJ86hsTKv7mVv3YEb+bwTeNR/b69+atUOiaVm/2AMbIlay/HKUZ2XGj
j60R9pqmOfbt+zka17lQeXZlW6KIQxW520cO8PMpk9S3pYe/uQ26Ts0xqeCX1ELBjjCtNl3ran4l
mTbOrCTm5eUa1ilSOQIpjoEqRME5ZobilGKA3nZN73jTsqej/59dzj9HisaHFjIL/QvBhLL57RHN
/OdyPL99GU6MKmoacwUhRja9xmTskfy3dogGeIqoOQPkquvqYDYPEZpgx/meaC4rTLFRm3QY6DJy
oVtAiUpdx/eNfsYMpNIQgOP/xvl2LR62XJ9GZtD6z/f10Np7Am+5m+uOW+SRNbVQcT/sdAcqZLk5
7GcvfP5XjEUxZPh41yg6MJrqGUcTTdYvozG26jiqXwyzyo61md/egkancag0pFk3piH/PTD0vVgl
6KKxshMCnB3fL1Ci91kiIo2b3d3tTWdnfN5Y+4z4wHLRubTIXvJkHhLl7UnMStU3UQPGYhVe2/Lg
u7cN8m33ibIfQQLgxP8xfEh0J/3MTDbitzRIV7pUhpgG07FfHhUj34nSOnj57GTpqsPCLd6m6pLK
+bR2s2TzjHnwobDz1lBynUJl7HbVv+9ZYKDTHFajyy+BcEclCByQQ3W1Q1mJk+G69+eLR67Tmazb
MCeA9anwzborHjNi+JwPbFQ3+iXVK4WrhwFBOZChUUU9wyQe00uFGFdvaoOtjiy4yDuGpnBaJ0Rm
Wz4FhIe5ixv77x/y2I1vKFGv/NBRSHM7HbMhjFw5t5vtf4YeCb5jbTfElSq3RLT4yECQ9j/cn7jY
6s247o3CF+VN5inR/oV9wV16Qcp0KCXb+4ZX9qzEwStbSOE57saoJuoBZJ6UfKXjWwPZSt1Nq6vH
XvdhpkBlDCn3BphH485Zik09hdTby3tfLen0Yn/NUrKIVdYSwOUy8RupZjDT/BpyHuB9NOgiHJvJ
IqY0R5OfRk+MlMSS2rR+VL1J0W/cCP9ZdkiiXIhL4cx7mutRabX68Nc3fLK6YpXUSbhwaGzWAZiV
/KtWu9NbX+n7lFdKqZVTbD043Vtfx5O0VguqM2YU1/DEcY8z+EaMgGURzl1TIlHMyLSm+QIi7Dpg
XD0iFRxl5BrN1RcQ+GhRT7YFtyAN9r5yFbkZi0Iv46rCIRsINmG8YJ4Qzpi73zYCKQkzYnUXJnzq
ZpLvPufzmyanjBV06qcvG7Th5EaOt82s0zP3pX9xV0XAolJ7J3BYgPh13+M9gGDo+DgndG/PP9QH
OWWIS8Smkm1YnbHkhy5yBIAT+0wdW6jmG/hLKhghk3+5gU/3pVoo/6rlb/dDJcg10O7O01V1Fnj4
xndtvhMtesYffJ36kXLaQWUXpBeBOj7EsIpzjpAGzNDFYz4Nj+Pfb/zpi1Po48mF0Ozr4av5eNgf
lSqUJwtQGJ0t20RZ2MoAfkngcAfUM3Te2hKEMU2o/Hsn0pzt8fhmpoS5tbJgkJNxtLJaGjizIUOn
q5D6VFe78XkroSrziVsYNitd8GqhNz4E1iNpj+Bcd94AOxk8RdlFpffLp2jkOCt20xlr6x7xfoMe
cOSA5ix8HfxDxiiH7FuNvAN9Ga3A20/Jc64BE/O+CHAJvCSuGHwtwCHcOFwNIO/9AjOU/i6CnJhm
IuOxTTV0joPBtZkJt4k6u6kfSD1NYSpmtPU9lGZFBUwWwp3ow5TiddW+XZ/Gsx+izCQzG2hLHIsC
eYdj10r4rT6XQ2tb+d/Uu2HTp/bxS9vnc+RR3AhhXXfYkSpQDJ2v7PWmuf78lb27eR5Sd1MtvVGK
XUiDqrJoc9x1MNLtCDka4e1Z98rxAXDQr8yvPGbBE+1LdRM1TF9LGPRDEIrz63jlkN6oCx9A0UQJ
yXyEzkJwrUV5c0wkSnWpm4GH1wv/XJ3FIksgZIchAIKx8ERNGSoSKlLGJCFnCKzfmVBZLsMhXbdz
qJd4ewa9tfdCaIyzJLnU+UqX5h+F+P4ZZVHXyKF2EgMiq6Z5X12ndsLk1NqTRVQMt61N1l/6zcwf
0j3wabMtpm0Prjv41ig+mzqNCZb/gVjuSVlw4x3LonJY1KQN87mUooo+07R6fozZso+obMKX3jHy
h0tI6gTFC0kTrfVD0RyjdABv7UBIZib0ud44dxWQLBjrmG1wdrvjS6CrCjxEY0pKp3yl4CbFkXsI
719YUdeqSuMJ63scNIUFATR0Hqlgy3mdYJgp0wEmY6nIGZ2FqC6NbpV3zJGxzrc6+oPvJX+NVr4o
bsTJU26LPo1Q92qQLiAtN2a2q2NFBpQXKunGREZmrxjk6c2Tn5I+KwJbHF6+OnjElV8W+eA3zzXw
JOVPb6GITZYRVDkUqB2WaGkE6FTb0EcitzF1qY1Q3GDSNf9onytcxO9UuEgoEYH2fJcVy7LdZWkt
DzGQ40yPTEFlgRNxoDDp1plhxr2WSGmn71ZKu41KyCDcxgtIFzxTfpXADurzZ+8DVtl+97X7i6fV
DIppHFO66Hye/iNaVp+CPTIFp/NCtD4hndlRRC7A4/dxBAejPTmkbUlRtO/ZRUe6u3jv7Ii7b7fC
8NYgOkC5xbly0+UR5s7PtTlCVUhPHwMLX4QkI1DYlQFaOBnSvP4kPd+bT0nRhhbcdttv0Zb0hRNC
HGb01zL49s2xcf+2qLnYEVpnGFft0lcepBRJRP3g1hq/wR3F/PGnUMKMaqbzL7s4iBJ5bCnCEWLU
EVkddLUXi+Aanuo3SZ3GSJQSrl7UBHtRM+QA2zr4mUUiXThjOhszGjqoPRnwg99HgyWZGHR4kBuh
ZdQ4Qx2whG+CtIHAKNE6wSGmVnIoxJsTEL7gfS5Qsv3wHqoMMI6D50poiEOXGja1ojO5ixhg42CA
FkM8zrbuysggpKepYoOBNqu+vW87/+WVOahRZgbAUuciyVye5Z0gn/ruWRFQ0U/DXI+cVuiImsCx
gc0+45HV3p2F8QFXAC+Ws3m+d+xVw40tUDgNYiSSfMcV0glO9+TAh5N3sa+Vznw9uetQZTJ8bQ1D
NPqQVMjhJYhEs3JpaE8RO/o0ueCPo1+mj0UpsWnU/t/pPPK9xuM+xuhk+1wuSyobMJbo0kJzvnLM
sxC2AR2mXO1FnGQ09hEzTe6dcFZc7TDvnIPR9pF0qxfLjxOvA0LTDaORLaG+8w6o4QlicUMPqNhR
Vttn+6Fbv5BNuGE1Q+OEV2WGvpcy1FoR9n/MtD0E0d7YOz4Wqd52eioT0hDwA81olRgVEyWGbt/v
6Trtj/DavM5nkm0MzFt1jC4oT0QtZyggLCpzrKKGoY5ntlr8Z9HW3X3Uf7+2L/jZwDyxXLqWVWkX
2bY7xNExz/x+JIiviM6noQhqwePOIeS8NokTlSez61RPzV1lMp6NcpmnYjirE9xOj4U9LQvkf4I3
kr3/l8NtbB62Nk6aMQYw+ivf7yk/34B9md5Zo1y6ZNz+YAC7G5CLpTepu0mk0O4qqY6ZcOnstK0e
5fsAujhK1X2iQngW35NSfDjpEksERjyuTk2BnjlR4g7s04nKofFGsb2fKycaJyz6J7PaBh1+Wi6e
W8xu8noF1rvuoug/R7rGkcS11EntBl7olDcUwtDI+IlQYY7NABZyoRADmmbjPPiE/vsesHz+9mVC
TjUnyeTI37ao25dnn5QvmRT55bonWXRp401x9LIsCu1iA4niaWiuUPcnfnzHooJmS8ZTsBzeRXOH
fT8IL8ELanzE3NrXB6KpDMwK8YN+uD/DBi+0pDokU3Jm7Pmi0PBnbH5V0nHsMMqOPU7m9WE9BX3s
RKYrIYuV2zFpzKphiFYHZyZKXxOQT98rffIO9P+N9vULuk+Vy+lV2278ECicuQCpHZ2jdDc6XfBk
Y98GjGWUSPr4kNCpGuH+UcsVwg6uSvpPOQtcxXE1scxl0N+Fy1O/uBMa+yB9cPkJCxBbAPDlMnI1
Jbq/CLo4zeHKhNclUhZfcbxgpT+yHfrQRPYD+f7spoyy+7mh7nUSwqLKFAf7bERCUCvZMztCxLea
xWx6ez36LmkEejnVfCaX8QrMJhmyk6XuHihkWkaCOJyj2MW/faMdCRNwJQFYY+DsWMIfK9vkH1F7
419Sl0rpknLpSmE83bz50UKOab5yQHa82sk2uNWrtRLCdfnV6XqU/JnmN0iK/56xhIrlyW86+c4f
oJAQh+So95jkJBW4nE6wzkSV4yM7C0kioNNfudSGXCLNO58p2mPrrmnpE2BOTSTY22RuzkGxqfNd
Dahz13pcnQ+7crajQXqftfLtc8YhpDJU6sABnJ2fCKCaxJOSHNcpQp9DUQCkLgqxrGMwfTURBC0G
p3mGpFrlD2MTQumZyEU9UMEHa20Ce2dvltxr+VkwXyt0iN/ChvYdv59zxs4dYWw0PVsbtAWgpYs9
FP7cdGNJETuBs90grUeKILnkFzONPdNeM74HDPJd8BlgMajXF10BSXi8RDy6MSbDx9q6pBqKqTRC
yi1FkkTRl2OmxXjxLJkv7owiADo4gwyROcMEbQSTsHzUNbc/Xwd/tQfCTK/L6L6A5/Z1KR1baMdM
kOgqNzRofalQoCuJ4VaclOMOiAWrPCTRauddjGuSl0Pr+0/CwUQQWRHFjzWXZjYMxfNUVf1QJPVR
/j1sdpGV/YI4rwusvkOtBWhMBBnu1YumD9KosNVaPKqdsHBVyD3G411MKRPVC3CwrIzubgHS/IOd
vpe89w/yLulAppFconuqMweMsD6yiz0UUXlgxnOADFiQdlwr0aLCUsKjetvXF/LD9RL38Ynxin9X
vKdiRxFwDCh35q913ytYqfS3EnX/1IdoVaWnT9hLqDNQQ7+TwzI61sSqhlCyYQFVLPM3ZvVsTCq0
bZLp/KbZkNbws12crJ0BnzBHv3ih6f/QZUyA3xGURytUGMJXSOr4mD8MAMEO6nxO3/FdAgIGJ/sK
X7UiCmqif2+w0m/SjJ0rxtowFNIkpj0zUBLXyPg5T+J/Ekh9Y7UT50ySG1hSmTwSWFetEaKsm8i+
j4WCsFUNTs7FRciFaOAxx03XL9yZoPmizvygrFN0ch5JFvGeOF5ocBpr2lLYMTYh1/VfGP5KqmHc
hCe43V341Wbj9uVtDCQm1y5uXZlLvHFj8IhoSISaVwPaDDuLvWLJfZy9UwTT6q2/7y07IOkFoSy7
AJUTTu2HLaKQ1cyddPYBLKk+lF1yKyGWRdQtqpvEtf6WVC5HdT93mnwBBVHgVsZRfHp5Px3Ld7uK
ArHLbDvv//PZaG0ixNWgHaHudRAjyEssKZicTto8ADdaSKTsKUVbyYwDNQulRoPMPFaXCE/aeTSl
4CSUaAF/g+GEVrVVIRcdPNOXV1mstIXBs9km4WU4dAlc4EanyDzlzbcjyaApwahQbskGZ4zWoIwb
0UdNNNQSLfOUAF+GMl6w39UVWKLrarhWYHWnPJwmEdaUYAB3isZ+rwHspTCc9Opz/f217yIAjphd
WRoD1piPKDeagz+yJVxpW8ljkzTOz3W4+DnJ7zmxGNkvFA3v9gfyjdUwqe88u28tAn4k0hjAHCrd
/I37hrMi4dWRPXKWp+n11+yrWoP4iL+Ie0D3cwyW6gX2SFNjHLNWK/ju8dlLQYfOHs3yqHLCMmmZ
xEH23UbpQiqpBKdMpsige+PVoDOmFWnoyfDksHZIqtqAhwXA7zl4wJBZpqu5ol9C4aKKeenezLjs
yz8rwalI8fOXsrhqVdNOwWkbIMA15GHj5jnLNv8FlKg79Karj/JgBcnL/IUYZVi6yReaPw7DwAg+
QyW4LIXnbQFNNGPdp2ottasRne+5jSlA6nFHzxPcNA0wnKKFn8KeCexulYXw06QNdQi8dDWdlb1C
FvvoUJUFliBYoBu4tDPX7zllANmQGseRpUtdOSwRgS1XnNwmkxL8dq3PF7MxbQT3P150wHM34Sl9
Nrtlo2+HOKarTMaz7p/IPEIaxjBj0Wxlbhxn9v6dcGiBbGFVWLxR73OmtvGf8Nsm5w8TEhnGN4qA
+3IQyPaTiB8rmGF5lcJsv4b8/7BSjhxGkCCgVQvj05K0DkiaKZtymcZdbXjsK+Ragt78YU39Zchm
SKHzcdFBaoeF9BzLeuLXAKq56pHf380hBE8XYJ64BA25qB2oRZbwX5Jw925bTqqbcl0yiFOAH8T9
nwTAlqkhx4FDzk6C8gBtQUZMIZ7XzK20OBqrLlDeaJfVhzxGf3n9domO7h1JHiALALz+jfLbqZtL
YaxUvSIPxN5fILbm3hSqCWcKWK0UGkgojiOJ1Mdcq7xdEWaFL6OKVjfGlyq2JPQD3jilQkfdhABZ
PboOMxVpC+MPToDfXaLJodSeNkOREwb/n94FARsGvfkPm0TZqto7PPQ0A+QdSUzicsSInTGMQa1W
Zo0Jqjd/ow6ShuedkafeqtERb717+NUnoI5vFYPKI/sbAfLKtgT/VSCCUt/H6/vjYosKGVLrXM7j
Ke9J45/Flw6Gey6UskN50c8QcqJBP6ye83Baik1CNTMNti+lnGinyujnrePZSPixAn8Nei5h/DI1
0evsfUIooUiUFUYFOYKwJQ5kFkKRx4U0jsy4gTDhF9ON4cweGl5tHMGMYo7njALjqaSWCHhKtWio
eukA5qSO07rd1aVjgi0TdA8Ih0X8/YCWqGPerGi6T5nwKIXDGoHksjwqGG+U0EECw0gVubUVuUXo
KQSDFaBpRlCKGlLJjSxNtWL4D3qZPuMWBUt8AuDojOPyf1E9JpkCcxvb5dJKM2CYekJYK+F4XQQy
ccvjNDetv9z4UH23X9k2QF2KdCj4Z1G1HRuK+MQ4Zz8nsRMnW/NGXs+4bzyOOeVnCQ9sAioD3eO4
01wLaftlLcbskQ55FrQf2nQCrstxNYq+Gv3Hp5PqXYD9Z2abrSvad+JaPIjX14U8MMpqobNZM+i8
uO7DH2KDeZGFN9D5acNXh/1lqudAK+09vj5LKNJVhseams2qf5S/OD5ZVBzD+lSWGr7MlhE99gEe
jXnralxF/40Zepyl6qYr1WF6XstnPAwSlV37JBdi3Nspv0EM86zBWnzoUvSs1k9m+/ssvOo/7rCw
Gt0lErxdtjpHNcckCAoW9U0YvY45oClO7xweVS3Y8U+VuTW7ooFE/2CWnZzTmfTFm6KDt+Sh6SPW
UlbqEPJArwPbXgZZT4dUhFPXYLQj9KPQXuxSlhIWlSuyaxP9zchnzING6PrxPh0Svwu5S0BgYTKB
xpNDORK4E9qURHzTKg5yraIDjGGe4ZZ9pDA8PkEwZEY9Bdy8d66TdKb7+u1dqHVEJryaya8xT+up
0ScVNjbAVGlCfcnzmPoK1vxNblwuMIO4eApnGs0Ftfw4wYtG8wslxt3iEtRpAGSUO1Rw3JUM+NDZ
uQ6YPKvS1yygipprK2sTCEmuWdFZSyQXOXg7u4Ga92GPm9VF55RNowfCibSxgxjUjAIffbNgMBJR
Sm8Dv+s/Xc/bVdwOBXRsRwsx++9ePMbgOnaZM0mASHjBdjswWzNjZoffHAw78zkkxZK5swvvnbtL
UxG5OEH2UFdU3lAfaYbxk64+IgXSzUyZhSaVsG+H2mEMDq6uEAV6XflTM+vQ32BdB1RjN9QgR2CB
EHBLC5Dn6sYGLsZwmNM3Kf3lmTD3hRfafLZiljFpGfKmEtexqUNFvlMK8OWjnt4InJMUazcTPuz0
qo4jqX6JkvPa7+14XqQaM2wCb/hKqHMQxozqVuQyCfIQpoKpBpDSouxbwgBCjgl9IfHmN34jAwdv
P2eeibhFPlVQ+EQnW6FYQX9kG9c6R9DW9rUCW9TepTgK9KAOb4DpjHNiUGtkk3Cs3JrUHWJ46/pv
wYdBkVERrGVwgDqm4dWRbZwTUx0PUSNoM8uHRJinyAMdVaNltU5nte6A44IZvSz7VsbNnnPawdEw
AoZ3CIdZ+H343CbIcpUtMKO1mifPx/4RVo1z0xegXIQ7UmTbp3VL8R1tub6TWiycMWSs41FUlJly
WajKxLa5LW7aWqJFgeVN3LubcLzWsC5YM57MGHjuYofVZzi/GMK2QBGgp2z5dyOjSPTi2o3uatCu
NKQTZfXtcc33JHsgS614AEA+au3zXe29AlBYiuoiK+kzHoS+TJosvatMSNxOxww0/tsELEqJYPMb
xnoza4VNs5jJNG1qZ9KZGVaWDOHYt/+B7sA5QnJOn4/QkUx2cv0sM8tR0AQtpQBr9xw0Mt424LSb
7SnXsy8orLYQskF+Ok3SKRpJbf4OnEWPFgZgakgpj2xf1HTEARc27yYp/L59/bt4iZyccyCtfr+O
z4/wxIy9DRP4Lfd2qQiX9QCYWqEmYvBWN5y57JpKWOJzCwZeSIpY/LAuVuCoyrCmiBO7J759sToU
+/R60CkzyXL8WHn8GOO10wH522vNHSPIruyF2odTmlR02t/+ZM9PYx7lhN7M5iQV2Q3YNiDp/+wd
x9eQWoaTftZjBtQAVe9TGZ7nCxekpsVy2jcMBvtPlgZ9WDg1zeNzcK/addax1wp/vCF0giW5M0Qd
rrsjzcAPR4SeHww9j/PendpfeG/NNEWKpmUN7bijBR1P6Rjb1RKcA3LlzF40EqsgSLgWH/dgKQs4
nowJSt8zZ/xFWtX3Di2Or7SajchfG/F5QCaiNffPLgIA4v3JwOvln0n8sb2T2JZoyaeWM5tj5ARf
xdOTKrfs2869urhGsdYl1YK4M0wavoDH51AX+wUKV19aThY1xyGnGnK33n1uqBy1PFpjSlmloVJ9
6bxW8vVLFL/80AleNTzkJjYnrfYPDg0Lw4nKM3abC/Mxc5hquwzotsbEwMojHDjAN0vyFTlGiV4P
CRALd116u1+8XjElxuIMPKmzraiX9mVlWvmvdBpdbgX8YA74IISU1SQJ8+EHnO4dI/AWKhnQXvHu
kzxkJL99COnYDFu8YrUwPzaIJ8DxE5jmZ875ErIGRLnUs6KvApVbuMH6bl5PbneOHq/2LOXXgyA+
tAa/P6uR9V4FpyHSaV95CmdSkZqLDBdaM/BZexMM8ToLw3GjA2CNtUTEucgdV9yZMn2uePo0MUYc
3dKz8aG01z5wKh/M7VMOCOh1fO08ubMfTc2N5AhoEX8SZDOp6h2mkRPSSoueoGkWVDbKREvXiFFN
3hqT/5rjViUdy0MGWwc/NmGDgt55PGQYh+3VPFsdHWP8vlcPplZ4v+dn+RQzC3HgdwzshaV7bjCo
E43cbRiehggCAThrogE68shrCrA35znGaKPu5pYwwD0R4mLey6d9+XNmFcsgZ25AxIJC7D5XMty+
qfruw2jmctboUWlDk3/5NJMwAa68seL1iJqCNgcWMfe0Iv/ocpUKIhIhpk8rO0ThzKUCxBuqvb7e
t9i6RNzAXl41UkhtcAVpk0UycXLJZ98qOyw5INAitqKH9xoc+CUiyFD/uZgIXiubh/SV/275fzYG
NVarJsdesrY2kCWxj1ubudX1R6KRqFoZTz/c4IKDKRDCBIs6Yd83/dNbd4NyEIgDFMR5q39jvkk7
TGNIp3Qkt8dTQ7uwkX3qLOkHqJ/aOT4NpxGP4j7SKKEvXZNoSLPqMRCgp2EGPbiUdq1oLtC77XB2
KjyR/Y2VXfsN0VjU0Nmy84xp886jfzeDNxFFjJF+08BBjAnmhSc0WHPwl+a+Von9NF6HTKtWNUfA
PfqM/ljjIgm4HhkAICziAXahhJiaxfSUVjryQG604fH2qC1CdDKsLNZRobtP73fpuxY3L26JR2po
oUC2kbJBR9oiT4XS2bky+78Ktq/lr5fVEcS/hJxlw9Wr82TgEIFeWCgSW/YZf0p54Tjz+OibYmhf
C33OQYNjnh8GIxVh5OV4zPv7xYDITK8IRgiS2i7J0GyK950WBZL3vhgTfTdRbDCroKOb4lxzoFH/
HrAm1/sREsl8ViOa9qIAjyYoIz8uyzKTei9tfj26bFPBfWPh77H9kSb9f9qGAFSSmD+2nkw/vNoC
QPVI2MLzIqZcGch8AFZPzUzPEYxJDni5wgcuVxOL4n0MaM3GjMou3dpWC9boY9FmIUy1+ath/I4Q
Rtigo1y8P44OmdZN1sxI3D3ZDp1vy0U/3jTBDbYuSG6IcRzMdiiiYhL3cvP5Um0+ZBJHoGpsUC5a
6XdQTPSKsv8Tzo/9XGrQ599+ly4mEFgE2E0Tl/GPBSuN8koVlm18ST2OO88kxsRNYYwZ2t+BWzT4
w34eP/XNk2jJlZYWOMJxiff9H6hkSTBhQI/nHrG+xkAjxsYQQHaIJaYR4NCUs2ErFtLRuMguHMzB
q+vD2dYPewJir5YxCCyseN/e74jijP+zPUJTmzTBXZ/X6z24JTvJucZWnWjRmQ/MyNAtjze+nNJu
93T4ldfSC/2JXHDsvR07E6lqOd2Q/sfU29eLCsG0uy0J8PtUBkg/Fl3sFCkefdE38bF2wL/VShTq
L9vqn1EXTg3mQU7QZviOIGyfzxIdFCrWNkGUa45PYs03qIgNGbOFu9tRAvzkv1ppFEXPerefXFY+
v22OICHX02hrT2ldD4H9QiIZtCM9NVCRtr4BcJAphk2ek1CtgM+sLTNw6sw3NuplnbLMhWD2BzIh
4XHqtv+cAgJ8LXMgpZ3YZEfC+oqQHOHB4IJr24/v4Xo6TYiMMs6TSTppPeK0+s5NSBbAFRXwelpi
Ab7qZBeJ4hutOPyJxOs24xrt59spZDpFz+dVHb5XlQYLvAKivOzgVexZoeb4wu82ms9hw6Wo8hfZ
dL/g9lKxeLSDqSOq5N2JYQ9az8gCpQWbWcD+dBhEjFDVyIZ5YHF8g7BRgRZzIBlgyaEqgGpRL7U7
t0YdpoMUR+xCYdnlmxV+xhofpHHLxxA9ra0ulQhtVzChbQ0mFT0rce8m4fRZAgT6GuPANwXCJ36Y
hMRNUN5FHo2tBFo189L+HFESIZymLwri7sr+oM/I2/ma3pNOFzUJIw3yzLqnMc2naglyLRi8r5QP
e4u5VQOJ3AhrDDDVHU3SDtevA6ckNE+fM9MRGnwfrYxQIG2gqfaUMaL4VkWXHF4BUNLg/MusO1JM
fcYsPSw/v2RaQeD9QQkuYJHx/d4IeFNR4sYZljv1sTscWQCom7ZESI6dEQS2WHQPiK10PiJz4ToH
I2XjSMieevcXVNxa2VfDewvCMfPq+65b+ssvE1mtZ211sk8FxOsy5I1nIU91n8rPLrc21neTupeW
zeAJp2/LUODSVqX3c5bujGmkKFSwCa3j716/4rR0t/L3Z9stR2EQ/Oc1mM1AkSokd/UIuxYj91m0
ssk0vFIlWQeB0InNORTLLEnd3nJ2Ic51qldp+gSLngPi7qwNtVUkAxAgsna+ARfNMSio7PJyl5mr
QjOJ08AXxnwi8Jzjh4H0mZx5ze/HFk787ZyXnluz4H/Oz7wzCkJNEXnXFer0NGq5PbcqFTYPW76o
M6556SvKneN4oh5EoJnNOxVneGq14KHX014r7e1sJPwLYWjLQTlQGhemV/lujSfh8W5Pe+l0S7Ry
3jDFl2g290n8gIPtsdlepj4DHGFbFiDt8SFAznv7g4RiN1VZx43K0dRuRtC6GJtTQhbp1B4s7KY3
6WPPDH6RMA/xrOrfj5tZsGlkiqKHBVpUb3YFBGMIkZLvDTHTz9jU6RoXneTt9czA1k0kc2QGuRwn
Cg1/NkeErZKRjF+kiXY848YqiL6TQGUzp7T0hFZq+WG6bH7DliagMWqlcI5d9385T7mnQ0dasDrA
vPEmjjQqitUpV62uz/1WglpB6cNLtyTey2OcKbUV7oo6GgjRuds91AoEoLaogcALBe1mRXBY9/KK
vu+It5otrgitjuGYt21ZMfWwY1qjGNbglJq48P/sP2/lhNHItpYe7R9F1Ds/4oK2h3WS76VT6u1n
qQx2SyLgCtzqgh592wiQgwTly7TVTKQui6hvNj3JIZYpsc0uV7kpDr0s/SwRcwuzAGgLncYu/gEF
FUVbET9D/bLYIkLRmQiffMrLjbCbdk/4+TXnarToSNRx5FMT1W9NGzqvNA+5NOr9TxFXTo+Ul7AH
6XJ8DCNm3pZ+AbNFvv4oA9uBd6T8eJseuradm4GiT5yICd15G6zVm66JTYe4LaBObcffKx1H90Z9
sPA514FGkWYTCC9eUYs4qFikZlImmY1CijczqkGQqyiIG5TcG7RpLqTfQU21ffQy28AT530rr+7l
Or/Koeh9nbWglMQtmlD1zqFzev40Bo14l6OJaSY88nqMGVo4qPnx2czjH0w76ZnIRNRducymd5KX
sjcWJSH98uzkgKDJFVl3XygFqZ6Xcr8YZFAaXyBBZqI15E6mG5IvSocD7FWBcM9hOzM0V3P0oc7v
UeraYhjeU9ie/qCByebHe+Uf/eNif/n+xelQh6pIxsVgNXevJKDZfiP3inIZcarzeAtGJ7nsZOgj
8WuBiWBpx8NFjfZ4I9Z7sQa1XZ+WULtJNly4iVYnJRhYtBXBjJ3BcaHsppEp74FHwaEf6q/GYa/f
ARgXvBwlAQlTtdhr//pkaZW8hhBVYnizv0RA07c66xIqof1loSgXRqCwc2q7a+gmCIyaQUu3rFPb
imBRTX18jZ/mr1Cg4Pd7yNVQq1W4zaY1Q+Hco4tYglVktUJsYjTByUgYlxL4WMQdjfwbuDbxZ2uI
vJo7dZMNgPI3F3MLMouRaa0HtKKSjzafnoJF9CTQ/KBsGk0i4DA0mNN2YcBWVvkI4O9SNeYcIMN1
vTv7z42EZBQ7U98S6UPkthr5/nfIu91s98Tm8v7qs0GLDq3eBbSkdHq17MOL1v7uze0uRXf+zPJb
KSYLrFzyjkDBumBP+7/DIlVfaTUHBLZgXJhNBF0DMtOVs/WF4q/lmijCtOsWh6IXAlgTGNaZbOPq
xqS+7B2JynbpXrizERGtHNRDH+Omu2B3BsQplyP6GfBmcbT/omaqtpPjk1xJ6qerQPWxlIMIw/xU
zZ+Yy3h3RQxXD4ypwrwZiF92vf8hpv4ai0qpouB3n2zcHvunKQQBET2MWMRGMS9s1l5CLW3HsXPn
kmkzgS2dt9GSghndVrA1gE/NkuN8v99a/tVbNjSkSQFb7V9WuhihCj7I8S3cgoVab/Nx76fTAqGj
OQm5Hmn0i+FcI21phHaH6l2vyaR05FSZMlOIXUOWQNh7TmXBJMpEXM3BnAnOIppE0ldWSu6oUGn7
9r8RsNcNyB7MDzhlKP4GK0zY+WjYIuk7NRArkthBVWAN3LZLdix9aVMk4DKH85hjwSfr2Ny6K3nF
32B3Y3AX2JVsqGjdyvWUaT7WdO9wIsVXa7jS04Tu+DyAhLgwJJCCJJt27gG+YpmLhL4Iiwf5BEdV
mgkimpyjDdzxRg2s7CqsMQeaM/b7N3lOoF0ZorfGG/kWeQ3RoKlJwuieoSN9xxI/MJvsP5d/s5pj
sWBBkw0gu3mL2n4nIf6bXmaGRS0Dp6Fsc464J3PknfvbZW/jlcrW6KzoG8y0G0jnP2hweASdsii/
IeSePW/ljbFCk23DTt39+Ca4r4lPjSc7a/7pIqlnkNxEgRZzuUIgI9f7B7WVbWey9bqQRfpHQ/Ey
dYNWRnGQGi63tZL5ZSrm7TM0jlwbX5Bvd6iA12/Csq//3Y9n/xxF5nAteHVQYwZQaHuxt+I5D+Nh
jBKRrRBA0hPRnsa8MscmY/Az0g0G4+6CBldFUh2fDRFBXdymeQ3Fn2BjHyERKN9GUq86pEoVOfOR
989jnZ4juHaeOVuzUaO3AV8gdl5Jk56xb0KcZ1LP4OAGoOGKFOZRm2iSMmmMjTJTq2M1WhxEq1m0
FLzvQWXIf3xFvt1xTrT0uJwxp6Jv4xjVPhpeI9S09sf/0PCFea1pWrnXStge/+No64xhhVmvLfgN
4mP9JF+rGqcqOazL/3lPTgrSlLEDW1k2uR4fPoNgdp/UPFPcUtcLrYdakzzqmm2XWiR1r99FR159
A/zVkJRS7Jna37Uw+wFCGcVhhML/S2dLmYFQbtAtO3o86pvjeR1NRB2dSEvLSR2yNid5Zucc1Pb6
MaIfL9RU+5bGeLp4CRtj0z97fTEcMTByODVpPLvNzIv62+ca+q+hmACJNAUq1psoJvUWQe83MaMb
GlRDmV9ufI09PkecC0+sVXnhWjQTpW62aWiOKQtrQ45lQoV23q/tP8YHsluoHUg7TQ2CBjJ8OLwx
YQUNWJYLp8kEw2R90YzZB6jwoc0xN6glQe9is9jMuG47Z37NkzuorWz2W+Gfg54ucQOz4zVNBx5K
AEnQViPLkLU08HjlEu6lDhLcw4C3UJJEysk9Hf8a8PaILpIhvVCPk8P8KFY+anjiD5CtSikI1Aco
jTLATHUq5zJSSpU9mHrZbKts4RfiO9VbxBLwns86SwBPBP5CKFBmQt1spxWkr7Wljz7PILJ+qj3k
bU0galKrM+AlptpwQTTh23oGTvvfTCwjgEWkyGBJNHZEsxoiyoQAW7i0z5wgQB9J97e38jTZf179
ZLSNiKVY/8yaxoc+bu32C3gdKRj9dfWwY2qa5S0aNlmwUKu6TIuI//ug19723AYMdmPQtVwD/cUb
S64ODLsxHOM262OWAFE5zEVWQAxd43HZokdL+Cn0vEiS13ArZ1PwIWqdFOf39dlLXit/S0MdEhEs
R79QjlR/1r33lJg93OJlHZjDbKKoBoZVn55ljb2Key9wc/7gzdxL7bQSpH7Zqc0HpJ8JfXzLHHCI
BouZ+NcoCJmeEb5a4xzsq5iA26/hL6LgurM5sp8SYAr+Sp5NLzgO4Q9drIbOxq4BeSPIdxce2OBg
6FTEEBdaxqYO3idTLD1ls4Bf5lOedq9WXwGI/P5ESovY2GybvlzaR12/zOddM5ZHsRliHmCP1OPj
lL34DasHyKSC3Gq8tDUetJnN3wYpkzM9YaNQ/B7EoIi1+Ofnf732KnXUwikZ92Wu1SEx8aYSuZUU
BV58iGSu6yc6QSy8uUBQgYIo6OAVxkt6uvv+e1UiFcsxhmxh+lQ3Vw8i/KJhkzQHZJifap/qA9Yd
ckNkyBrcgki8PXWnrD99yykPhAZ0O40rLTU9VuYSiOg1BiJs6K+nrK3SWL5kTGc/zTmcbx7cV83/
s85biwoYLtSP2lF+i7diGC7vKHgzTYOh2dsc7iwtsK0SbbcqSlmCZXhn0K6PXNkki9l0wVl9MGb4
Fo5uxowhHdAZAJrweOj23PCGYl71THmeesrInn2kGQ4iigzquuZTqBuiEBNJ0Ciy+H5Hr03hkRUA
BPyllt4TK4LL66sZpO/ozdlgXVFrfHGeqqze/c2oUDE/YZbf08ZLCpQQM5FU0741GW5+VenrFH8m
AFbMn1EjS5uIc3PHoxmdCs29FXGB4M6XGVMCOl3DR/XMMopf+LQRPuvp5kUiyPSljraBgqS6+a08
9XDKfGwPyowL8LJTh+IKJvT5SeWEyG8zNrPCKzZWj7pd0sftsK6M7RWvwjMB08PNVphHgimnmdlu
vv3/jWvXavalLp/S++WTWqRddpiRL8/OGL5POcpllzwzFJ66zQyKjamTd9hgUV1UcaEyQpvM3n7S
TIav7dYn3p5bGBKD30+cewE/ZNZb24zlAvhQaWtSyQhzKsB0xvxxVkbjoJ5VE5DFECXaNNadtgtj
keMMMRUsPYzTGAPReu5fjZhOOWB17XZk05t/LAJ5y36TgWOnMOjtv0aM/3ORymcywPbMTjSl5VhQ
TJJ+pbIze3NZ+e861VKFlPcqOUYfkGTkhxv0BcJ1zu98AjWhd4PagE3dW69AiWtWujwv3p1aqZuC
2WwYngqzjVky48e81OjzdvXGHr2+MSgfAAcFKSyUHZrmZep2Vqbio4Zvpf9Jtd/xcVuyYTLJHHYQ
UJBpa5o3fRGdCxozVjOHjlePVZkHezhWVu4ck0QeCJZuCuCQjCYTBmlriIioRxNME2J2QIrcgE0o
JWFTe5tyXsiYDHNspyHC3cZS2cfWQtyITbnP4xnw7A7NYaIEHA4cqkpnbzo/Uu2DfcFimbYE/Cm4
rgQ7wSycwYQXMZI9MVoC50CxzdUjC4UojlXkhgX8YXXbiBs79KdYYfO/pKdGRgah0oJWDkr76bDI
IK8LdmzFeiFUnZaNkdGO2DHfFQrEZoI2/FzYRp0hFHmlvfEQ9wobBBBLwd2MatZ2ZY/wIpAKg0Yz
jOQPWi7k0N289p96dAUpGivW/PHw8i6hpev2tU8gV/NTdfW6Qv8Eh4oAYIJukwtZasE8TSAHeI0l
wgTAxZgaBetTllLHzSSxZxrXumLgFFZH0JnBqP44CeuHCpclnKEU1d0/0MqBlW8SDR+2Tbg8/hUU
DsZKTFWcTRRCuMi5CXwZCusjUV7BUj8xnY2o0wg6kWNMiXTEzv90fG24JKhoXI+SGK+4TgpAv53K
DQEtcbtr+/6chHDajbn7T86E2+8NHTOcvLoatijlrdcYsv0uxNR5aZDlCKYcK6Ef1lrsZSKhLUF2
OxYWpDRwba1HiUIe2YByKljySyfqAQyE1tGFPaD0UUQD2oJUlDZiCyIZsOn0pfdgtgXixRO5c9Uq
A4kGTtU9SDK0srODYUPy113pPNYCbRSx3anxxbw7nhD4ZQRo+ykAAqiohTHYj2d95lJEuvFs2G3B
BKEUGPqlRVhfKlUXs0NaxdnoNl80OZiYNVQKDnImxQgQ/U6XP25Q36pQGQadbqrKFGugTKfHrjq1
lCpdAl/OFyRY+l4/csRKdVIjgzDv8zIA4x61AjFHdhDP0vn105/c77UCBhC+trQmrlpeNQu2vjBQ
eV52E3P3+DZDxjVKGuWoI/0RTiK6+iDbR1oSxZNcYEAUmeEU60iZFj4BrAIEZ2XlE8GzcQcWCTDS
BMAJGQyG1Z25YPjDIDBp/Fg0A68ACbm1KpjjxuJGUREGYy7dZfu6hy422R/Ex2QbLz/s6aJgoI6y
UXBqefvnha76ydctqCrLAcGda3VEM2Cr9XxGvADogMiv6Mha1mmi48YDBiuuhHjzCJzUzKJ9zkh0
O4WT5bURjRwezfMUozr1OfUa3/a+UWkhZjBzUNAcD41xpGUyj2JZjAUXOHQnTGZN7ho/0uKOVViW
SZAeDNuegLbSWEf0Q6ciYkeq/SL6ricL+Nz9wI0zj702hMbv6NGMw+SYAU/fYmB1bolN01/uOq1I
2UqM4fUZw+X/PagHeYXLNM0wVxWfCs/BXfw0U+ZgWTXd5tPM/vSZteDAaWYJeMjj9zWn3sRFSO+t
+Ia+FyhELJqcjOpFDfJIuc2wrRx3GyybL31+rG+9NTQX/leUzO8Ppjeiuo7PhcG+URge0EwbVvsH
B5UyDuNxFtQqlCg/NZay1MPpr2wTWm055S+YJZ7x8MmvVtyxgAfnNf8TGbAAyBeW65wfLcyvAuaR
lRIdbkgB3prgFEwSbIkXFFatHNfBxgK4hBdVhTgrjuG14OAkmHWV0zV36qTd3+Vvb581iWGGw5G0
3qWMkRQuicM+aDs0ywPNR0VQds9emikbqWrn/Qg76aPuDTvWlfx9DwKyOx/ztHiXfteeWlDGzGaE
eR5Hs81z1IIOBv7VYmzN2a4S3MXWChVQZFahQTd4C+gOu37Ku9esddlEszhlqr0dycSDAVHAHHuD
kXE4PY2iti/OW1A4F1IyVJN1JetcfAWKRBQezwbwt+5lNUTuP0p1bdeDbUjRVdvIEjbiksSOApdw
m8XbEMCV649HIw4W4S4M6Fg3jESHsC7MSbxzLHCX6JPfEAC62fyFDdVVVkO2Z5FkPTx5TBxVt3PS
DhwioqPLJm/hpe+E7+1Ev6Kq7EZSwUr8DddGe9Wu0ZcY/ivCWfehPE/P7vUqR6hR44ENxcbRvzHK
f06UAEp7Limkel8pIPVp6MJIbjrekLEyMFw8AQALPApjtZf4Z6czhsUHHYp3kXx+FhYfuOGsUMhb
ghQwiy/UPO6E/Dfk3qiCou5rj7pSCpV9ngHBMitMSGyuAwNMZd1GwQHieDZE41yiIUg3VDNSiOaJ
+6kwLVd6H5OY03cSBcQ9as30UjoSu3SqpXeP1OSHt7/JMBCDTg/DtgdfccpoGkcMbFz38NKrdL0q
YWKW2AG/DRi0wkRDT/5+EM9FN1FaoxngQGZFoWQfdr1dfl74RuvTeJ8Lz0Zp9CwAHMttXH9iOk3S
6bVS8Z+lyJsf+f+dB/tggIydRuyP5i2ihl497AT6eXZBT1f4dmjRVz57G2+diivdqAy9TrGxi8eq
ZMBuotYuyXQxuIifE5zgzzYvU7a8Uy3AqFL7rQj4lmazHXZNOV3zQVJg+6wzuzwAyWBLIts7/EMc
El+0Aj466HFD04OINMNyBf30EyIyNUalxhSPKPT5DPvKSc1wwiry3Tdtaak4tK4qGq7efKc5saUO
mbCDIkoqeU1afe7+ZxaIqSmSDM6FPcVG0JPzps/PtYjouR48szzTSXJJFYvagSqIw96CFccO/w+T
Fd6yzxFz150gTu64XCwN0tEZoe+5DFl3Pxh1DOwVDMGlZPb/iVSebh78wIi7mP0wlgIsXh4dCBcw
0qK71xXh4V0/xuwSfzWL6x2fhfcIGbybkQ4RyzByRjdHlDOOVsrkTK6vF80iWWpPIWb6C30gNXWG
cygqKOxUkJlXCrd0y3c3qfcdHpfiC4UcnvUpfrPqBe1eYe67X9jiOAq9e6ApynsIhmCOMXaumWsi
buzcNJEN8ez3LrAnOBT67cdQMVZkSbfs7PjB3va1+gdsIm3p7HccbLGRxCTQgF0hGyG27XlE8e+m
JzEmSIQNS33zBfcAoAhWgLnXObIY5hum2z35AisFefQg7O7WzNnNLvIkUY7LEQG0aFcTgv+INavu
hKsDW11hbl8yIaZGadYw4ivC4hembhj2kHLPENIr1n0mp4u91Kt3KSCo2dzV/IQCY9Q0dRHVJH6G
dEuYGpKCD50p4LTGWMCgVguE9ec10h1r+CZfhRrpp0waLk2eFYoHApYVEofAxgeI3CzJ7ZpQ7qIy
+FZiKyKqFu3IMcEnoIvhl2oMr5uPVpNqUJsjCWtewCaNZRi+KqiaXrz7KX2RFCww7/2ScIZj13GM
Riwjipq9UBLArJ3viGN+7UjnOGTPc4DyOp18tb19etlyv9yL9BGCdJ2u/OnPo/tGeoUCFIO1XAg+
1c3ND8HDYvIi8iKP2vyJmTEpnPQ7pAFa66AM3+qltYQyvmN44gV+WyKIH8HFDE3iRt0Mj1CHNLyP
y94pusDbkwcR52Cx+lF8hESB8Lkwfioer306qfmtygpIUs+7Y5PtvXS20gBdUCITOZ0rEQ9wWwoC
+pQM00SyPi6smGbX9UfCP1hwyhscLyTzL9GiteSERtJRtt3zCCJYKHe1HL3PlZURljP5x12tZC65
98oRJKXnbzECe/D/fCMAOzekgwrMxCIZzs6VfpeVz/vitLgN23khTpw8/uD7OkTgj3iC9lcrWXWJ
Dv6aeNp2VAllT/6IG8daK+fA2GadCXAy7tbzokxdGlWMJKYIPq28LDzKNIdHy888FXXm7lPXsaR5
BwsLm9i1vPojO538KBPLM7oqi1ecpPuNPFOhjbSf/kzUVnd8LfnBdz5U/8LXR94o4JCXz29OHM8R
Vv65uQHvpet1kEZJZQpOfNlxhZKL6ZYrX/ivVot40yfNrvqWCnuRgyK8RAZabNQFhYok3Du8G8aI
U8ZF90ufJU0DDjjysytCw1q7SJEdhRPDvsapsKU9s61pPnc9FrlgX42ACuZyFu499vqEyzATJL+m
G4ljqalJ5MEv9dbKkq16MNWYjgAeGtT1xW8AJ+xj0kNFo3JBTdroB0Ux/o5Uz/JvxCs3BAGoBeU3
nWvsJPIzIFdENhTSpX0R943hp6VMTcy+f5tnFrx8G/mC+jaNdHoqR9TO5lohPNw1uIE7cDavuZnk
JnQghJ1ykwc1/hK8yZ87cCaEYMy14OYwmXJf7f93KYzoqvjeNuylN7bdxstttO4MIj/CyvH9W2a6
aPV9ATmW2RC6s02POxOEGfjk7oXWsqmTgWe0ZpovLo0Bk51zbbAZ99+ZIHt/FNSJMd4fxr+PdLa3
543oxgvov4bBOTvdyFnUZ6jug+bXXAcdLAWnWklvofwn4uParcfVFS3js0Xi0MSwFCXCo+hefqd3
jDfeJspNT0sNBBqqGzrPar9VN83qVzecHTbg30VIXnJL7jVOnq3UmxhrV5iO1Rru/iY6G8KgA5bH
qmvle8gwJN53Hi9LtrPaTTDnL82PhjmSyPqtRsavymHplh5D+yAyoCLehnJCwWVUoNgml5NhZM8W
5fSEPvWBV90Tq6y/xQGxHcyc8sALfeVuprNb73DhFBYVymy4ycmQ1D4woTxlA7gN+FKQUGM+vz7/
C9HbjTKr0Dnt9/WN/eYNYgu+Vk0hfdRuIUc+o4/9oK8SJEJXN83VY4GLzhoHSXk/KcC4FbFsZokw
Zjva8AyIjTO3/pa4QvAxpSKT2lYFJr/iE9sKvO5a3gPd+DBTEU8sqvGB+wEIGD1sLg3P71Vg88Va
0eB5Ksg5nlbPzgnN4kwEuwlKJvfYlD2qc99fkpCZ8UpfuQPT2ZYojEGbl3ZETVUaN3eHrdtwVt5R
idVydYnWJLyMEVFlxlvIjNI5vJn1v46ecjwGEtmgZjGHd5dqZ7O+0w58PPeKrUwgMPpDQKbjpNK2
5krkAbkJi9Iy+zoN9JIZplod08PrTeKylZLVI5baFUEi2Gah+lJkBPJdVvH2T0tmJ1Q1tCL3WCnm
yMMTuklSgo27zJG5yV7w/uLLcdIFD7B3W2xN5H5MVb3bjx9CCtkE86wW5m6ZExWtIm3znMrsCjiT
JxMUIa/ZDu7IwR0VE+FTEheywprPp4Tw8+xXBgrLHQq53WM7uU3zv+UWowYn2uIuxaKGUjxYazky
5fni0qLKsJJ9ITz8mm5CbJloXDLM0KLx6eLt/OchtTgPjl3bOZoLT6U5/70pEXgO7KRiT8llpV9D
7ZUzEqgRh2fheDuYRKPU234TRRhIi03yUNH+XfodKifhLoyc/NS7wWZuQlxxSoGbzAMOEDXd4KWU
zYzpUaiMNubQFB18DfQIUUxWYXCCtwh+pxvJCPZhWhF2Ha8JwY2frzxWtxDbjija316K+crFvIgw
TRicrq/CxMrEhv0Wu+zuSlaovk7T5P6W2YEp66jRiS1q5oD/nc2ILS159c884HpjaDjo8DSl9ccG
hFknG58SYkT9BTwtwLXMbI2oYW1KXfRVxbs6C6cXR/yyRDyU8DjFweBwENyOFUh9IUAiHfJZdCeR
e6FyTg0H7VKEwZvsxDV+TZHZyf77mCDk6Q2PYLIC3N59qBaIF+kl+MU6EiKfXZoDqO0rKJJkXp4K
3YTflrgYL9N+CThBLdhY/VP4De1OqvaevdBHzRqD6FONKdMAdUp2L0d2O3xUyvhIOx771cFVHIyZ
m04B2OvVVhyo2+HhxtxrC3/aN3esSHPsnrBZru0JTz9hj9cPSozuyBFCzKcra4ooWxIOF6PM9+fS
eK4Sx1ldX9byp8jSu/cA6QZw+igbLdTToseYFnpIEsE7rd2bqC2WTu+M4M8ZYdcaL/rgSFVJ2KgB
sYmSax6eHNx4KbFBv6CFij8qbF8IbXy6LVhJnbDq7764u3XugFk1Zv4sMPZdD5j3rOVlw9dRYLCU
cLEpOD8fz3dexQ8wF4S2RzCn4GC8rPQnsQHdaQ1EVu8v5y9a9ccvyXeQcThbt2MLunYV14+Kb8Hm
doKAZQpVP+OQs8o8oa0nEdI0rbSQLdjyo4TOoAk/u82yOypRki3fi6OAi/YGQRr0TelHo5LJufsz
KRSDPyyVjebCCC8YAx+SowzStJzM96trh/9lbluILTzm5o3X80Uo7S88S3yBqEG+oqFStF8inhQf
p6GeDgFaqrQNwjDEvs/JSw7sNuT4Hcjwfp2G1B5SpOZEnXgcFOgHKvz566i8Bv0aO714+MJlSP9s
0Wdr0KMwdEcirmBq4soEBBRPyOyw2fi0Gt2fVpfGcGuwDsF2c6i2OEUfoT4cbAbPX2FqsIyhvKXT
fijA0pwg0fDTKNkENKS/CX7uNbnM1pFJhZ54Q8iFwwFWHv4hsjbO/k7qGq7QSxYPJ7cMt275ro6L
Xs8WKMQEDi66LaC5vQf/myISwksYVyvzBKGuT82mSXtrvVEP9YhIqMTrcQTHPDM5cCUz1sFq+j2/
Uk/yNyvrafSkXKWaJz7Vspw8AAO7DNB/AEdcmfAaMPrLAbfF6wICgzWUSrtZ2gA4rn+kCwPMAS5A
e758RKglxyrUa7KEXibsJLqapu+pgWLFNN5sO4cIpNVh9F69qCirWEmM1A6lhi3waXe3zZzYIsJT
BOF8Wzl9P7VU5YwDt7um1JWc7fJS/Mo6shR8OkVhUw1a98yfne6mfCiV3U9Lmp59H5NYYjJ9iFW3
DIkmPQgWr3qFU+Ctk5JJchyKvD+7cM3BALOoJMzpkss51Sfz2xkfkSiXojCu3ssdCWQknIHogBoP
a4x2+8LHPQZKgJNy0AXgGu4WpaLQWBaS4s/JUz4GKcyUDsAvwPORX/QWY1piJ8cRRXBNJNQFvEO8
unJXUlIPmz8SpRYjLOqXGoqYBrfeTpCnVIMxY5VQdZKpHwct7mHIHxI58rESJyzyCoU6Ka9DeHCW
QVH2P75s71tW5t+eFKxIzvx3oRD74PW9jfB08CieqjFuZR5NtlfMISqKVRZJnscIkVWZtzOOCt+C
PPJXscO7FnGTjxTrYgYfKTpnp+6kFhAQX7pmLJAwW/2JReCxpfjZMxOLlHb4zYXRFlg8Hr44xv2T
BTRaYvd8s2sd9lO1bqg/lUUPBWUwO0edM9UUVUhJ3gUvEPGNcDjiHE4/MFWmr5ZFECCSHT9uScuR
HDbpEkgD+BWK4V7slLovgcKIP2C48wwPiseR+76wgZRztd8q1NMd6loK8X6yJS2g1+nFwZKyWOvJ
qxEEeUr/313jcfptVrImvw4MX69Iayk0KKJYSy0BqU4tQKTT7Hcftes7j7/pSdx7lZTWbb1i4Qch
2FlOJWx2k3TTLVwYzk8jETRhw3YZB8Pi5B00C8PcL97rtvSQzYxI++CzukVz8FRPxlicflDxTG9C
FDkBR4fZrvLCBe1+gHySk8ZIlzfDtPo5WG+/rDsHR82AsvEKYTShyQlPMuKB+2q4w9SUw56eNcew
dVjH5XfKfuACROrDRibHOw4YaFcxl/mXVlBbfFxg0GBSyB1tDQf6BxgHFFFpn4zTvpDRD3NIVNtw
1A5viR0bje5CmzWyj0GtrUz6GEaoU37ubPd1ZGlet3iF7umkn3r9ELq9JLbdWx+Wi98hOJBhNJZM
D9BE31RcGgLd07yIcmQ+rO68hU/RdPwKlAii6wvfBQcINCFhpuwB2vUUZ7M8dEPDrlwHqA7yTux9
xgMMwqq4+sHELteMG9yOKQGrv48V/TQZ+as1Iw67UX3CyRNSLbwzZIoik2obO8AnJutVw5qS3WI3
rwtXrecYvsSsOoY4/fI5vHGmqAbFktyHk0dgrAOIpiivRBYvY+jkWwLqBmHbmXcYQsH/WR/SJP2n
qpWk8mnMCybVosvDZibnMKot1vE3LvoM7gGTPIhrnpE98b3NPVvIydbteoz9MKHWYQa5FjNL88/D
ErDaifCrnUk+Vr3CjL+TVjdsdw42qMRj7kE8/wcxDdHDj8FqEnJd2iGGhx7wK5gCBA+F3qmrQyRd
lqbPt15cjYQs+sX5gzdO3767f/V65cmp7k8UbAqGwv9rgs1K74g6a0nboWyjWUUJ1CU4COYxT5nS
G9CXikxh/8ewge3AHyzLwwMhBo2HLcAxl0AdqeY6s6SMbEvWhoqt6mljiyPKPQbNdyYFQD5PKP+a
99B7Kvp/Xeb6TzBkVqxvDc7/xkKweW+iKvsCxNXBqe7MyljtwqLLu00xAYc6JHXQrwgxq+ISjdhB
dWD0+BlGwHmRkEWSmr5ZkJ/Onqk9Du1YGUfb23vPvLc8fB5eESpaKoQzyn1vak8IyAaCM2bOXdT+
qgHr7iEWZDp2JErr2FI2tns3FrQHxHviIb7Bbdhx0JGMMAaJKQ7b8CxdW6fzqmJtIhkBcFVmm8Ib
osanoLH7KVlnrQ4/zRdGnSxLNvOSaodfmZU1zqyidga1NxFvnxVNtxdj96RWOVK5acxh8X6jLFZR
nPm2eAuHey+FNJCKXSVShMAqfsrlK84hvmKIKydnzgkIDJtBTUeryRYDZUfdL7XZtFSCc8s9yISV
1tFNiPMr1JnxMLDQnSuudt0btCPAtVB1/TNAwEpbRaJb1LKtPtn8t+6XJpSqwL8+ABmaG1oF408l
Mo9jwvPMglqb51Wa4IxYESwuW5yaqUCWPaZVx1xdc9UBFEygY+5zXFQed9KB5tKGXFG2cENkauPo
OnigueHSu5/3dvIYU7oha66IqbyyxUDO63xXjIIa08nB8QCRBC7xfMIH2nMmMhQg4ksTULYLs2pf
d71NOFtMARSdFMQnmzCufeIz9HW412VnfhsQ9SRp88lGfbFIJY9nahHio2eOpYH0dGJ1IvBgMAjg
UC4I6g63mysRykyFy0D+NsrdBnvanz7On69eslFg0kfF1+571D27AqTTNW0RytkT+obFNfW+piZ5
VOuZiCHuWIwhUuyYUZtSY+qnXV/iQhlndop7Shfx8DmT+ykA5zx+rbGZm7ksgm7p/sab4hvEHeIN
rf3xZcoiIejUK8NFNavZk7cFuxNqj/rYbGywNi9XwEFr8xf6du2DjPneo7s6a7i/DCdBBtu1uC44
9gkx8eSGAWsV2Ul1F6ieYyQxIxjEEulOrRXmJgMKGNFJxQVrEU8j7QcRJ7ZU4idbpdAlBc2E4lp1
9u0lAczmnm9xpRVMSx0Zjagt1SqO+tgeOyR4BJ0nXP93lC/zMZYZKWMhuVD5fP132dcBPjd99L/k
FWK/QC4dK+rmLoSLmGcKOYiyDZfUcvq+E95+LT33zEy6AbWd/IwM++uVHI/XjLEyPQNokopvuK58
PafIgpi/KU81J69pO5950JhqfCzW7dNNssYZFCXrx2UuWYbyoq1xn44ag5N8Iaf7nsRpUyMoWkpR
ay3seqV2ue+sIj1J8kJjbNUAhog4rvcSIms00MnIJq2c8a92+tXEJd4JsuOZJ+6GvL0mazCdNTNd
639HKkI02e1wible3RAV7gHDcFBE+BA6XGY0Pjml/gbGBbs7SwKiYXeHkkUaoEJzN3tGK6bWPzo4
h/CZ2wuzYJn9G+F7JwYJFdMlTgd+mzciH0jtAKpvLzreZT4lSBAOefV1a/eDBjvm7H2jajZnebzu
sC8snLF3nCZ0Xc698pp9DMnAC9690dpgIs5F1Uk6ATTXmgPF3xJUjhu1BquA11VoV5Sl86U0cVBx
9y6+mecOhU1YJkU1f2y3iTIjvIpFJyb2EZ6hvRMtRmgmExc5MdcPLb97PqFAtNNp6Rp6CHxUlVHx
YhDy/Q5n2GcnXPXmVm8D3MCJvwkWjXF1mdqMIsRYPPzzCa+Mhp5IiqmDL/pKAvVCqUm61lzmBfe9
Z8AbJx/txTy2UB5XrCfgb7tddxu4JxbHBZ0oqWaz+9j6GAkRWD+YkV0oKRK00B3esVMVullaU6Ts
DYBil3QCEIHUP0kUssJhBiVaQiPdt1SFC652yTWZDCH3w71yObbLEeFN6fTRX76BXONzwT8q6hFf
vWcH603FchSH2Me1aU85kkKyrJZ5tBfdjEIbzq4OTO5dVUyxXaVo/TJ0HOP5OqIiPYlw9X+Fy23L
GdazyBkxQPgWi7ckm2CVZl8eesQds14xKT4nS41OZ3OcR0V8GpXnj1uoo1fOcE+wIg0IGerC0yHz
0FUA8QZc9vZ9hjY5oi2f/guugD3RX3cYdSnJ5nmCTWiCPTRPZC2zNYeGvihZNtuTNY7myfuzRvdP
VjDZWaVb2a6W7FefxJoTPBHKGZYr6vmSMtCY/Kj+WkWNWY3fpQ+rdg9ztHeYtc56Pw08h9U3HBiM
hYDfn9NmOJ4h6sDyyVJJAOoYyC9CbBnFVWEQywCouyLHfCDwAEg/NQhqUDkEFXlyPgM5GrzxltyS
D0iKZGtIxMoxe789EOVmz8bn/G+hoozIzhFSlhUvWc0Ta7tGgeQ38S6EHbgLwIHGnAR97hc0yuEi
axsepIxxbuWtPa6+ijx0NYa88zvlbc2HKdS50qVlj0AWgy1ZnmJ1DsHWfX6iZe8m6vmUzrsnuIfq
3swTCaz9hdnkNC/vrgxij49GMP6USEnnjo7Ltq2BxKbVVghm+Aae4bAkFof3/zDB+flPrukIJr5T
7zFKX3x3KGTCXQwghmlH7XrwGGpQntT9pqtQK5D9W0g99om0DWKyoTZTcv1Y7BUwHmmte2knhOzi
OtIQdK18RBzITLZ5EMFvrPXLHSHkcs+m9jYAQpvg9D5jnjG9Q5ag3NwlV8QaHFMe5uLKMU6E4col
jQESj1HPeTfqdX8R/Y4r9fFGcFqQauGXh/eRTojL/6DnesWxU4TytbowRH0alwBKHF+wsRka7IIG
6l5P7GVfVLXvpvygY2EueWP91yom9jj7X/4onNWdSr+mnXxS0WXNR4giJFvwykTNRwUgNxQsr8FE
KoOaMMEffWV35wfeA5Q20AInyiJFzS1Lkw/k7TubFs2eXmZ+F47a7cuV+yKJBuaEs1f2F75fgTYs
AOALdLWcNhAGVHUUxVB8M3cnaoPvZwfNlyEcSPgA81FqNDEPnJjP+/zsawy35yPAKYqGBcYQ8sWS
CToAcVRP88En0a7fu6a4jnEw7QWl/Cd+YnLf5sDFhVJADrjG067G+6M1jBgiB5QqHY3u9STS1Rb+
TVXle7DA4CpRCg04GgluTJ/8lZmU82JJ4o5afwngrk4LFJRro+ISUCz0YD0d1U9VYEyDOuzCg07J
cUKyP3+DYFmG6GUvPJ0UZTVoFxFZasSsAd1QDK31PgR5136KYzr6g3ByOJXEL7mZatA2tLbRBVkL
OMSWN68/j5eB5CmHhe0sr84bdSnecwP3mYDDVTnOm5OdZIkCr9Fl9Ly9J86Wbl6IV5Wsd3ve+M5B
ccif50+40zpXhLexr9DGxpS7JdV/zLynNBSwPj5FKR/cQTnAnbwbikVnrGYF6J1TwWKX45sMwvt1
dQAAS9v43JFkgGKLJoAgGAS4CZJF6D3R0Doel3Xf9BfPlhci7Di8Xrj+p2a5JgTne2OSsSXvgcU3
62AUkSIbKIv9CDbClbTFo4zfwH0BmHhdgNUkNqapAVQ1Ww6tS28JhpXaw20Q7zZAUpxOKiAn2Bxy
voWLht+yC6BxB4zKWFKzzsI4cBVF2i06qqO06C8CvW6vN1Ma6VFN3V2DmJRlasQ/QHvm+nevJsIW
YS0iHIHMeGZTDXP/wMoIJ+aMR2wdWr5I9zUm/nDP9XHUuVXBnE1EI0lRm1pXkcu25QG6DEEOMVGa
/9j6RZZP8wDM2ErveGtXILHnfXSRWYCN1NaWxKpmUluWXmgxyVQaCNfiK1VePonpWzLJo/bgSNT6
LKpPl7RMYTl7Wg1s5oErMP+xc9LH/qFth9BAzOMgdCsUTbMSpClArqFxe+dUl00qKMkiRNdKaCGB
rkhKje7jgVOhR2/NZ/5+MaX5Ss/qOdJmj6Kw9yxlN/l4QSXvfz9LsizO7OOLDk6rfE7/U9UilqEE
q6mEOLbDgKsoUGg1AnfpR+/A61Y4ZiNTOk3DOF6YabTy2ZH1X9IEXZ+yRuwkrnarGlZcg/9m3Y9R
w8bBgrbVEAKapXyQsnuYUAKvKsD/4nAGLWAneMRa77VS3euEXaSJyHRQee2jMRwtxm/ABxf4paTV
0Qa3W6Vc7H+K5wbZwjYTloPsVzowe5EVDeJ3awR0pAVAM5qK2mZ8MzV0fYMzN0i9XrJ+cXdE/7iv
QoTFK3UHNftFltjzOWbyI69h5S8fO0Nkur7xX6xgjwDNGPUl7ekEsAi2Gil32S38B9VmsNfreRkz
3wx+LgS6Et9yL/HPzbU2moUFbkgGWov+OO7W+t87ybl4Zwg+lh7mgjrMqKqag71EUMGNC0+eH5mA
R51Io5l3lxEnR2vaT+DFaFshtaDFxLxlIdF29HDOap0vX9pdTqusMp249QQCWHoLmJ66z897fTSd
p18wefCwCLLKaUcuVdAhW7kBr0ZyPM1DA/mcYqwV04xe+2v2wInBKGOzzmWCWXfsCdCk41QuRfcw
9Yd1nmU9e+y1/y/AHmn4lFtpC/2+sBQVX6j50nvtMOx7cZkuLmtXOOOZFeBoJC1LUAtHj41wBI1l
KoR0B1Na5uMZgLC56fOgIHMB6OJFnA1yAbyaget6r8o78wPXx4L/LEBGPXzLHdHxRGpF703pxhGK
rw5kVrxdiabAaeuduowllSxr1RWw38BHYfhxVJzdKTwK5jFC0S7+ku1doWh6e3VkRUoeLoIDYKj+
d2FFtXWzTn4cXEPzuH6kAVNJHucy3SUMUZtumWHAxFvRjqLFUHgIEnpcfh+g/mbuNb7UHY1yYXQR
CngUHbNyM4fBkD8bk/EUq/AJv/ar5A7kKJTAkz/jxbygPj0Xv2Cz+JE0oWRISf0b0izMU+pWPnNt
LaCLE+j1GcUpMbrwMp//+601gZAIMDHU/nlsbvRD88OY5zP4su3B9YcXHY2zj7EL/rXBXvopFlxl
87cAkg7veNuvD5EiMdv21h1ROHaN+/Jw+9HVMGEsEcoxykmrJJBWDyumwEU692KDgaC8yq0t75ED
9vkcIrkbYLdt1LiUPk6Eax9i5d495BN52N9WQWNpfLuLnNrRXW5oTIMDTsSZTtj01U62lMu7S4+M
O8Ir9cxJSfZct/Par8+TN0SNG4tRNefqlL/WlV/lUp1EJxYw8Rt4AnsH3Y9EgeuImK+ts98uEbKx
ytLk0rjnyQ2zp93UqFhzIigDpLhT+rghNv8/0yckMAaqxZK93Es3HKkqrmFIO1Q+2/6lS1eAAiwk
Zeu78beHdX/vrRm7FTL/vQOlQfiMTCWCepwft+hYxQr3AW3zN7y4ItYu4OFehYLRnl1Vlqss9jjh
idx+UwHpSLQcIiKcwnbBavO1HHTSJWphQ+/A37fdp++WIyzT5qUKibcCl+zx9c0PnEAIVj2t8Akc
bZTv+vx82zjPFGE2bttymV0h4t4VUaGPuT/cuKdT2Y5WZikhmnaC5OeCHZj8jzb/ZkvhLfOvHtJg
K5ra6VIDEcVi4lUZPuj5vPPW026XaysmWsPqzxFeTXPPwTXB/iLSZc6wuIvj0ZmpKZ+oCbjsTitz
WWNBshxJMOSb5CXG+e0d4YiQqPyHui1gAX0XPOrW5F8YoX434dXHpDlQjSEPr7xB7O4YnkZCzSge
7HjmQbqijuHnRAzfYxZvFjpphof1Q1dbbNb+pUzImhGmUpZs3L6FNERj0k3CpQndUTZD/0pNaQ68
SvxuVlvQ4cyYHQIu5mKtPdgVhtUXBX8aY/cEpqx/j+Wmx1n8cTFMXQqm0ExmS7nJFv1ij7rdOW1g
4zbH4ayqlQ1gMIU5AVAzt0Tt8YENsCutX5XarQtzBuqO46wKheTEyMnwXG8awfYb+NsaGyGyecyv
fLHBkPOHU1+rAUv0/nYZreFrvlpD0ijuqXRbyLd2AyaE4++GUGPfweUxQACZKp2OvAcg4NAEoIdP
emBq6+n92BZwKzcnPByqcvXLKz9nHspy1i2BiR+YsouEL3GtQEKy6x0FF6poP6/mzGgaYtUvv8T3
QOFYGWKfdbLYWcJxBX85jn6dZe4R+W1ATiWc++umeS7QK2EcWS9/8F6szMQ/ym97MaGVMpv/dD4w
RTSTS/LJSQR+uBcLpG+64O0CAHeC6ai3G1c68XNXSCZY2fkGBIc+48BfvlOczOiaiukSz1PAzOfY
f1o42KJ7NP1Ua0/sAIfRLuJSCZ/yA7Z8ZMqueCkM+e55cQ7QzTgm/JUyM8SPNkVU/CGiNJ4Imz7l
UsTi9yuecr9WtRvAIS7M4x2++7L7XUm3waHY1HU1+JES4MsZETWw0ZJx7I6HFAMOmyc9H2pCZs1i
oT5xoVySduTmy+Uk9ka9ozyXRZpdJ63O0ue2BPM1T6L4XSej1ePQTUKJyjRBMF2A/j8RnMVwhIun
SoRZCJNDqcpHDQlgbC2R9athawNHJAZeHaoA4X/XsKRacXiK6oIBma31FrWPnO55RrF+yRfH+9Nz
zb4sHHujVd9GVzOM7NA+dLrVU46xlge+WphIE7yqz5oblEgvQ+PS1YeYHfyN3ETNixTVn7xDIlD1
yQmdjAJpPbBlWxHvNx7E4EYw7rAWa1edkGArnVb7yh6QfJUNLfVerqjLMk8/LtiKC0hxv/gQwuZr
fC+SM/7s2hh2dCqsS7CjLo2v71rfjXxkJPLvFgzc6OL+Jp4+HCWIE6sBnWVy5xM0e3MfjZ0ZhWCr
rnq9Vwzy5G5QZOOzbcJ4AHYrQbZJaHylQ0JpWnw/zic7Txx1TyNIrdt4eu5f5oq6FHHhtrwLl1Rw
EAlpGymUI6GRWWXmw8cs6qnnc7irsxkPP/kS8K3/gfSxUzjn3YXwNRLHeDC4xXOEans6Nhq7ySv0
hoBVukMLezKinPPV0v3rpM+YgOG1hD+9UXsnYahuZuv9SUQW90shwF5Ezdm+1w6m3BmQjKaxWVg9
gYPigI+SuM6nKKO3Z0LwBRaCc3pAV5R2REmwLWYqeFnwW9YMTEKmGbRRfFeUAoH5Jbz2m8vcGZgl
avq4LcyGwO0zKY12sqmo9bs5xkFc4onf+WW4Xp7Mnc66hICavB6YW9o8v8Jeuii4Rt9pCo3bmtHS
X4e/koBEPwJlugRRouMo25yBh5H6HlbaB8K9OQvt8UWna8pu9iBsj32P2TOAIvmc/OCjZfYsJ7oo
xSQlcD/pS5Y9WVVObCw/gGzvo3VimS50FQTzOgDjfdXhBFfgdMCBzMUvqdnGZKis5YULQvNdxkln
qhrqY1ARgKmKhPefPblIU8lYw9bQQQ/23jzt8TRCVEJFv7/0NWFMkOl8+OirjiAItCih65mk2PBH
U0aKeCi7xIOwsfQZoctYfo3h/QiOBOB7RZIeATR7C6LFJvanfU7io+vJyDxmof6wWq862dxM8xo0
fnx1d4Z1mulT3apjHO8x8EiaT25YhZDM7ZhpOIHHn+doB/0C0sbggnPcjhU5soYFoumGY82/nwMP
DxCHBOgDrveXImDDDN3Oe79aW8IUjxUWApblXdlgmTispJ5wWw/FqXBdTv65fYXPnCo7jjI0sncn
93UZOtRfUQQohMffT1A5/tafrxex0N7FMEaxEV1qZYMe7EPW1T/d6sFmkixU2CgoFZzk5joWOWjk
d9jnzqWRRMAUxnykc0Qf5OH6lvjdUAc0AulCxZGTghjl038oGNA3WHk18WTfGUyZqazmpof8i8zU
b15DeNaq7FDumiMPsYjtHwk/6+OfJ9UmYCNkA+wEjJtFGk/yKELwMkesnWyJYSo/ylAKDkxVyLa9
VTtDzLFpVWSio3yQbjZobK6yA4iVdJEdBZMWmtQ9FyIXRR7A5L92G1V92zvb377bErx14AYjm/Ob
/fmoFHTMsk+KeKwJZN7lavKYbZQbfvuF65DPwBC7Sok8nLyXehKZBZpWes+TbPyXq4oG/sUPcLu+
3hFs+VeRF8YYOolIi6EP4jRCsXac35Nq4OW+Kk+K8s1qQRgVbfMUK9FlqUCNmttHQE+22QSSmDoJ
Sh/wjmG77UxYsCIebnZu5OK3wIJpPpbvPDZV9cRY8wDgf9gUUPJkzz1qZlvWbPN8gpU9wdatO4Vm
B2KVsCqlnldp3fmBzgt1rmwPsm3xMRCdwhOOt2YuzWMbWR8FF6Hqe9Y7Y0ZnpF+x6oWzFdl7ZpCo
NBxFANu0KKzszQdyxfJk0bN87y1X5/FWA+DjUQitcGrVA27u0pAyxbx5pesUSO8nSPk6PTAbRsXD
lUupuzQ9vPCBtc1ELHfncUiL+BcutLErIJwo51D6UXfV/k2BdCIQNYlxyq5EdPn/5cSobWISvOpT
QyuzdM5w1nNli2UC6Hh38Xzp2T9Np6kHI3LXckSuMaFeu0PZxkxfWGlQOyGQ3DM+54ob92K7QLeo
9oMELPMfv9JvT7NX/NJrYY/Ck/KcxTRuzQvbRNz0910YmE0d++CWHJOk/l0UQYyonFnDrUE9Ij3f
ANx1OnHMlUl7BKJGRcA0Z7uExnwawudYwjG86Zm3LwDpHl1zo40SguqcmGmdEtDQiHUQ60pO6jOz
O+gXrxUz0ny5pt2DvFxahn4RjFVzp3rYUxaqCJQCBHrbZ8qSiByCWAZyefrz6cVAq8rITmPHYLek
yszZdXwxJHo8EjztXIJur/CAYMbnXiscGKjuVkGkTKMBriOQ7zyIHA1YFWx85wghaV7HS8OBsURH
mK5UI0hk9ECMEomPnv9bdX1TfFl3h/Qp4pn3l+jq+sEmeufX20m7i/FIyzKSemjBzeUtMWgOgR+3
Yb/X17woy2ZckcqAAULNGomdc//9afzOvj7hnrjMt6D1R36wDVHgSVflM+PDvmWEbytpxLEJxDTA
mAhPkblOTZdjcWkj5WVU0IMMWe3I1ItczEzp59dw6OLrMSvqTfX2OECO/mO1lmDvQjrJaLbsHllo
LNGzVTp6qaU9UOJm6VsbtRHXWXQHWHBmr2qg9i6bhdCMuQ+8ZOsjFDCw+CEepgnVefyMQhlq7aOW
aO7sqVF0hHiI04dWb9HTbGAa/ujTkCUldowruWVJ07D50RwrRv4ALS89SQE1+/Qo5JKlRAC895Pd
I/bZdXQ/UsMNSMBmr2ge9LdP3/+oj+MtP90BAXDIEKOrb+eBZ7LEbnjowM3Jvp3BFQam0lNE+pPe
s9FIcIYJ56JSxyMBy/5CoKCEwR1BISe/w8c9PlnwE43QgAkErXUeFyozsIbm39djAqGXvdFaMs15
6YfaIxaVYYmoCrdoDSEhYHGFGgwcd8T7Yeq+onsEQ+BtHnHRNuv0XoZwhnHXCCTH9f6j2kW1wS0F
1lBdSTQoJQQgh+UhNZ1NQkmebnbBqJZiq+5CWMQTF7hHqxOPBSm5dno6KhTUTUQwdFZnN7ZF2I4K
VWG+R7VjV9rT+LxfP1fQCl+tnM9eqlgnd/R7S/kDd6PjJn2c9xH+cGvb4A3euUjiyJK5EBdnawDZ
T/bXNpWsrA4MH5l50drjnW6s6JuUOXJHiYJdVtUmudp+//6UaouT8tEBOeIkUK2wJypk1NpUu53A
a3GnP/oL+UwnP4BHukTh93csfCHlnSLkkU/iAXZYBXdVBCrZwto36F3LXgAe0+i1UzEP5WlL5EGj
1Nffmde7H5pYpo8R1dD1v7ZtZONJvoWomDMwduZdDnm0mujx4LgjFfWi1yUbZdNQASAOtSabMVWG
eOyy2xzPjJAvYazoKbMs09NsXN2RDIoF7ej/LLjY2Bf07jCm4LWfRRqgds6C3dB0uZtj++hGJ5y1
2fYoGZ4jEGUGdPRQ3QoYKeI16931ONQ4j8pPFU+/sbA2SxrGjFgNXw+nJ8Wl6pK6RiZG0BcsYpmH
ZMfWsYOft+wKdYUMt2tGNr8TpuxEP/5HXWA1X/ig2BGwb5q1MjF8HMN14rv2noVp9FlNJc+5nCE0
Tl3wp8Wv5nAzyUG9cbOSEWellVAVYqoE2cmyNkdpAEVaZxN432nyhMQpR/Tn9/5NhFad6xr38a9g
JGZbcCesEq6fD72tKzXaukPjG91ukF4ORHHdHqxz8zx0iiOX65kK+Es+DLfhX0G13NpQJpDAfB4z
8uisjYWL+Gm297aTuCmarBtk8e3XAA4ErfUMWM8pAH1XCH9pn08YHS9dhQtPNy75tJjCRj05/WKC
b27KizWSS7H86sm68jM8yNQZHEi03aPGtko6qvELjvNIxMrgGlNGiwNA3rS4j5YaHkLHKrs9cnLZ
ZtHZ2cIm8uJgEaQ580HMD7jjD5Cg3WaNV8bq7/+Zay2m4FtSH57dfSvv7twC7ivFH+Qlf8QiSK/4
5xhBbEfjp+VGWA6QuHfSnO1Zr+g4jUyxhVyOENrrpR4zzD7q4+xtuTIQWa/oYKQ/lWF46aq6+TSb
FONve2g3P/umH3rZ6IzTpUXtXw7DMHX1AV+A7xS8brquPYt2IK0UpdYCU1uZuzbNmN/iGXZUleX+
/YurrOHgFMJ2k2HxSNsSiMyFophV90XHptiP0qBromCUkXpqU/NrpuwCLW2TfPAjF0O3m6UFwndl
ywbn/KQuF5ZtrVJZBG6JCyXS34Z1T+lHyoU6z3JwrE9e4iw+tbv76R/FRD0h9nccoInp9D5Ga4tn
+q3SQt5SXC+poOIrvCemhoMaJj6Up9pwtP2mJLsMYTykG5vT8RA8DlNbJmcUJty/IRTkk4TEiVDD
ibKQhbY2AhEk4/mRMrmNXuwXtedkdyQ4zsrXTEWInhAhcw1qM4DR5ka3xKvUuXaqTIAgxG3QabA3
E/5InAGjSYo6QMv416MD5q0Yp39nLEmu74dPqHWSd63awAex45ZPEeVagkfYly2Bj3AGZNzKF+BS
OPjY19YoQ042hz//7/Hi/kzRDo8VnSM1HSmsc8u75UEsZ9tnCIYqs81y50S1cq9O2ZE8sKVEoqiW
DuT2tLJ9jU0qdObAcUHIwdqeLxwjk6w0v97B6sTtu3jDhs/MRz72FcLxNebR3exra33fjOo6o0WA
MNlVwxG2+v8XvV04lDv7dzOAWAticKF1C1KEeu2KufkKNZJmRCa9HHvLPO0LMHMF6sDoiYuTyLOT
pxfEP6xMdKGNn8uBEQ6tg3DXpqKEm0RUtxqeOnLEvMA1NeWdG0z/W8m3/WE2/vFvGm3T9xgBg/FP
zk9hxCPemqslEaHQXdmT22unr75axr9NuJyJNzyFndVitIVBasZQE47j+7EfctHf7Fh8/NLkDz7q
FdDravfAmmC3JAhyWOS7/xXPGwRkwN0D5h1ErqFqB188qWrocAW8wEWSH/fyOnAcQQ4bU5MttjLv
bMMiGJrv9UTWnzoXgbyanY5Op99v/SWDYUdwq/CNHfNp3AFUt5mka/7d4lBYOrOiFy9y+7YM/lrJ
Ve8CTRVtipV4ewxxqjoKLfY+5ef6/xvoJNURukDPW4gXLJrnQYj0vWDHhb+7Txd6EVH7Aa7ct8eQ
3aLpME9IGVaIDWuzL4h9YwRLCX/TDZY7m5Rkjbs076uUx9UXrifG2BIbAgozKXuIhvtiqzTDHwce
jEAfVfRCah7TIPOJcHinzNIUEV5fzEvQzbhMN1nDvp1C2vblAzISAm2bq/1q1r+3tDsMzOYBUgZ5
6j3yPzdelGELZBLp/pSs1MkX4im5uKG+SwtEL6yqIeF0adtCivAXOzhWgSX87W4DgajPBT6fJhNL
h+Gd0dsFkPly99UAcLQHFPpzG2l5zRnKzN+Z8aX715Hfz+mxCF0XIKT0l+Raku/1YpgZEuGRkHN8
atwUJBnRYenCfKjK8iPfDyiufGnOmQtxwa0Ve+X1TBgJ+DxfmqkJ1k4H8SKyb1Ndi/LpPOvhoo1d
a5BZJ2iAVvBbxKCzPQzY0cJAVT0Dnty/F+kxUwPSMI7DCc7+YcBURXszxUL2H/3G43vXoQHSjnfP
5wqdUI2eyWgoJPSBX73gqUnpGp/l/SmmQhAfW9C9aze9lzVopEGn5+HJaqBhOkuSHeqNxOeziuRI
IzpERCpwdGDh0UBAghuqWfkV5DJhiPO7y9DbYMv9dcKs/6o1lcEwZaAw0Ark7UQss9hz00+3CAWr
3Nr6nf0gQkr6lIKUJ/Dr7S/ON1ytZxNKWBFSBJ0ci4t1Ag+u3cyquVJ/3YbG4XYuAfdCtsPpvBK/
vZ0aEce+V11EaOFbX3bMbyF4jMSZQyPPaHcjTDRdK6/kvXqXqn/Hi28CpqpLO8Zr2Sxna5v55MWo
8Y6HWR3qk8qoLvWjGC3p2vzN4v90DpjScbCkx5LYgZveZSAkfprTXoU3ZubQp0cv8gZsBxoR0kVV
HAIQBJB355FNzLvKyOknqWFv1T9qHp7tvxR9f2tJWGy/D3RcEoXOpIy61IjeMaklQtPT7JEE16K5
+/Ng2pZpxk2scZzv2SilWZsUYWp1SeFtGZcEsSQpIwPLHGn1flFW2bZqZX0YOeSI4sC5z0fqjmQQ
kLO7rVysV5/mif4dbzHRv7yHwddUk4DGYSKZzOjFP4P/eF3lRJ+nbNjdVLGxLceTWzKXUxCWigfm
9mItHAoEVmHQpp7UO5r4VvnrNrB9uodf3oGRjsgC5Q7t3RnIToqWfM2ISmvdF1tMHhF5jkn0YmRS
4UtA0eAQ0X+3yEF3ZSLN9L2R9dA8ARD0uye+Nq27+LA8HWx8RoiuI96zi7IHHm62RxeyADdYmGxv
zQmW4xyz1MM4gY74Z5/p9RZhMVUAHL6WA1LqsfvVKZtdbKBTJAHrWbvfvnXxSvzfvwrFBUW2TLiq
a52sILSe7AlFv3BZlXxw2cIYHT76dZsC1jh840n7mBSjiQ2c0PV+0xNcMMt2YPRi2e2zd26ng/j4
chVOW1E6ZZxY7KHf1u1j4JhdWFAVzR28g2GKs6RMCSVkMyKLIDb//kqsFkjdUR7ArOB59jQTZtqP
RCG/jr+yxIJDw3DWDIlDP4zR6LBajlBJZpU4oZ1Rgtbi24/IzCNa8DA5wyQCIHEGPtntal3dkLNs
nSSb4d84h1n6Oba/8YDhQnzG2BRRaFmK1Wpa0O276A5ZHe1QJydEv4vglzbudjWJx1pm53K1siM1
yzAzhvy5Z+kIjwliEW9iDptPbpHjhWBPqRoddPpbpqpOJ5EeTelETUuMkD4rHMiRDjmIPZ57Jx4y
5L8qGrLDwGLkHqpnPALSPoueaZ4wf626Nli34M66xn6eh88ThOD/cmjzo5cJ1aR4AWncelbFl1mM
i1/U6Rg5aHtSIJ4lv1GVzJTVKNt6EDvh/WBSFNptIUUNOG2La/sKWBxfVl77pu8p/+++b2sYfsHv
2nA/FyqmRJf+1dUWc1L0c8DSwchYQgk1hMWGWooeAYK/Ws2JYuhuYXjr+oXFfIYQollnlsHka0Bj
5K7+0WALjQKkjSWmKOCjfZm2VTB1TdwjnuRKkpohxykUn8behRFCTkyf3jvXIONNee+uiRahBVyy
DMR/xsc8sVKveax7xEI0B25N1efzyq7TkAnSawThMrd/6ZW6MnvyeY+NiiUbvMQfpTIbMjI4t4z8
So5CJUuxoqiOTpymXb0sj4nds/JIUypDUiPeHeSzhrUlHnCeYzI++Xam/GNdJ/NiZhTWhBiod9+f
Xro34qvRqCvT3qP/26wZqTCE/ey8wHXzU67TM4YZpTYMl9Gmq4IsN9I62OHaB2Yk/2bpCzKevZQL
UBKrQIR8am4xIr8vWf4JnDdjCUGzaqAMPqfQbGyKO5zq7FhUgYWTBOKIjUAFohi8wX/n4OIapoBV
NF5PtapFYjhIgpZn09ibG38RdujpcxwV1N4aF1WvLCIwGejTik7k3VM0EVSENEm8ob/x7lf281W2
9vaNC+zKkaWyf+mIX7gX1wmS3sTu2vkjf0RjM8L+41pA+PrTWcDQ1NSIbsB5tdNn5mEZwNZncDyg
yMdPvbYWlPClLdgjReA+eCnXoZuo2KE9xBso+FQ5aSeTnTBiqPl42kBKIQ3SUZh74EPTy+eq8zKw
JonGxRNt6UFrsKMbERcq6O3aG03KrTPKPl9vhYcaPOxiiQov7JAmINHg7EkaXthpF1IOeVF8stkI
6Qllg1oopISTRGZDb90Vx6IFedQf6KD+RAJ3SY54nSF1IHXfnp7760OXsHCX0+eFDzqpXXlD4c65
h9rVUdISQPD/fwVqexkNjAUSTHZO+I4LP72xvMkObwgdVSJObYvfOFNy/5uJF3v9LTYNHRD8QcAo
x4sSWhEmn8kpA+Q5MrIE4sfAnONEz+6e4wafjBj4/3DZbWtEwECY68K6gekePtHc3dlbfDfAfjOo
V8TyrTDHP9Dn80Y9VGwnz5Sjfk4F7DlEFtZp2o4glFY4rdYdYj6ysCKMnL4EJ2mTRG8ekcmrNZLd
rxD4pEHJP7IBDyL9HA0b7C4uOFKqAje8nmg5wDYnhzz/p+FfOvPg9yJKqaJ+xKUiF4r6VFA/p09L
qw20WgjYoWw8JoEknNFRLVfR/S0s9L1/lo63+pd2s1C7CtbR97qFsqy1ivOQep9yfGjh/flK+IZF
cANwpb+yQ2Qw21Xv9yZOsgj3QGbcU1HgcozFoAG77Cahu5OzZ93h/OinUFRW/1agjOFZPCtU0iD5
JjBmW/FpMYKSpfUa6eKDZyU3/6zyfD3BYeQsDY/3Fyz7ewreXkvEQosweEBk2PR0ZMtZ7+QCYXCC
HGovnMbJSun2+fMIYqIp6VCJ34+MHeoblv1GbyzRyNolkGWmQ+3IDzdpm2eKc5NOrNMLOHzAJeL7
C3kpM8lNF3fLznq28XcS0cNkY9w6YiptoBNOIJNx6nWHoVrRO+hnZnSuZjMeZa/Li/fejzTf6HEK
gw1/TYP3JxJedNQk4ztiO0sYh90MDmjKmQc8g355YBON996UfCzVczjJ8iU3QonmInhfjnC1avC5
Prwe7Yu0wuFi128SBj0YGCv6LvJPi0tz+tqLfT21algGyNBpTPa3g7k0DdyWNtiAClfGeoW33kYo
uzyLOS3M2HbJdaUL3vHKZ9Eu8zhFHCJDgwvkItXOx/dX+M7OljCqYcO08j67FRhv6rijrQZpeQwO
7RhofbtPETNA2tAcEuMUXEXf9e/kksmYEvETRMHpLjfidZXNNgaJDbVV5mREldOc1+ylEgivxipU
TsrVmtOwxfAego5JueYT0yOjMrbrOKPPUgaq1RIg8ERFJXmnj4n4xC+tNmtbQJ3Cky24rVHG6PSy
LMmpwwt5XwouaBkIMpoqeHC+y8ycvrIuYhYxi0fCj1vgCAjy7SyMbLGRgiWTFOoV+Fb6CtuDJlnE
JTUqPUvzWY7WuveJwUFdo8IU/V8NP71UCE3/9zNYGIfGQdorIVagHZPMwqHvTaF2AYn32x7mZhKt
SMb8TtiYQNSpLkmtzJWZcHfkDAn3q3R0biQixzlly1tQG+fhJO1GTN8vpcyCMGrDODDPMouTHOMG
nFyLYerW9ylq5f//2fMOEmSGB/xrqxI95krBJOwHCC4SIQfu/6VIJM5TzBIEOMFXSzJSdDUzgcdM
pmZc1dK/GVXcMYKO2m+8ToiVXz0rm+hwMCJee7ZnM8ZjmFriKqTMDOkxy/CfbPJXPQCQf3toUXZF
jU9hvzN5zeioqTGjQeEqqcDzyl3W/gQOk6gaJ+e6QvVIegM3d+2xm4D50wD5xoayGzrZ8Gp5Emj4
86QoioWx+F8Uq//Zy/W16JvBFcCsFCglEXhrt/Fy4hOJ1F4OC3/pH5fqWzhWk+slB8gQwyucjFlu
IOEtS5yW5TopvYaMgu3s5o1fw9Ocj5H087C3UI1rVHHRzGQka8oUq3iG6D1O/UjswYB2YD/spY5/
+P+a1bzsKlyL2zRBXvNS5Z0k3wR5f3z5wv4WsvIfYUjDAIVJanuayoBu/lHytIYXNww9iTdghPH8
7J7QllsulvmYi0IPVNKSRJUjjaqSuT3uqu8GSrM8xmTXJmJR3FIwgoS2z4wQqzPfenIqIEhuF0Z8
ZRkBzGFL3L8W3XmovqawQhtdloOXfJF0ASOYApBHlg98Z+Xpw/YWQDewJwcAx7ZErKtKByPnVi3t
8SxPEsc9ymAbbrz6ELvmy0s+K7MmcC5ssREvGfk1KfMe1DI7FD8It1JScSKkHZ+JL5e9e6A1Nyt0
eq9zyCIZGAQR+bu2aBSxJ7caLrrC4Hs2tQkukSrPLlichEYD7+WFBGPWnta8AqJkr42TNwqSsJWO
iDdWhST2o3IHKWiW2l8pVV/x1BrGNVLRdQMBFt66MRECpLhXEb5b8MDBuhV8pIdpqObm0eIY/fik
CUef14RsZkxSMtRtzRoavpfDe/mJND+gj58VyPjKakbcJeMcOD2ig5r+xEh/91zbjBVLIOnTG2hM
CQlyNW2gqS1MfFBxro/hWexZWUar5FhstsRFKWcgY32YwCcQrAq+hRoLWZXmpF9dpNSZdU90quQ8
faFAtQORY1MGVyTWOpVkulxqMXMvnXlYqKxhI5DwXHaGB22o8LtAb4O+mrhZOltZelJZ79laYrg8
i46R+56tMm7lygBrH453ajjA6tNDzYOC99AAhNm0sGROpGo7lsZX8W/32ywY1uzcm7n7tUZTEq+O
+KOkEVaR//rRc6DIwWS8vBW+GmDmXzoxmix9Avz33TWPxKIBd56HusOVmCgcarLzQpHs4Mui25IY
MvAgdABNiP0VZNDg4j6RQRkh0Q7JEkTQyjSg4xHT5Ne8W2p2G3e36XTFwJSTurcV0yPsL0npuSmq
ZXJU9J3/btWM+MqvvGoH+tXX2LgKOTExpcHzMUUznnOijNKoKSCSlQ0aosEAfk3Z3Lo5Alrn6Vvs
T0DHr4g+P7GDTO6xcjvx/+083i0yJSKDm13EcZ3c2dyl76/uZUtt47cPhqwJ0FmtkdfJSVzX1L5Z
UQdga8qOszkfCUmvzvko/1i9lqHtmSzkZCbJ4bNMQRRsvBHo03k5tX39v3wV1RuFabOkDHB7eUWl
JrGAqaTwVFJE3PWDVee5SMW8hP0vKco+gE5MW9rtAytQGx3du0f4Qt2scJnuXTaw1/pq8Gu3qb5Y
SyTFFvKWf0GxiZMQbvDeSnKUussQeCKPkuKjuBnMHTS6wXSbHdwGiBJ+A2eLp74ifyZC58G9UTqm
+/lfeUZjvi4g/C232mMzydMqArU0ek3ep0TiLiFjHpjesRhEaAx2BsGHIgb62hV3Nk00IdfqZzXF
gqDlLFYAbpRSxPUnoHHOSAYw2HSMhhdYgoIqjE3iZes/c8O8DCIWVngnjw0018Y82iFvO1B7EIz2
9WzHayXv2Pj/wbmpptkLkL/zaLkQmhhibYTkvVmz9bhJq6hGlkem8/x9j3V6pd2WuJj5lUyv9i9o
zDxj0LGDb69tC32v8e6BfQU3GlV9erC4uaWGjGHWkCYYD1/XCkRkUrtfbYfoB9BGXRYfE7pTYnXO
xQpwiGtlBSYz3Z7JAsAAnY87RWJ9NFz8NCqt1WV/3DvPcmD6/Pe71K6xCDuzuOVBAg/EtxO7kkoA
mjclWBQ93V9uPoH+IAQaT7S97NPIHojG+gcGQti+mSAlLYCNJEFVHZs/IRUHEuFgM+P03KS8s939
4CljUVozdX4V/G8bHx4LeG/XZXW4rEvzcKOb5kShxMvHw6291m6UN8K3onTeRxHPoS6X5GEm9yal
dkRaIiFqQNEevmmW3fApKj+2iSvx6uPxeUZpRlbmJ5LS/6dueMD3HS9NQh29Sdr1cnj2ZxJzaJZF
7nacfiBW45/3ap+8TChydM2+UbMfUWSPPwls5avatTyE3nt6jkQCAmJc2sXhW/o90VHJ4BFmE+/a
gQ/zbHlPzlOY9IdRapyHvqMSTVwUhaj4h7Bk/HesG6gb8gAEjtkolPxtTedQUSmyfctuPPIS4UGL
LwDwNN+RYWIV6T7LM7WSJk5D3fDV8bVhrFaVM2rKD7+yNfbUacm04j54vdSOQJntdkPaWA4eGlUF
iyhrdvw9u+gjolHemFrhtK85cMTxgyb2DC8PyOMxwnjEJms/xytGVgmikcD7RVw32oiOEsAJMeou
ZZmJ/ULMNKhF+gipS8jatBr5leb//tx38udlzN+CAVd9YkBWPYbtIE9hkSEhcMQZE8uUCvFH4mfM
sAmog48kkpFpJPO0V8UipDy0nYkaNFAIRlycp/A6ADLQ5y+Nq7/TaewlBbyoyrMzEwiS8QNrQZvv
tGaNmIVkBuIYwczoXZXAwZSkXquJUTAtf3Z+rBTrwF8gfFaoCXyAYUm47RNPUGS60qn7Zy7gdr3N
7guXDKYBFO86mbeY/as7UiUr+lfDQ3wJRnlBCsUytTrQvTOqknHCkaO7G3qlmBuZZp0fLjd4lACG
5WtvCqWaG4EAz+hJi8BONJD+Ie4IgsTox4sgaldKUyaqlLgErQWv6b5vWZqsnLOip7Cr6Av95Xar
J4iusQUM764lWr7+L0NZSf7lJBPxZoH/IPBfLXh/zezRL1FxU9r36R3FSj2NvEVGBejFjwiGjsKi
WMmCClplMMaXlWoP3CfzEPgreAWU03b1b0JvzrEii3EoHzC6kws5PP6yaEIyHAbm5TZZtL7ue4Mz
8sn0f3ZGU7hWWuDkoxpLNDgxNFPEq5uECUE6BBiTNr6ZqxB2HAZ5u4F2EczFa3f8RoA6iNLHP1IE
arbJr3GVJGNEyX7NFCkUYCOTX+rhQPVk7j9Yo1ZA9BEeGU2Jklq0MKzVq3oBSraUjXkLIb9sy7zS
W+CPTUchoWWvd+5KsB+DJ1VcT5gxgyG9uQBSidqMQzIY/cNHUsQe0fQ67ELZ8GB/X/Socb+yeTYT
GvHWRfH4+o1WeQgp5RAFbYl5nIUpiGB46gNHVkuhxe/BBlkEOemT0yHoyt1hSs8lrq7yFwfw4JIW
9U4vI+iRO3hdwlD4aer/TzsjIGomVJLTfw/bYCl4tfmTCUSf0TsSusbkiihoKFyKfCdi/+6u+jk9
38BeI8yZE7of3RF4nceWeoIIYA95mpL/yM7RhP1kMvDOAVXCwdea5QPh4q3AkkR86Zx5cUhFjJf/
WWFaAVLYr9NVUHL6m054SXp2uW8sAWB4JypNsRBWn1SqGs8b04QO7/kae3fSdRDeF7pbAf+rojVm
6RsO8J2yMaHtGLuxM/UdHfVng3ahxiF/wl1Hg2GTUoAbnwSwPSwlIGx402hY+UrTJbDY4LVSVNcd
nfeenKTOu5kNrXdrwj0/w5iC1irucKQP87CqRBGmqvreknnM+CsA58bMhyEXugHg/jvdF48YPpwZ
QmUonnr7ry55wIB3UQea/wBXSc4L5ZSHTOLo6SANhnTmgKapW0v+zfg8UI409FBrltL6zD8jvGaQ
ph1GayjmFNBIKpmKs4ZJxnffxe7J486Zb5Jh4XAC5i4LDVmnlAIYODfw9vm4VaCnhEFDi0ps02+f
6YiRis6y7RDMVeIHj6dpQmD5eyTqTuNj+6Qy0lzaSBHc/5mPCZ52vJq/t11Jpwfc7Iv2IzvFnccL
bkgyWCYnN/JpH9PvAPFbUwoQfizBzREV25BPAW1c0zleWzkZJTHuQtpWgt8L2jeSATw9VFgo6ndz
G7UjBink8RBCTBzwLQzysrlfK9bvi0vhSF+AMebTv5N3OWys0r0yJu8wJn37//InvI/RDYOyk2U0
rzcjLCFw/YOJZJZssRIJWPY6Sn7gGmorAdEGO+sXipq3PdvYXn5yuikVBviKxfZwTxpdfxywN+2N
hztxSyEHuX5V6Jl5OSkbMMdUUjy49o6b4Ff6b23VXlPU1/3PNy+9SCEiSxSkCvg3nX2IVtIt+zjY
hKDIPk0gZY1h/JEWCEAEeGOK6XoAOPy/8m9t/lGvCrhWt7mNXtQbcKZ+XGQpHasY0UmMcCVjzTXx
ezzt7zLyoUEizOBxNh9l1DKjA7HlG5zRraylthj9pejOSNON68fxIeCPbJ//FyM8hHHKz10p56Wj
S4pAgK765RMYtJK0IPaTs6q+gJ6o9ySYPE5P4KInYpTwpcetcwJf0S/hQdx2mTjtVU5Qs45s+x5L
evDmVgjejMRJ//JRJtlEfXJWdJcxmURyFKSl737JFTGCQ3JhFdclj9g6CGl5eaSXyuNMttUuy+s0
6yqfbxv4390/rAtSDjavzlLqmNCDxuEjb1tLxt9vEeQY7iPYcAfuIUYVmNez8yyJYtbXjPrU18hB
8hPJ+sqNK99JSuDBTMGhit/A1O2R0FjPEp3Hl+QrAqAdgz0htnxlLEPqfgEyEsynRA1xoX1bv2P8
22AFXBUtILOsZVaC6rGs/5AWrtfPGXH8THi5qsskCZyXYDIiXvjur+mDFCZHr+hnYyVMxVryBRBa
jsj0rOuXuqyTJoALO/Z5BqrP9giomvuVBfbdksv6iJwEaITkuj2aJ7Cg0UvrCB90aQClmpJZMfXV
ybDq8Any85bRmi9t1Si0XXiaWTlTcEytVUYxu77ndbaZNiBudM9FQRmv4JbcunBYbzMa+vb55dXe
vVA5mv4FWzgSEVNZqokww38L4ccWms9n9HPsZ9Lqr+aIPurmfh4g5aZbS8s8nnyaAb62gEX963Tu
HmmPCCiETFH0z2CogZf3NhsTBNxTlXIhe+Fi+IgH1EmWH4T8iqGSFU60hXnuVj34OTN8tM21zosp
rHDxl9tw2W7rdcK6sCg9abTTj/ww1hR//RyUShaahrCSdFbCIaa2mYXY0FnauapCJH0tSpAK6j3X
tb4bf32srjFIQJ3qd900nNLxCcGRB4ZkGGJc6uk5Uo1M2j0ZQpT2ixFYBcNnRs4KUbmRNR0i9uZC
MuBo4HgXIgT2EF2cUYlmm1DY47logsLBnXJPLE9GB6BOMmHE1lHpdO/aYLKJHjpRxHqza28x8HDS
EHNPpGxUXF5byN78ZAIYKOCs/394G0uPyXU0QE+z6UBKdKDNfCWbTm+bx9AWR7G3pUNvUVOI+wCU
vwJJNoPeDmqeKA6a0zCDlWSPLVwoDKs6ReN59RqTE38iztnbEVnm9ywOXRP1TaHcWWn4Tnrn1BJL
v1MR4iF+rrpgrN1xzWlAN3jEksS08BQhJlgrXIrRZZF4JwtQkcK7ZKd5pETLcyfYVkfVAowmQS5c
tTTh/jwNhW53UIj5hf6MVEboXB/CkdLpg9ep7vocmIkxqwsB5OHn2mULQlG/cLmTnGRrg8YdNxHI
6LeyZd8tAVBfSRSw3S1DXLTpkUERSmXvQNp0u9Cl1dIzlxDXATIckmCKBsW0mzIkRNRa3S+EsCcS
uzZ7DLa1XRoY+UzqXVZuizRiqJTBd1OmfCD6QDIhQN3XYhxGdHYzn62ppIPsrsqDNizKWFIAk6eP
hOGvUkwKKXLqec/yOmii1Qui3kJsYNhZdCbQzZ6oJZ6585TDoK2nXbpsW4v+7Mr3zu1oRU+5UckQ
ZW2kzI/x8pxKkVdCZYXNL+DG8wrpDkhu2Cj2NWKxJ6/RngHwjslMROX4O1K46wrioUWVgEBRyhs0
l+QlQB547e/VXxRgKD5/O7xe/LnMVMGomYq/13GOHIcqppMfMl24WGgO3z6vIwfhI7R8EmF8vdzd
kvULOCoCw+ykekZD6jKdfBf0qWV4HvU7rthWEwKCd/WBLRro3gBHqhaNZCMQlJ/rApZKGEAfel6q
g9rNwZhPFNcx4GsxCmwZ/0o+kRrp366/kcrV3RX2X2vdTB0+o7MGC4JLXFYKJ1g3wm2Q00JNPo5R
iZsVNG6/SbChcwQ5jsJdTfhTpHBInqWN6G9ZSZqd2Evy4BCdNOLi4XiQ3e9FF0QDV4hiti5mPTum
+vXEkKWc/9hc75mpZezcECei7iE4WzmPavF39KPQtYIrhz2TwPYKr6ukw+xSl4Q0oLB4l37gvIFt
hrSy2k39At3IiCDQKH+/88CIyjoSbjRvqUT6PheWuzlLGZhB6O6wue+JvoPOkTmQTBSXAeNa+DnP
MJMdpra65UEbH5970QiwwjIDjoA4B4zqJHPQHdvAqMDVejljffY2fYA7nZV+xKGeR+WmS7rBA7rM
yGaAlBCYIFRVo3AoZIX/+eCZH5TuiJ/+2WkEwRAQPj6YTL5jXYwbP0E/R9W/9aIFcKiaKNhMeNTM
hZaCgbjtxu7rkGFpEixtd7qpTaYe6Kk77NzIA18rzhYFlYPk2u5GjSwMYJfm1Jby1K0436855Nnj
iTP25GzIKb89ql1Au1INsdPeAtRNRsSYhjaLcpZaxHWcjO9Tvye4dUIr86C3rimLIMWECpB79WSv
4OSsLXACB1yxl/uWZAbse1bcrRwVqQtlH+dB1M/2ujQCuhzksHZe5tPXCXbVA5mkzoN8oIfwMuoG
YAKydOPtI0nUN7l5m3Wn5L4+/2BJMUfU6xvEI7pqzdp7hBwY2+2bku8WQq3fppUUZLgJ1Mdyr7MS
Yrf3W2l1JW4jwY4t00PtF48r9cfMNi2dhwyyL+0lLaZPRQomd7L/vaLPE14FcLIZrhAiWDETbKsf
TyrjrERHTpmcRpUNp3JSY7EOAl4uA3nXx8HskgAbnjSaPndEKYCOpb9uPQLQTnOZsfXOMTIaDVLu
htyeyACA47vp2AGRu2t4fK+voAlidVI4bj/XnX5kW0P04hRxx3oJiXy7rRwa+QThXyyY6/aU9nzp
LF3DcMbSuK1s5+MEHjAM60clVKrJ5EQDoBnRaARfkqbHgUCXOe4Ep5GRqn0Ptr2xPv7EvMkvn/uo
pkqrIcDSW8K7YpEcjNgEeLPPI5vo3Bg9IBSHYi0EstrVU/3aJd6t2alsSihAKlAA6WrW8Y3hX6Uu
W+4MBCk+3uJAIlZ13eswK5UCSDe/jV0/ZRzpMzXvEPq/VIKZJ745oBooUernDp8YPIjM2K1LmdQi
Jbc2lqR/cj/9yvzB3OBDNoFvCqvXwFZ+uWJenaYaaKviUZ2TxpAk+fLhWp2SKppxhlgtlhErsoCf
rl9fEGEJKW0EOqQL8LliYivYBoCDgLuXVo9KXtxaThrBH539IaN280ewQrlWs0tE1qnwQIrNRxXW
8ixuqzq1L+yiSKfo7eFRL7GnoS8fLjVG6LbL1XWR1MygT5GL9oNDYDqgTckMitZdBMoqOwiZPVhV
UyDLIE8BTKUjD4QSdW2ftpLyJu8b68EwVVGuD5o1+u/kViOw2DKeUomK/p9SjRRkw/kaSEFKLrYJ
GyFseHBqZvr1yzxmQF1kGltVdfJSzyI9E74DLO4tlRY9Ym98KbDVJTTzDP2kmGLe0YDryaGm0iQ3
F7okixoxEHHiE7umYTdQB2dYvcxGoX1RfECBsC9i9oauUIjYC2bh+HRaX/V6V/U5yPOwCDpzI2XB
K4mFkM7bsWZbvznDwnIAf/Vnd4KMsLa2sn/x6DfryYNQTpVHH1N5QAyE5D06DYI1Rz7WSAu+zXXi
wdy7hsPh//WiX3jMVgWgVqbPZdxkAELSuiFoE9ZtwOqytR9zFpB73ckJfCXbPXZPg0ocghjg1Vey
4hUVgLe6p6ym3NcP3REqDD/6E4+iuyQojut+WB6pY4v22uZiBNOSGlrf44fOhvl+/Q6unN9JsTa+
44xL67ENS71M4FduUCHBfNU14Bx8GNhN7ShfRazqkH9cyuwyCBVolDETBBX5LgnYdX7GvrihBVEw
pURbPAZ58WkWw+SuTXgtnPB8txGZOzMT7xZgyPF7uZ25SVS6CB4SKl6nZeXRprna3r8zFRkMIIRv
3fE1esA4TDvLDgb3uue8SPkmrbih7ifChHlpiMxFLr0sKmxm/vjLA41fv/xC+SaJvCnrzg7RT6II
u2pwCE6M2eBvglvyiXe98bM4yiz2CqyIsTbJcO1v0x2ZG6eaSDtNcyW9tngHdmro+UT63rGAsJ7+
Yc/Eiv7rhgG783fJ54pCWJyrEDQIK1LCCTenZqKQbrFa1hskAAAJOnd/VDsE2RtXcYxjAq6v8Rre
74D96EGVD9nec/v0o8rEcVWuvOT7widGdZz1BTJrniuav/1KBjf7D8TvwSHEXv+s7+BQvFSiRtkx
j5oNbAsLn2fWHuJSofQ1/lp5j/L1fTWhpGtLiZpHOv+n3T6OZnxb/N4+HkkzuWeeljf8+VhkCEXX
X7vAiBybIlRdINnEFZ2JIQJU7ILHvmfQ9erjmOiSI0kraaGhHT/zRfOLCiaFi+SiWeCtFShdi1Vm
wpWZC777/MATt7MFdRhAZwt6L9Yu8M+Q0RVXlV8wYxgLXPUJBMcu2UNySt57VkkPX8NJF1kd88El
GMjBrQ4aO7F4IqanyhSWkZQ6z51Ilx/yxFFmyaUzpuWkdjc6ZAw1m0njmpw7AqOO8nbzxPHxAQkG
dGBe8BLkldWVvJmQkBnm6K5WNW8DhkOiXOfHVtuH2ZE8ooAfe/cgg74rOsoDLerCjnTccretf/Ml
jHI5Jt8X5ZbbgP5ymSwOxCT72G2lFVc5hPGH+AbtVjmC4XyzGiz6a7cw4DaZNktvwKHzVMAJO61T
cHrRNQsz2TXl5gY8CvNF/shUUFO4oG5dAlYettJvwqRjsbD46RyZoOUJtvYZuqfJDvQXgzNt7E0V
56+uBdvlLXbM+CrouIg+Qkj1KA6bqazVriRENcgmhonW9QYLrhwEFPUjOijOmnzafdcfeXgOAS7B
BBdC8uF6xE6K58mRAi0R0OqFg8iQT0M8sqD2Bgzci9bcxUuis299HQPi3o3/xzB4tMMDqKQoldYZ
0vT7bga90lPPkLRxrigsGWwALOVVYuJKX/NtkvJQWtUdPOVWmI7PkZhQaxNoNVrho2Rea10coRDT
OFEO+F2fD8FW1tCnWBxScbIaFyY7BzKc5ke81HA0nlFnUvW4AxbR60/fpTxaptsK+DdcPrELOOa5
nYTWBOOeaAtqi0IGHneIxPpvIJzmEorxU3uS1n2KAmwthueBGWlqDoQcBYB/UmPmq6JKwf9P2WkE
WmLSdBxJlgWQXP4Va12iagjjnXTySEUyQuvxQUovdWdSixR1H4Ucw/9WNPa9ept5Gie3RUisihZC
PZPM9eZ27lrqKUkkVXqJYo7ntwWZLwUWPLPbiR1Wwa8Wpd9EyeVB7lfieppPXpySfrn6ZGdq1E5l
v9V2IGMVDWjMJ+5+3aSBssS0PG/vCDc8Wwe72oHcNfCfAZPJpYGyX8Jz0A4M9mZYEFzOZ4A4S96h
ECiXCPvrMYvMEEJZqtL0GthlYF/s1RVQ+pId/0moGW6o2EiKuLcWIrZytfExIMlbwjcJGY7Nf9fX
h4xfOgdLwfch6VY32dycqdrUD8xoagYr32CxdZvAJr5IPPuhXvuFf3uIDECDcz/gAWA+a3iGiTJ0
uetl7Xr0HmTnehcpn/9c7b+V1uv0iwVhWMDqAenslfvlmI6X1fTbbHrx3ZlxBJ6Yr2oKZxqs6Y+0
+SYrYwnkA5SeG7NIbLEjEe70DYRLjm3gsNeuDUp/YBOppl0HQpTCGoHRduHdPr7OLSLSJGjvvhdI
37L5XEkiiwxHM1PZgUps/+Y7pfibcPdZjMJSnmEpuJTlOmvwZr9yHmPmS9zNpmdVJ5maieadndVg
cqc0RbDSO0CMmxhRaXsci5F9wIljF4VvAYLI2ok6mqYtd+5vwiEEcRrVBmNXWIvCwYgFkEGv+aEZ
WlTLfXMpHI8pNxUVT/vMTaDBoQOzzcpLEcKzMKmFLLV1TLX27nSlMB2dO7ehqJlrqs2RqOMa0LAj
VkI77b5Kx0fHX4Q290kaqyHOuCsmZiPCHVRT0NdJuw3ttSIFBHYh2/shEjl6Fold91j9G63KfZjA
yAVKo4CS2Bkk3mRpbQAdaipLzpXEP9EP2EEd7KNe2qOKrVVjXKCATBwiZsCHXuU4J8zAs1iPuZcA
Ij0XRD7VmryVRo+q49lhq0row5xjQrMGOxTl2fniKZqIpxiQEHlavcEvT1sQsCTDIwueBuGF939j
dAdH/P6iHUAoWyHVjfBu36oHGsto/DbCmJs5oy1juVhNjesFXfPmz0pD70FFoM/qqOEAQknZtZab
A74pVX6yif0qKjtYPPfmSGLfCnyUO7JSL5AOwchmfTn6EOJg9r/gTE3Mk96RjRDqdf9R0FQoRVVp
sJuqWj1E6TYLZojngohOq8XJXdpbZIgZpqa4USWnDUN0ar2tEU/UvCXhrxa5CkR0evD3mk6OKN0J
VEgw+tuj99JlU6vYpHb5A8VHavYRrOScDRUn+Fzasvu/QCrAMoTWMZwUSfmESsZ3N+U54PFTfSA7
ceh+9NE3AD3Zm/fJUwBNON2oHDq7hlrFK+Sf1+7gXfR5fg1oMhkbzfHxsARA5/6+huAipTSKHpR9
cxn4FZVVltJqDh8JMX91rrpdgNxg1KX7sSXmlnzbpQNoz1IPT28gdHg+9Y8v2ggu8up9d3Z1fPpX
BQq65kCBgy2KSo8VlK2LXqlYHo8PSqYsnqGTGdUrrZ5LRWdHQRw0Z9xRtqHK5dX+P35BTuGgfLpt
TeVLgTrTlr0CJDj05SZhYpVrtAMs7WZQxG9nOCN404OTQz6pj3h/muLAtVYqGOkp7znxlK49KDqp
favWA4CqqFH8DJOzI+G5hI9mDpN7F48PJDW2hUHfyRM1bURCStk5b/J2jGMHcL7txVxPAo6B7c1T
IxH2W+qCS9d4YLiAGQIfOU3zsVGilaVQePSa2QKFM8vhA2o/AdOuJn5aOX++JzuswwL2ViC8t9fT
Y25pv4y3KdWBDZgFqHUv26geC6zBEsGHTTO4y8uflbrSPjP5LTKWfn152wW+D4q1ewKWm32+HikO
mGWccF+NBlcGjKNfWPXQgHPtuxysiyF89raYDnyRIa249IaLjFwsYDQStRkjnN1hHtWtheDbG3QW
C9HviiysywWhSNPguBggqFzF+2wkBowi3MyAVmSeJR+bzsGjuwbldhrSAfv+ySBd3bWFI3sf9AbV
btL89lMeI4oLAtw4QITuJ3Rea2M50mUyN8RFTgrh8B3cCXH6Dl64447BKJXQHeUs9eUT2rgmfOLJ
I/Wb6yFeVER1eVElG1Sh3YIBpmyiqLFLvHdFMG+TWmJLksQm5L5kB1XVVoOB+ZJ/8bblqYJlh3Tl
G9NCspd/LVP7UlkoiMk0yGsiBvakeNLBUAiYqDvn9VlzOaOgTmpMXveip8H5s5zCxr/b0Ax2LlT+
3XRBAWQQHtIu/dB5AsJJCAzdIWUws0mFFZn4+2qodtI7EvtcDJ37ZjViW2w4anSyy3WOqsYycdVZ
ZnH+TpgLEjRDl4RADmq2sORXzvGTKS98gT8Jn0ACjR+pD7SBzlhuxkPODNMQA2oDdS755gCqxTWe
XIxwBiPkKeYlSE6Zsebg5afoPB2fL0RozfOIzVHMj8RpB2KbR0pHc+vy/yab/8JBkz+HMwB0b4ET
oku2QJ3bZ5aCMshyaZSC48GT4gTeygh1OzVBONTNNFUi/QJqIZaSXRySgiNYTyuOqJ/D7XeRjqrR
X4Yu54sKOG7gdUZ1IPSH32856zr+0WoNzHwXB/ZfOYy/H6m5sQIkw6Nz3aEkO19ZEMAFg503T9JK
USoKP1Zu3auEcEe4+ovYqkNyCNu0hOhPPT/57Yw70qspI8NMtVeRIKNmGj3/wvfGcEg/uB1BaH8+
j8W9L3GBSC0Kv0xjYHA15hE3HVesE9YFmSvrqu6WnAL4Xefub0hTMWzo4lxqLWLASShbYQTxDfYZ
/oicP4Id7KlO1WTNXeLDf1jAIRMN91azwCvDMRIL4ALU9I+rI+L6x6DV5gs4RPtOfR/2F4dYveyd
0htuZoEO4C3KpMS0FemQG7zg4imx0LkeqWGbvbBDAmTmHOZpy3B7he2K/y3kdb8R7ZMTi97srQxI
og5I2HyPf/hRaB660rAVnI39DRkYeUKYdQ2wZhq+A+sZYFNXvpKR1GhNlOu6/PZWu7aUmsuX1sdD
aCR9ngJT7Ocj3k/2XZpWZoDpQRHTUClkcrmWBqGn6AtZdhic5Gj6ZfQ1RFJVtkvkO0B2fvShs23C
U0wQceLj/QmysyY3CoPnuApb4WDDeoKlh5eVNGKrT3hXcEmEOxGFhtp9i57S+1W+3giwVHRgsI+n
eEJ3zYKIha8Vvov3AgeFGK2b1kGTOUeRL9K0V6WFZmLkheJiitDpn2muLoGO/6+Z9qK8699Nl8rw
VUoROoL9JBeqJ9Qyp4WOkF3IyIzTIBJXbcGT6I4cWT/ti+kXCYIVeBDbDLWlpU2IY9Cer+QV22Oj
ZXdt5B7iAr+n0GaSriNHFnt7JQRr56sglaaiCRZgJPixduF+ruUuWtYPHKN4IhiOCnOlye7+7EWd
vm/BlbTZ4x0QQGUdtvYyc6YUyO1lQhWdfpgXvAJhyZeE78qQre5i3L6Xo38B5T5hZmRFN/RFs1Pz
VNcDP5EzzB3yTdBtJY+eORGVrANiWV+zF5A6x2lCep1Ik8sjJS90FinH9yrSq8lmuhc9xSJtrbKo
gACOerYDa5oAdVj9xGwy3sjTYaAQtP0xUA2/UTyNvFpDUhSSTcCUgwI2MgW+OnxJP4DtwwbjJuep
XHlskz2lzvF9iNcZFs9HgkOqFPIvi95HcDaJ//6O6oLEVxhnSJVkB+TsYTYdKaIdJlsWM3tM/Iln
kWYI5M19u3AiHakFneAC5bURcGxHipm92YRVWvgDdsScADwIraKkwKJ3m48bDpYvZhMcyDq9GbpU
IqotEozObqfQuf80mSAs/aFyMDZOIUfKcf0by2k4uZSLUROhIbstzpRMX0z4DhOVpJip76Rgkc+m
WJftSMF4gW+Zkf/hts0Y1qB9wPtXXhxGrkRhRgNcyVO/qvA/zXY8vPcaTLL5qfB8LiboqPUKltwl
366EFn7oD5sexkKpP7EKpfBhvb1MJnBKlrDQ12RS7+pC3l6PSRBOtz/us03nhT8dRu3U62nc5Dzk
2V2EV97aavNuYRCjYE4W2cP1PwNlV1rpPhfkFKxjM311c7WrsPTla2tmvOQJtrXDY992vH1AZcSs
qze9632m50sqCV/r/cskGKfIgw3IBTYrmSLSBHw5PRafGKdHhNn6B55OSsQaqIvF27TdUdv+5aoC
hIEhX/005b/JPHdcseGcFc03eTYSn9J157XL296VFGY1rhg6f+x+H6bcjHei8UKdRBYcJD4l033e
oHldyw87hOb6BPOZy5SNwyNNeniTHiF8ujR14feY9+LiAmmY6JCfihP0X+DsLKNKZXh/iVz8FTMQ
bs6tYK/DH6pNds5/TeEZ9J7I1R0N94FtG4DKw/zEyLw6zVg66A0HG70Fj477xYpNKXRz888M22SW
nwaeRjjinI0W7SzKASGnFyKlq5I3poYiYDs8wr+9GgScg9FraLBqxtSuyitDXFEJ8vl/asRkdwhz
+XMiyqrkliLJ44vMaS5DB3cRZCXM67IIXi6SRHC0Ik26fcAlDW/kCjkZ8dM6kG1PKWcgXTs2xlIn
4V69vjxNB2sxJLLQPW48STnDhsOdFN4Xc4pd6+yqIEw0Boi0sc+7kULW/XRtGMoOTHgvlygSw3yS
Z5gcY8ZlzJQYoSGrsDnX2+vA0kVs3v8j9y5jA7MFf/UJj5uFz+h2vvQeedttys9JjiT/EcA2DJik
CcALqA3VGB55x+y4JWQS1o4BXWHeFSVulV8pGuSZPSgWm4lgoCmwoN5Vc8rwgnptO8dR+LN6eR6V
tJM8Rm3Pjg4bmGin9dRex3H2TtkcfmcjZcntsRhgFYhA0niSGTAt5RsQVurDH1KxErLERU/6i0xz
hpQL3rp2dOQY0GiUSQm5lQqr1yqeCGwRRsJ2t0eKylH3/IRapUnI6asIabLlspoKvC6Nhgg8yYEI
NN2kDJ5u3qJoMcIjrPr3JuR6TfWMUTALTWfVYTmRij2gS2GUtECKLESBPJjYM5niqvwizEoV75Fi
jR4nVwLga3SrTbEkeR6Pn0jjSK2VIlIoQtJ0TihsKZCfZBqWCw0mIyms6cluTLdx2lq/QvJW8Bka
wvTSKztzcmtXZBdd0RTdvWB8Hp9MhjMyLtFKOsB0PVBSn33POvNLQQWMIzLAy56B+PQoGH8owXOG
PXRjN67FiAXZuLwQfI+8DaMw3ablkAMuvCgs+TlEUrYky+uKzRwKFdvAKBpmkxV/3znQv/vSWnKv
E3Ta9w9lo7Wph7WovNdo0vBPNZMTOCwF3G1LW6Wk/887npFbBsX5C8LrIS2FhKzM9fIw3LAgAWuH
Mgj7GW1FkEdnWJjpSmhlmCl/g2H7KsLv81z7S9KfCPzqKsTxfv7LuiEkIjS+JOUeu2xoZ4bTUG3J
iV0UmLBiA4jde9EREpvBM3a2qgcrJq4E40U/i3Qv7T+d/hoFzS3gHBJTgHE0ahCYJYhxMyxsAO5v
M1TXU+iRr/rgM09VWwk1rt1KhCb/BPlO/x95iGm3u9vBsf3lNjfs2n/Y++yzOScHaE/c2QrssOz0
1m+xaNQn/X2BJ9mOGQGk6DvcziBXhG6oPwokrpwbVWKhuG6WQyE6csYoOFNNDR8DZeJrc3cKb6ly
GBXnKuJzg7Xn+DYzt00um88bZueO/u9ERLYF7RDSvChuT8ww/CQ/UCpgGDp7VOxOZ+YsYxtR0A8U
zUt8EjvR2nXUNUHsxedG1qr2fQJDiEHTj3cvbZMfp54/hwa4ZaC05cVrM02tC6xy52DewGmD7ojo
5v01PQ9WHmv+/QXV/P042WVznYK77u/M6oyKI/k5itVmiY1iXglKVLU+uh9l70hsXsugXVMVOmlz
MT7HARa7mYj4gdGGS+8AYw93ecZ9XfTwcRFDnuxiib3FPId+tL4uROu8Z7S554ojm8BZxTvLtHCU
9qNxVxtrZ+QPNwxJOCniv0dLE+r1Ym0YHFMXIM37LusW1elvjUICGa9X2f55x+ZW7i1JRZs+IfHx
M8PuG84cnk801kT3/i3TNBENDNIzYQLUXiivhm4NaKxAXVJ/ESlz6aPbRyOr9grgIGMjw4jpWmBR
QcXq2oFOwuilrAePU8724QC95zvOzE8vvCNWZk19tpolog8Rg//zb3bVoc6X4s7wMPI8Ss3oJ2lO
j/Qfssb7fBti0CdcUnlI29TM6JANpXvh0CQT/YS5Hl8m14nAD4aJg6sI0pxmorqx/wMCZwE8Z8Nk
qKiC9lYclLGvdRi0z5BXmL08sn7d+AE4BRTBUAQbBzwlvIuL8Mg5RYxK+hYeJ8cyjyQfIkRTKqPA
8ZEZGjnL8DLmWRF1k4RXejNBZz6wx+ts9pLIUcY5ppUl0q4CxZsRAmsTNL9OzKSE39rV9lI7/24q
EWLxjfZgk+0cpVwCWrj67bizj6YatoKLBrgLzKF9oi2j8xNSQOE4az7N3mITB6WHNT+SVzH6u/da
60bbaBU4YbbUoKoFOuOqJ1BvXF5OdLTUGYBHCwMdKbjRhbrp8XMj31TAyTf8VhsvDsWn6JpZnL2l
Lw7UbGHKy/6XOLOwG+sXCtvcFxmtipWEfanczJekDlTKLZ1NpXSGUIFyHr8E9rnqE6OnFJJYJGQ0
+0UpRAKmcL841+brdyLL7zQzhlR5JkCZJyMBHGv/leimCP7d7xnMsUUbQTRLFNVE1zVBW7Gvno/1
KV0HvhKYxIb6WLRpDr4R4h9smRUmbOdlf9zEMm3H85UCddmfHI8Kt7HBQXaBF+IQE9GaYWiQ4UjL
bV9oNSHoW73Ir3L2Ew6D09YUBlZRENCGfKK9BRP/hcruCl/Tmd1KP9RoFCG4fpZ/ae5r3/6IM0nE
pKIobXSqHnCdkm8Zru9VIuZ3//u5JYbcwYd2Kweg2CmBbJbQfGSrtXmDJ2Gv9XQwe5rt3R/tdBTI
16xSyMn/YVpKtn9GgooQMmgo8cIoDFUj1wOQC3OUI5N7KXYKf7n3ZJfGWRYfe6waMmckj3TXIbgT
3UZj5iRS+JTXBZx9aMU/MLNqI09UTARtjeSGUDwPooiS5eiqDEPJBioQ4ucXSxIVuyH+lBNZ6VMT
u9GOaAEaY1mg0ZF6c3bBro4HA1UhTgWvMMPuCJOrfyf2vC063KSZEjqgR/BOtjtwzWl2AVh7AVn9
IbVgQj6o8D6FgsXNfN5hUMbuJ9xtX9CL5gXzXZAEu+m++HV7Qh0Atu1gC8XlQjdC1cGnIxYrnT+o
8b6URzmaJCcwY7p8KNhWLXCQQYaKAD/fsObeOroe5l2UjAaLCA37pjCAQQR9GrU1IxXE/gZ1XDr3
uadcU5UBOl/t6e4dLcExTYBTba8iGbT3F69E3GE1VOth2YnWdYrra1cKKCjrhzegvKHaUx5R/N+x
t6rINl3SWhztrIqmZrzgjdeLjU28nWbZc98pik+HoC9+So4efzNbwv5FG+q41rbnE7bqpN2Hd5YJ
XWb6IzBbRvoKc0FsGaeA3ukuSs6qVdhBfa7II0x3p9vMxabYjTc8GzBYLH/SfbBn4KI9wquVjeD6
maaJdirvXtGpMlmC4zpGrVZbz13SRVfim4MDjnIlep2pZngnI7tZDoi/woumAgGlzBitOpTTuQtE
rELtTqK7qDYxgmFYXX0CUIejMf6QF2wU4BKBMSLCJ0kAvS3MQZ58MdbQpOcscWdyg03sfBJ1+U33
uLuwM1W0fzF+e3p54F67xF7fwy4R0QSWEBUZ9mAaZFvhSmDQneKOu+NjSaFo2wEjD0X+/5I1uFsA
Vwnx5UblgAPEjezgsuicHouBtz4LFERghMnDZSopP7J3vMhqVNDgVa55T6YD4dFd9YNR6msUlQr+
/DTFQJOH9Hx1He05Ihi8CnWBPhe0+b5sAea6dJT7YgzhIP5lyf0IeTo3RwOW9JPfz0mv5b+2rYfG
4Rh6k7Rl/srVDnngbrLXa6D7Xs71cuQbNrw0TZfmse079Qc2trEph2FA4tH0IKnPa98767xpGoZ8
vHsh5IIE1PQTGr4XSVifvOFACxOMEeg4LaKlY9LhhzHjGPo6hhTxDXWvHxYJwoC4rJzVrQMW7TYJ
AIGQ9O+FlH0LmhLasf6znsqvXgJpQiHuNOTiX3OBBVW5jcp3c35Tbs8uKlZ5DoNXAIdVPGxvtqqV
JeVkd/+WK7+fakZX4uWwDr881gd/2SFAcMC/GL9/9WhRkYSluoFh10xtILCtq05WC3qCVGXHALKe
zdwEnG2olySE/bweLV3XrNB0tX6v+p74xSnCcdsJGPc7x4dwwDILyXf/TY40datTcSWMiEkUpowi
bWPIcH3MCD+MC/G9wmErAfwj6aJpCKloqYho4ujZAHJ7UVUrIjVnQGaBWIRkSmK/up8GgqWZEp/B
eK/0Yae1EdBpe8wPBoRgGl1/JkKnxbHNq/T9husnvEZh8TFms+E56ieEsRHg/SOnJjmcREjMD1WM
t1ITDxHuAGTOW3853nG0ySZot3/4jTGRzTHtlD7swWzxIFPiNvxC3/5w6duFM4SVSSTa7N256KyC
v857oebg2zH48Q2pKPx5f/eFiZJhjzorPa1zuA7DRC3r4ueNhGJMoVRJyU9xuCIuyqi4Vij8Vk7F
FE/yUsUrUcYyr6ijMo2wcfYZHpYpTjNU05WtlWgoFXeSlHeGzFjYQEa3c1d+IDykDBSMI+NLo8OO
DoVFLTb8AXwU3VjdHAYnvZfWQ+RVDeCGAw5Hx+KJW2j70DuqlSPEiKDNMepaT3ISYls1I3eAVxfq
s9183L38ek539Ig+U34ZWAfzc+8aZmFYfhyHu17bMniKU06DX4bxilBQaARVNoREVszsaqJdujOQ
8O//S1RLreTUigY5Fc7RI3QtOg1gCtZBRg1iV+eXTzoXDW0tpfgSb06MgD17smZ44jcyrJ+LFOra
1BLCPOWY6OmSawBh+Iv2WvGoWgPu3QUMcakpM7Usue5aqlAKitCPfMrs8hPLMF+GIShGXBC5n/n8
kK0AIHKlgXj4NhR9ktFwYkO2escSVTzuGqTSF6VQO35rmJ1S8fx2YUyHAVpfsI9Po1ZJHL3ffV3G
eUK3e4N20WvK5f0yGCJBpWQ8DaPbg9ThnunSW913obND0ROYY+yYYfkrEP5rIOh/S9dnb4tq4oir
0CNDqdZ1F4K/4FUprsB5bc+IbvhBT0ObEjAfqFeG8J/U3TZ659IcIAWkPnPnR46WdClNwQdPARJM
U9X5H+e9iJCnbE1KMwD4EO6fSvLTh8S03dCFJwdt1yRAUd47ZyhZMrnSCOPQVEA3ydpnmN+eZxYs
iAVMn/Isx3kyu8rxBr2w92INTFAPJdjs/ZF7HDnwwAWsDIeDj3/6VZJakNbY+FwTp/p90KArYd6A
HOK0ZiSpkK+B4AoZ9M+9LWT/2xcYAUEQ1gX1HQTjgaCGgRxPCg46BTGLbVF1rh5JMA9Qv8Zhswi0
TYlZuD6Gfz/k8v+NzT0FI826+gPhCb/a4TMQUTb4wo55bC3Fqr7wQjyylPK2QPW40UAn0eziRmus
Y8sHYAq8RxubO9IKby0kxPC7VvqQ5xYker8X8wpCA8lJaxuB9luJEdRGEN7QnnWZcFZalyR6W3bg
l4c7j1WeOUSaj3JYyR4XKry6avMlGpnPOLk8/V+CCkvxvjJhG/xSr3moNsDOYobsY8iNWOND7rrt
fmE4fNjp8pFh56twrffkeccw0UALG6v8o7Nbd0aRaTEXcMPXEMwRjhCWkHGyWLOdyj46mbzMRoRk
yUXHEXpJs9Y6HQS7m6+C4FlGdMBGQ8RQn+4Y88wQ+U2bZD+AvCn1fXg51zskL23nxWoGunPRZqzT
15EKZH2YBHIaPIMMzrVdzlL4KlE2gA/eHVW6x8jcRxisnTVcHEf4zk2z8iQhxM90KPHovUX7SVe9
JHrOcefphfZrRQMQvLcDYAJfZKL7yUrvD15K8ObeKLXnkzDAIYHur4+vFYGwr8oR0aj531l3M9Xz
MPWWXHJSgWm44Dx61qXkH6Vl2hYoN0/PImB7WQgx6lEcPGQgUcvcXB8inSihhb+twpHSmhrZh7sc
NX85q6YmAJ5dyosWlBUfvvASxuCDaIIXIcgx9tOCJz8EUzzhcLp1kWsNtaSbxKsP53i9OBckQ/e9
poqaLB/OO4yD2/eKPhCssMznFYUkvmbLaequ7Ttb3I/uWxX2TljP7jB+rZadMzo6Zas65oujfsqT
HWDlSvsSh6CLJZ1kZ+TpPDHN+x6B4J1YnjIq7WgieaXSFpxm3BnCvyPR1mod/MYXvgISYT+CMf9Y
RCcSCgVaFY9qlp4VHjtqlxuSEkZIK7SirBrSqIqDp+Vg0XH04m9Gi5RNu2EQNd5PGY4uhI30Cdox
4aQZsqTjnTMzxYyqgxe7P4mExOvAXbWXW9SjvpKuypUdJJ3UCbFU9N/VE5ppvn/61iZ8GOR4aTEx
2lnug15I/DiuDlRofVtQtnKrgIqUasSOpXncBQHL7KpxirMQJc10EQbMhIC5qHLLB3tNaFriihHu
+k7IEJRQsd9BDppWI7LFajE+5N1KjcxG9zbvV/kG1oKXNGJhzdjOi+IS7fxn6OKYBed9hEL3pBhq
x7XL77Ix9ibMiksMfORpu4FA5ovP7KTnvcje/xEuRTww/80iKVMgm/CFcq1DBZ6niiUEWALjrS/H
56vHj59AHDvGcfwmyfXcmI2kUqGWGv+0eWwT9Aur+7h7vR8VipNrfCO4A71WTNO4UvRgoEG00a8P
NM+eKM4WiZV9o3/ymJcstq+aFWPwZlt4ZRYMjgNOLzbBY+5jEZ0VlA15sQB+nDbwdZGj80Y6XG5F
qFjmw7nP43lFE+7sDbJEeqKNjbG5djVVr3ZL2YiGLI0xifYoDVQwC48Ket/fLRfU5LYZjU0Gm3dH
srG/7jp1H0xn9BX4NiaE2Fm5JWM4tFrZM8r3DRYcrl0c6nuGEgIKpPKuHc349+35M+KINSbK43Xe
2svETNJHYsU8CnHitGuOKKWhdtAd52EYX67ymesqbyeqTnRe6S9RpSCq5KrsnFatFTvHRdmI8sjT
HQBM5+Kva7tZcNwn/RR2lDuD2cyqdMR7TtJi6Oy/+HYtq8cS07e3IeF/xeZ7amONGce3bIJxObLU
AyJ3W587M1y/QzgqJelSJ5rpDQ5WjaaZQhEcmgCQLIksS/en9PI44fOGAYiETKkH07uM4KQOQcug
Nqdqnhg4xAKajXVEuyAuXhBSnDVwtesq0cqo1sKGSUS9L0EL5DUawMY5yOZfmbL5BtUbTcEN6wRT
HXym+FnrAh/vbxMRoIaH1F5bfmfay1D9vJ0+Jjek8k16xDUcjBC0FTeYtphBjkW/zbcFrm2sU76F
izuRRBDFo2DTI1BFnnrg3P870Sf8Mtb54TOkLppq0dvnrGwin+KyrwOzEiVb51wCPTtH3XqKA22l
ErmGNSfz2VkilGCQ9c+BU+CAvtwAIRJ2zISPu24j6F/nP/QVvbusVysGU49AthieW6ESi7zbqh0D
XqZsUVO7oXtLrHcF9BqDrR5sJt0NuprkpsQMPKAB1cf4GvLpEXA9WULirtAiUeKiv9oCLMLbIJ6E
5eVinWlgpqzbwpsiLjhSiuSrexTeLtoTI/5f6wcJHmyu6WQysPdOE8o2IEzI8YFG+1RcrCqmVSIS
vXHkCbJyflnpnpFibm1p9qRsBJueE6os95Qj6UKDwnCH4KGYYd4Mdr2OTVevhk/+0Q38u2Z/aGnN
tlludpPEMIpRQXa2wa44nAFmnuFTRNXHtHFBDflcNwoj4fsXec1zS9HXXUpaX55UBnhGu1HCEaXJ
Ci0HJNpFEPYIjP11s5s0//LEjukIZqLmmBAEb596vjrvPAw4t6lHrBOnA8iLMQawj+QrrRyYq+aK
9WCvSvg89eVKDHtxD5ThZnt9mYHcgQPPSGKa/NwGQ/h8rmZefDjcHZved5Ixw/5vklBPeUfgoJH7
1dVJyyWLbu3Pqwr7UWhGaNlAs3ArsKpFjpgJNrJFgsLig4HF6g0ss+0GbnOSvhrWiwwVwquVCOgQ
vLQTzQDHZ5O1MLoBEdbG+zEgPJbRDMAZ40jqGNgtJEdW1G/gG8ING7CWblRni2++mZdOkDhtbFC6
uhnPqVxDlJpYNioUmOH1s3PuBoT58/3k960jQ3mKvvHpWzwDLm6cUnvmuQ054/Vbd12Fe2TETQs8
JVAseCm56joGK6YwxJAwdRK4ORByWvgWyA6Ggf928VIWtm/uig6xOJKJ1r05plDd+mYNDQJkaxe7
IvPLULdeuF+pu1KOpnMxNEO05qJSIAyXsE6a3NdGmBBr1nyGoBBxWlBEihL14m3hcHzOLgcN97AC
l14/w/xKuGplKaAV2nrLwD1IcRddG057//UwCU3uQFzYN2N1E0hJVLe6p/WB+E/k1nWxn/Cr/2nZ
1/SXlANyLB5uVgfOdd1WfXERLbgnckmrwtlIIiCi58nh0JiPY+FjCqE1tSWQVkUvjn8ISHDgCWRP
LGoto2dzxNQr/nU3CCuohpzDXf1WHviCE9TkmLEYNslNNOL3P0rPBkAB578Pv6ROtprSRejADAMF
Fep0+pDDrSx6znIRO7+zqn54xeSTczSJP8YsX9AJ0E2GuZfAQiGCEwuEhk97zYLDMpG9/R9yCfIO
3xbIQiEoGaLqfyDcLxwBf6H9FJhhgq6/KLyTKAmPLL2pMA1WbPU/uyKVcZW/TDGY9qfUqXwLhS3b
gkfnQpaKt8he7/PUMkV8chLvwcELJby31IE6sGzPftb2rBhnM6NayEh+R5doAEexGmkpQfNbbTiV
/xjmA0m7spg7IpBUCY8CVBCnAdgPI3WJeE6ksgZP2b6c9IsL6XoFei3id+XZ6W579QNQfXDddXP6
O6chTQRWaLDxEppsmpiMDexQEeWg/G/ua5y3+LGsrJaIxR4isxDcznyE7+hMiHzX5tPuoazc/q3M
mgRDv+i98H1rFK5lb9jYpuzxFrRI+CIjccMnjDrOMwFDFjJHUykwkao4ehpCugWM2Tu+Sr0RU9As
nXDFaWxU7tnpGRHcaeJ+lJg/opeGinfqz6l96yk5oMcTuYG7vbn9bVl1Yope9btWx/sl5ilW39Kr
NlambKGnUti0dqVBVLhHlcKEQIFoVf8FfQA+GRD3KVlYvxn9K9u7VlCrDXdxQ8V//8DPXDPaPuUL
iRCKM2uB5wkP0KsaTEYO8pQ8ok8Yh2BuhH5Fbx6t5mNmSyQTNlrEkWH9787fNrqfh6abY7NaOhJ9
5pq0mVLbNrQ1gJ6okifU4lumKbbc8NnKnX3KCbKQgYfXZRCwY/tHA1lcirN2XpZiDXnpvc2NhXMO
aNCxZu6aG+OFjI0053RinN2lgIjg/gHFtErn+ZqqhMI/wxuKmnYnFvAXcL8y8EuD4kFAdeG4/hAj
Ams7+OQDOVi7Mh1kWaENaUSCWHvBBCacLqpJ9FG4OMUtptx8feo1dtdDeafkIet5A6ycGTyjElQM
+z5psq570ayvlE6zl7Cp1zkUW3rIQjrcUAVd21igd961qJcfhzPr/5qjGWMZj0NprSUgLeFGbFxW
FxHWrVga8XWvBrWcOLUjnKGYX8cymB6VGp5LqtqUzEb7CZ34uY4zgugV0tspuH/Ps4hhH61gAl65
0sEw9JDoQ4fNPaZPSCH7e8jTOXAz+5Gn+OIU+V2RZofoF/a3LD5IXpTLVwGdslG+yf4/a2k/kLC6
X7MB8gbcOcRXy96wovcbtQY2+Z3pZ02nD6qj8Wy44w4jPywBtMDI0vQSbY7EdGNdwS0FtadyZS1A
W0SVtFSESyDCJUabFE3upj2nCJZ9UwqAaFa8BIms+h52umFxp1W4tRcRhxb9jBgPojl0DFYXVC0l
qhKzFBusZe+aTQcGkfk8la/1+TBKfpUugFua+NRASUEPXdBJ7tA5KrXms1swm+0J1Job7jf1aZgP
ZBGAXRsE4ngwcDBM1wdfeBCQpzAwquF6m6yfr2DEMq5MVzeWg9TjpXju8V7CmWURzrxe7YnI0DkT
HWfdEJ8waNSHWf1RF1L1kPO+32KoU7nDXG+pndMCzjkX/FZGli+2A57clyTgCKcccg/5NYSk1Q7N
AmF1OWKymk5WKyXTiydKnKKb6K2K/HH6ZOXE+xCwNnb4suIp+YAtDlBaA7MUDT0f6bCaec5eVLTz
NjM1IDgovBIoyWqXYIjdK0mP13hEpgt/DbALvNbolYA9mqBkUGYrZ53XsR2avXKsx6hve4StPU+i
O1TWhqka2Qm1hjuQM0N1bT/3ohxLXGBQh3AMDlZTwY/AkaosBlHKFoEzj+BpmJJbdBRR4ngek7/r
CoraWopD1fPvLiUoAppQf3DJVJq+on5yHzUEamB9GVftUo+7KEFM6i0TPsLWc8RxO1x1ishnsGz/
YjRbv6l6qkoIBpb0Bdjf4OuKNyHDm3QJNMO1sP8q7nieJtKK022VriNceSODHRUgZ9F2erYFjY+B
FBETfgo06ywiTjqp9uXYhZn2ebK8eE1nVxW2mMLJma5twCJMzV0Ttf50ngp2ZxPsvAPXsTDVu0Gp
mmVQ4L59I5Hpg6HnI1Jx6Z0fgmwbuncwH2gKq2rwBsJrQVed2O/GPF9fiANnkR5fzaVFcZhMNjxV
0Zrx4TTB1f6tMQY0ohFB+s0zBkGFM0SBsDoIdM+NoIU1Mj7abXQEGD41MwsCvJAZ1lP/tM5+GYSl
FrONnjKcOcC/rE6YvfTn2AZlCmZYkNAIznqG2vpMIjr5dPKLxybnqPEx+4CTlTUK9OdH9UIWHW38
QMdiiEgrCTTu2sGXu8aFFrIStjZPAuRRo6aR70GBYEAAVrOvHbDGkxkY3GlsLfqST6Y3M1SQK63n
0SDEZQe/X0rSBrmBn9GSmLSl27O553gRTksBV4hIlLrwIQPmN+1vFRCSkmkROj8SM3P8UphYXJNk
FEkRGavUp5KiBV4xWrvBENeYcrkIiowwuU5Tp/pZ72W4VNali5IrZNaeyAcLEigeKPgUPKKnjL04
zebLFOVf4Rl86RX+AVwqI3JbnROQpzVaHOy7XIpfqDGhKQgytC9WYTGTfPVJhZHYEvHbHCCudl+v
RNmfNhJP5pZ2vftfp/j4WZyR4r7AM1TJcdmGgMift6hhOC06lA+iz849POJKYN67N+0WZzDgctRL
trR8vgbreZXaC1EgXf33+0KQaTQ0AKSbnRSostpBgP4jKN6arBdJcMA622IcDapRsdbkppL7KU7C
88KF2MQAKWeLOBAgyQ2XkGp+iqphSILY+lUI7iklhmAmkwi9Lx1CLyxhLZ0N8YkBNBeU1IpH4d9z
IW5bhDRkc2/UpFhL2SiwIP7qA/Js+kKQgqB/B3+SbusILrbarUMLnOkMm4qG/RjIvIqnySuyOP1M
6aTzc+GwIBdGFtEIF0lytIWZN1ujJ+eKij+7+EXk03+9xpqjOVFthesCL10br0jpkkpbfvkm8z37
ymmxJEgUkoc7KFBqpNHFn7ZkmdXJhUVqE847jTqB5QP3lxIbwZTosT+/rmARYDZFrQ1z/5sCFmcD
iQ2Ork00CXVYo2/PSJrMAHLHTmTqYiSNK3x1GGIgJ0UzsL0Be7aG1mcsZ6NpS8BzL8SUU+oZFxe5
3279YfXuLFO6SdsfChUxEv8LXWVnZC4J+bnbpt9Wkd5gOZo0eh1DZdyZhaRMRUzALZ9Lu3I83keN
LfSPwqojxVWfhPC1Lo9JO6gMyCEPYsMO9jVOEVv5fvUNcSKw8lDJYMOcfNgytzkXzbLWXQZxqj7j
OpV9T7QpAePITPsETCghCE6N4jDf+jD6arGOSzsfdnghG9vJ3Y6lEcKwYaTMZAhp/LFojab0TlTf
Ta1Lat/hemSInjVm/xOW4vyNdpUQHoUObHqHIp9N/ogW+P9wCMVdDNHMBNooRKLtOXJTJs3VJHp6
cGLOGndhi51oU01BhW7QhjNFUD0kEVpNXWjhToUn04wmt11RX/+r2cj+acXwlvV6/wnxUY9D/GdI
L1cofq64Pgg6syswNSY0mdjlggmuAZdOoFcBTgr6uEabPmtSEJs4osGNABiDLB6FDb7bpnoQw6pl
dNOniFtiaPkvYi9yakpmAD5otlUVhEaa7xdfl0W5LOWogndj8ilHY4u40rUxQGva8rlpsC99PjMb
Dtw2MmwIi262H8s/8Mu0Da8lhZ2S+ITWCIC7daW7mJgeMiopS1r3jntDmsIegA1BVfqy0ts2n1+7
Q2vtWLCjn4dq6C3Vvtl3ddKrjY+ujxKwbGzEDF6zdCcS/x3NuB4pNopCWJnNg5ln65xcpwBiVHG9
PM6pDT6supwyfV4llQw9o3fCTXbL2ELgq0hAbbKTNh9qTpCdapqIHmzL04agr3/oWNUAHSeVu/zh
VLes+bEwe759spvXgmDf4lDBwUxG3JnqseUgSEcalrvdKyQ9dqr3IJC2U4XVhEuHtcKY0TdjRzzf
mNPhwzIjBlZ6aBMEmd434lUirogBnfTYu66ABXDbt/8pA4PcpvVwMuxH00wN3+SeEGRD9aOQfpUV
0xIGT88h7MINxCcUyFiaudUm1M3U9uzNZYMZevEVDKDa59PnHJOh5NStaIe+Dv8gaFLFx6eN1zmW
Fa3sYaETBlbTDUsv29BGJM8b7pWoJ2HUuyHGsOAc6OFjXFm2jjHLs3i4YmNUIFe66zwpnhCOAHyd
PCa86B2wjnQMCR2Z78OCqu+X56Xa6bOxSyabSQ8lX8M4G9NGi53DgXU7T8rsRMULh0Re78+ngiHH
aEinu/1w5NuptxfnLjkJMnhZ4DIJ7mAk/5sY2EC8wGSZu3/qqbpR8v31eQvUqOSKxHtY3KXgCM+a
IDsLIACFjw+7KkA4wuLU3tLeVTJ54meaSdJB48evcNN415y0yWRMC51GMUfUSlLZuhL5r7fT0Q3W
trPVuz9ifBa1qrv6OlyHDOhycX1vWbGMm8Lz6Lx3bjaMskgPr3O9WLdBeFuBY992x1ViBFmjXaBC
20vyJQjWvxuoiaR1WehsqPZZxPMTY61KqflNxwIeB3zexZFO2GfmcW/bjUgu3BeZlblXHQLfbclh
tnNTbYsli/U4s+G35uFFAmv2qdwvj+/rgK9byZyzLLkLUAWJU1FtZoCyThUztTxmy6vKj0miklFZ
IAVIhVgbM5431xX0Nmuy2BEuo1A24pvTg+CU0WflABiMyN9I83sO1udmOsIsiRdbrpAtyHo5lXam
hYsnRwMHJmMSHWLVzo5JsRR51E3mCJCqGS3UmBHR37uUu0jjq6L9kBoCpIvzDjGk+uf2VvhaJOhT
/lT/Hij2qbj7aUHXTiYPDsxe7jSp3mm105CjUC/yfLMFPhjJlPBR8f9e7TvHv9vCdec5wmxWmaHi
BqONNtH1CXH7eRiqrIjByFIdxQwr+RJZo9qUDptt9mtCsRCZZsiBi4zcwaAk2ZGspH+xZvU309UC
75v697TX04CNYJWiMAUJ+dnt9WhgAjb/tDZ54MPPBtP8VBiqFNp4bb3fGN5+VhIo8o9BQPBvqbXW
ti4fHTu4DuuRWqJvkGNSfm0m6RrjbfSXdomL+w2GnOzXx1nCG4WrhP+gT3tDLKMLNUogQxZ3dMqd
Dj3hH4BYJ4otTmfhbHIffq8fNCC9tjgsKaWSUHL5PesfEElb9orh2FXKlbLFitSn5bLwxK4lMZfo
waeehvUiRSNjv06oj7zURRr8fVqifzs5skl/BPF2DAAJce1QUeOyDw65Br+nGxXn36GKebcrTQy1
wsm3HEqS3S0z5zZpwiSzfHFGm96L4+kDSvJNB8gtv0rREHF6oxmUYVApTDbkGaWcgrppm4xdokO5
KN6XKGNTUNNwzRtaQejoFHRL86i1oTBx/RKz28wUtzQ4wcx1LQpRqRIMlSB7pz/euTfQR2NHw10P
msmggM+3CO0FHVoDlMEsET/KSYp+nL7ov85neKDYwq2y+nfRTkr+UM+Ck12S+tPh+NWXNsdNDcFY
8Z+siPWTGBJpuNCk5zp2QsezoUiWnvgvSdEHDppQB6h1Yb5rAUR56DlCksImTvVPPreM/WEGQOih
CLCcitPYDTqGwN+kOn5swCkKCisDgF6c4QZXMFDCXI7SC+YKfvBTkGGmwYFQ2ofYE6Pv/jeeKJp5
O1j7KgSvmn9MLiwuYEgM7O7N6S527FKHaX5krgfrsnvGuqvyXBa8ySzCd9l5fizaonqEewE918FX
EJfYnjTkC2D4lYprU5uZKVB/0dqAJqOF/4Owta/GtpdthUGyzSUNjgJ+5GFFQFpRGsGGOA+ZRPlu
CWq/rTpjZw6pR4L5PzdK+F261l3ZgDvowONgK+KpTtJu4hYE3tCugl/gvANAS2SekcLBQSVxvr1w
Tqd/NFkEUIM4s3320OcUahA4bgzlg/L2Up3H2e4V6i+POlV9pE++biPQh0WNXIGLiaNyD3LJQeYj
sLmiN3ftFHVqEWoy+ed5uNkInxD1IXzOnLkJCFD2QsDTfTIJ7NJE+zrqb9w1YrXAE1S1NlCjrbOC
C7uwevr9T+Vm7YASl3D7xd4qc/489d5Zh+mEZ3YJ/McGiK+gy3Uktfs2hilTdE0DdKU+rSlSM8qH
VyGC1fhH92W5XVp7atROUW1b5FT4nVyHp99LZbWq9X7M+Z9Jjm8LIWWvtrzdoDPOaPKtCwAXvkjU
YG0f6gqtnONcb95EdVOPI9fi7Sjt8eD/KQnmMZjHQspXGJu8td1MvXeLts5qJj1hQQBn3BSSTPCO
41CIay2aCW12f/HntadOuHBOzygunfTKgNtfeRGgqsF+5eMn0G1h2LHXHwYBaHmSr+cwu+6qtilZ
fxbz3KC8JDVD5cVnRQaH1N8CocojYGV5PZ3uNELqQryMuEITetuygfm7M8YegPm4c4WbtoyYQvfz
6zonp+kHsGx/lwX4DT8RVaA//8IFzDLut9A5GXdj3/0YZvkC3w1GOwE6QvS0AMOzgR3aEPad4mTE
QCPKXXLqmF/blFw0W47QjvNSYLHhEDW8R9CB51OQuN7zUQhQZz2dIGAVfUdN3awn4pICQeEXjkRc
AeZuHeujRK6nthque0EhDYpKmSKF+K9ga8H8GcrQlzN7VxIxMJTGTpyK5Gpm8o1RqBHA9h0bEX/m
QbYdmwS0GK0uqdYpKqeFPlwWusgaYyNaEu9sVFoFX2nvgqq1K9FvcVtAxPjDdBDnv+k1Nf3sipc2
/VGuXK2bR2Koh7REOa2r0M8N6yfxj/y0IJm+OyJG8NabPMlmxTS2KooibL7neng73P4aF3mnjk+9
Eyntu1yiR3+WRgUfP3Zg+OjmRK9RjEIijAKQ031Mrbb4ACC3njG/d8UWUORIrgnfonF4EbKzm5v7
WHuibN6/jQBe/Q2nEercxU8g8e8SyO+R5KDgH1JuXtxXcEXPqJajSHkcngl6wTvcLBMSLFrpWdn9
E+v6pU97iixHZ7zPIvwHHokkGceV8tERjWE31uoT8J7H3/Ye+R7GnZk4C18+QlwfQF3wmcYpvezf
SVKVnmUGb/73Gs0HMU/UY1p5ZlIyqrEWwtWWFEb1UA0xmICT5MKqXIRzLquzQdgDqFuWgfaCGCTf
y+XX+DBiOfuG5eiW2k0cnQOtQ2WfY3MjB0h83OaI5uMxjWQT6SY5WM4uJAuBSUC9RnXAoWyndIst
vTs92c4cSvdQUZ1lfD9iYfZ2ca4cBte+BEUxVf7T7NV8q3ztcISyK0DouqoI0ShNQmHYtM5b5ZE7
cBUEcuo7NcrT04Do9AoT+fzzJc1fxx6hlByltnNLlE5NeOybeHSbvBjk/iaZcmhsSjtDDOiS/HoX
ttJSkoRTujJ0R4VktdvDF9NOUOMfrg6ayJp81B88aCvrfduAc5e/qmxtIGanA9MyfengnLnchdgU
PmRX4nk+9SFEBih2+g+AO7TNGiJd+QudoNw6eAqAEa4/zbEKMGWkzS3gN+YpKzLn8OpHgEpNT3Rx
++QhaPD5OxLgfzj2wbCXYGyYMGXVVYFceIwPRXECmG3ZTME6wxhfNHRh+HiOQ9ly7CmIKbjULQpw
hZTfLnkxD05HElMqg74YwnNMkH9AAT4arPwnzc871C0ur258NYpD6s0dAwkXjTzduEMEiU1aR6F0
pqNOmV85RI/icCCpFzkupD2k8wcmtDC9wKE/IdCRB0KCRT5YstySbaQNAJvTH8kZpZ9Vea0T/IIM
lPjASN8jtUYDCwE7pCxsWYZR2PZYB2kara2tdfygfMY82RjGBte28w+GBIgfl0AzeWNqBqO3bK13
2/dA8P/icP7kcXwFf5eErmLEM0n3axNoDK9Z4f0d5YCO+412Y9ZB2FFXyEojbvDPBUbSnF5lnJis
awvOl5gsqcJCsm8w3POtTv6SzAxl18dkNViioT1unGJwBvxiylBDPhf75WNAk2fmuBboSRSguQUp
scI79duw1KNBQb5lxedQI1Dy9OUfJxel0WHMHbAAbgJmagC9LVSFw/lwF5Sytd74XfERvggbjhOh
V+o12gvMLT/psr9tpWosU2Z+VmgpiuHDFS/8Gb6/GEDELbJ7WGY8JSDW/+Xj2Psa1XnTHpQiOtX6
NTuttQl5UR7UZFYzYed9CMEeWRRkQtuTfb/ojKC5HUcbbbM7vszOHjZI2Xa9J68VdWvh4V378WYb
7TfaaknWeFi+GG7KZMK4nfY1dVCEt9klj2sKLNOyozuo3gvKB2xzPG8y/uD83obkrXeVwNj1FOSj
SHo8YK4+Re8sKrusElKtKGUfA3Cxx//8rb0ZPd27S8Or4EGCo2cIsF1/UPGwSKiJbzEXpGPu1pG5
0Lh94OAwu6QTGMnn7niLY6mrh3+Dq9hWNvqVZegm0VQyfkyficXZ+AYi0n+etgj4hnkGaoPiUpXA
8P7xB1VOzQOyRf2nvH2liuKnqfwqKNGiJQX2Md16xPl5xHzYLEq3f0E9/ndeUdZ5aYXOntmWw+wM
RTvvkrEBnD4WyaQy7IspC+jwYicbvvglCbi40C7Hd7m+d2Sum3KiBXqyZGPgd1B1LoKGE8btnKYf
uDff+Tmf3mCtTiOZdwZYfNSvNdF9jPMd+ND5+L2g6HfcVztlilSAyp1rOuI2qXPWlBixQTCwrLCA
6oimrnd9AFfmRM0Hvxcgv9pGCSdbcqVulAEaqnWONznWCGMdLRg0NaUciPCpp6SK7pOW3Gx3uf2f
8CkGX9RrHxadKIP9Nlv8k+cAhnpIJrNjDua6b94PY7Cgp++cdvXS1UeIOGf8d78zdNSu7fPP7unL
1KkAYrQT6Kt1DbaZZy0XGvopzTq9/I5ER1u8rcOw6eaXfLl5gZQypgnZznss9NSmQEsvilMv6zFi
eJYSEk9m/NDVki6UAoF2NnmKA+QYrdt0Cv3HzAP3RSEi3V2/AaYhza4JavF6N5I8MeDAm37+6+nx
TzxIR7NKZXST/xctmdkNDYBK758yfeQ0h7Rppgi9Tf67UKSBFnyM1vLoICQYsKq1iGEf1eAQM4Kb
9zornfQeO+ZdC8YcSwx6eIMzZlkVWNBnkZ5zSYEFZVTpaoUoR07Ai/3hHLGNIRKFemuukmmoR87i
2gmb2KSbeyZIyeym5Evf+LDfR0DVIehaAre+Tvpb9Vrda+1+I5OlNmzI3opkFKs3AC7G4qzRqce8
MfgGkaZTIt4vC31A7QsFZk1Y2d3PEFyDv5A+mMSNP4EyPW9gWfmPa/oXcovJwpzeYhPUXlAzWzbF
JtURZzCLJeh72P4J/uB7bhXqnNPDfZPkpX9ahUPOChpylh6LPa1dGis0aPMeD0d/cgTlKHtc7KfN
Lq7B61+zR0GHhQaabSYWoX/QsYZ5X9xOV+liglSKhtDlKMwdgDc7QVfn/lj+4jrEMDZmrQofDgKj
BGoBFKCj5AM5X0nKqUaOrQzBltfGO/ev+V3mtngKrxx4ySIyllidysoBD1VRwtsQlw8lOyCo25MI
Z8N6yl/bPEoFQdCdZuA3A0ysEQZ8zQC3ezo4dqwa06YPRXArw1zrlzlDgaG5k4FaOpvL8MK7F9R3
ehzFbumY4fCdvhtHUpYQB2280BufNvsgx+y+z1GtPrIjHAO6UbFuCHDxmU6NDr2b0IrV3l7Wat+p
HehEbB7E4tpR1++5EhqITg/+fWnuo79XbLOjcp/vID/0e0qSia8ZjfFi7QAKN55mzPyTBBP97J4f
t8LJp3LJkpLhhiXYCkHjr7mYJqwTpOoxy0LGyvT9Lvtyem9M0CP1yOPxlpU3QEsR73htoXIa4P5l
HKKKN/FXo5GSBCxOJlfH3YLvr7+qrej/l8LdYnZyC61weyz2ZgihxN9YBkaO4o0fldrFSMpK6Xc/
cJMGQMpkm+tJXKshOtzV3cgB2+2eySiZ3K8NAelzgQ2JIusqDr8DBRgBuvN69Fxf/SmJlL8tGzPB
+7Q8Y3jneaXig5LEaa+pBaYPwXbKDasTAoSVmZ4D6OOzJiJQ50AZZQvwrLw2puuf+QefL3YWo6k1
yJ1y3/L81Xkbp7LJOiSSkaKF9tkKLP47k8s9qTz6YBNyLbj/3/grOPKsHKcSXaaXscH2A3iLEr32
KiLcYzwb483yh+tfqsOHb+d9/n4DNZkj7XbptSbssFEj3fMiIRD8tbaGqk+u8fPPgK+UohXrRKdC
hJbF5k3STVbVSAX0vOplkGI/jHdbB00cw+y23I8h33bNvgxEotaXXtNOeaI8ikZxrlhUxisavWHB
0mDi6bLkFTyk3EgAS7iGBECK80+/KcysBOy55960FQyVBcA8tkT2M5APPd7qyBUgiHpQ9z9Jas8h
YEoqd4ZxRzSekthgONJ5T43n5Re+0ndqEY+DfKcBzPF6XGW86Pb5EE49Hv3iGDFAIgH8tNHXS9Th
zDBxAK+Y93XS8xr/2ER2dZKQSa79+5VdKKOim0LomIJVbHcj4/f60g3/NNJv7bYz96C0h4j69lpP
S+YF1fUObAJsk/B9pqjjpsUroVG+QFqtwxFe6H/xShBlKUjgst+gndc85c6Rw1UdhhWf5l93haSc
z2p2Ol9IcbKHizsd9t3xFXdv6ttPmFFjRhCit6DvAFxcagcRWoyBuZ0uK6WnpMG089r2XcB/dm+e
MApjyp62r2QdZ1EPqFE7iTKAzmHIoiBdq3bXoL2Lo+KlRe0MkNzgzfvFmjDJWM/KcAfVbopHj/br
fyUt6n5rbHJlxIPF9iQDdeXJceFZo2GFKz7G442PmwxR10mL5UUOn5oNrd9VpJT7vcoTGK9ZQmB1
wYceBk7AiyVVvhBpxylEyR0PyJ54BW28RbL9KmvxB51uPOqo4Coj4owQc4qlL6s7V0fzJiOBeESu
pUmj7PHeseqMcXuPMD894Zj1m88vQHRp+viNRP4EPq7D667QAIwZrFxzfCCCWT+jv8cXY8/uetW3
mZUgvN2r5KeS4LM+o3xyllHjd+mUIHwQzlk5LVNTGGO9kj1m7g2yxqlWvz3Ia1HBNVcmHZ/YVch9
6vWQlc4YfXLdXZRBF/BRikRrHqYPmqEQ0NH6PF/wQd640G5bqTKriN8Ntz3nZOY2JskpcxBkVYJ2
O24GIPmO+7+N5VF8qERCCUWbq47YXK02In4xuckH1AQDDDA52eQQxBw4iXQyk9lo+0SA4j6dRUEG
FBoWYqT0DY6TcXaRIYUx3Xl9/t/4CW+N7H6W6uNNZinBS1rAU+hFRMqO1nlbzEpnWnYZivzmJEei
B+4+Bk6z5YC6nmQ8FftKICcBkqFbmUBPWwXciNXI9aCybEwt1eVODcL8XK0lNKAXOilLvDIof3IK
Cea/N2lyQbeVe2aBC542s5fAwFyq+ohhqvrDopAUbmlnJg6hNY58+ETnASQrROIqlObBqQ5pmAV+
4f24/QnCILGxbjCrdvtVnY72mIsK/cDvWrNL670wyQEQgiGbYmrc+vNMGBlrsAji64+kC/M9XOVk
42R972jYa8Gr6fd+aM4oPT+vh1ncvv9jZ1bp7BhuaN8bElLuw2gG5jRpphAtgYUoyy+MzAiV4SNv
4LKaW67DO4Lua6/ULv46+fNxl2uzyrj0HI57l8d/KfyP1B/hE51JZTuT3GbArU7aPQwH97cDloTu
I7HB3uqbYgz9q+8Xgt4gtjs0uzD177pVCk/yfp8S2gTTuiPlYAbbT3MSQduIrVeO4Ixk5eyXC514
kc/xb80+Rz4whHVn+opnwS0ysrlA5OB7FV4Zn7Nh2nBokeGqmgatQ21CWbamSqVOTZTGjd1KrMaT
1FixKmAdWiD/2gHP2zIMIjHR1eUZrCdsAsP8kg9dR38SUGHCmnAXjSTBQOQBYHhEP05PcsPjRDpo
CeBsT31dQRyYqPMCdjdQ7c0ubfTp4WSP4oP8RpjGIdCRnXrVfogBC9LkemZQ243mOMncFc7pYloL
uybPxX3t2tDe5GbgbpWhKUrdHLoz8XxJQ4w2QLkn077rS/Jg5chzuJ2ZhyMDuPtBs8yNmhiX0oeb
GFlzvpi3ejyfk7sp9uiL3OUhOFnIP0JwZksxL1EJGWNonOTXZYHpfBlK2fZna2rvYwMNW+E+vNFP
Ccn3wRuw/rjbFnuxj1K0xnHYTMKxbYsANcXmvk3wzLXrcSkH7eUsPIBez7tLlspSJDkSXEVRnCHu
aFkGT8aomB0WUOT6TtBa/h7Xe+wVnfyYvbvzG9Ywp0xK2k+Hn1GJA4m+mHclGaq/JTY9eDb0ym0a
oa+ZVUdCadAmgHCJk77fP2O5NWaFMXrrOH1M7Ez3X+EcmEdP+wvM9vPOFwXE77aK+qekCofWMVZ/
vfqrmgYauLy8VzNtYe6FPrYfyem2u5v8cnirdERc4jaYhWDUKaVDu1P792xO/xBFO5+tWe0IFN1m
3nR8e4Dg33whbeNuxpk8XEL+hpx39cE4gg6nqSW62TXbl9TFbh1y5wTAljVVXgqFP8CkedA9OBDz
PG4v3ZSKeIfqagvBeBRLBnZD4yaMyhN8xfik+zr6mlUMEcgvUITslXb5N7tmTCvdVsDY0RmMvLdy
fWe27z0kDEm/0xNh/eAS1eN65oQmCBVjODxp993ZzdD+opv8TsPVMYfELHfWwXzAn78v63y2S1+t
IoOIkja1afJOO1Ai6zpIr7pv5x87DPTAkj/pvG4seILUgdqzRkbC+i0oubuOnEs/kNWMu5VrOFB2
tOKTFjCLY7LjSlam9vVjyyeaXhjzxTWlDcHrJOQ99/UOuwEhN5AJdq8vSKsyGy2D0dJluA2uDrbG
uf85i+nGD7i1vndp61lquxOqObYoakzc9GUkOtlGx6RfVDW8jAuvjEUaucoUbbJ0fD+D+ID1ZeT2
0BwKZz0lp9xME0pQPOd+D8p+Emm+lylXXH3oWIAFEDi3OeEcFWqEdEbV7DosZQlQTHiT1LFzxyv9
A6qqHlgWRnOs/BfuiBZKiQ2vqK9GccMRlykrPtjqkgWnUVwhdOHxwUhCMZhan306ReWyHTJQVg3W
m46gnIHAxj9tnELoD4dZnuqHioRF0tcPWEQHTQRds7U9x1+bLPKaXf9Pd3G80TZoXTLY8gWr4CsN
MnOOEg4tpeS15TwLNH82IOI15w3gqEV1pmQ61SRfYsUvTcUPp7HITQa9h22MIeCC+7LEitWT71i5
2jiteupaGUdcjoouN4s1J9JF8kUQv7fg40PiD35/NjhN6FvWNX7iLui+y0gbQckmKmmrVEENgXmN
H3vFXpfnDTaQW+qZjmC441SQmWRqKmOAjrWgfou2C6NOAu8P+UnSfklJAWjgS3MGS4i6Poy3XJ3t
hmOrY+Yk9GAzp2HmoN86OGQC4pr0oVty8n1/uK44Hemq/LE+hBiLaTti0c+9As44PFk01zc78Ftm
xXJHXINtRB0iKU1VtbH+dH/ypZ02/e5HdFS+UZZsjfeWWryDFSnSy+E0RpcgwmtLMqBsEDhuMtK3
D85doFnS2JTXqDhFkiQChaPiLrkkuj3rzRBmDsTy/Z3LrthueQD4kbZb7bRU5yggzYS5S+XAgMKL
JSo+UjR84IabtTA/DU3MiYAwiifHX4pwtjm/uOVtv2CEFWGuSMF00OOVmyU8WPLej5y01bA5UpdY
rAjbN8ynwSXOlhNHuaeTiGIwNbVN2zTH4MAc4tXiBWAcnK3mJK9VwSH8I+2NG6qGmicANJS10jRv
29bQMY41EfvLgiFGh6g8Edu1W3ej4EHMBScYXsoxWeuDQGKo4hBo5a6af4svEXLEkVXH7ptdq0Q0
p5aMgTBG3TXEMCbhpkIVDS759R0mjVh73NZFrdAsaTGFRIpQlgOXoTennJenNVvfBEh6Z/gFlAAa
N7qgSLNJwycuePJf84iPNhiWPK5p9NeNEwOy4IkcrTlJHNFS+83lMrkBqwzUZRPHUhScSHDZFAHk
qMma6BGuF7RWGdUTvJTCgCgGaDOleu5WMwEYgAxikkhG/qaoFnv+dGmQSTzySzJWNGl3wJ3NROBt
LuPQNUL1jTY2YGEgQTotMklm/YHfTdb7HExI8guasS7m8u0vtIVVV7Gjb57uB051WsTMtagN+RwB
/jQxKvJ4uo+7/EQg0qAVZVS6RWOAxeYJoQBC00zcnkkTy238xQ4vL6AJ9lOy2Vd9EeW/vOoNOtMD
0Ar/Yu+XG3TLxL6eIBmeSY9k+/vfJcjjBqwWgGw/j0vpu0UpPPKeC/5UY7DVR6owAOtrv49A5RuM
sDchvLqDbVLVy80VbXGq/XR0KViwyQmOestcj1/f7kWRQCEizildzz0Y/mZi8PCXpDUCm3BsJT9T
1omX+auR1c3Wze6FLQ5RJkmJUIxOmpk4QfgBF9/CYWs4Jj3dvxJG9ayfa4WZE5IuPkItdm3SVBE0
FvzLxV9hEkuSMMDq1wzSTT5Mo5gN86urVfTYFTCl0ie9/xXYVWrzKt00pKR1M3/VxCvfbh0XMubf
zwVtV6TrCl/0vikpL8pDGGyzbvE3UBxU+I31ewUdVV8+yr8MwaK/HxjHESFCdtLN8rruPBSWwb3g
kr4dPoXuKXWayR/52ZEp9OitDmPe/iZnLYzKUa8RgXvGEq3qqLSgVT4HhINbNygy1v55KatJk5J5
oYpYBAd47xaJHsW1ZN0vj9VUO3D+ORquots9IqtnWsACwskx7a4z5KC+dQFlOg/JacCS5PJBdYfo
8FweGEoSzQi3vgLs6mgRHVBdUCpbaVE5NJlKZRYOlozlx2asoyFFGhhqJ1BWrpfW7vHJhaFe1o1m
yXlH38h/uMKRcJWCbb+k5pIwakSeeUlGedKjGiNIxV7vc7t+CQcxCqSdmY6rQzDwZh0HGSCwW9gf
FPv0PKRLEFnHkbj1JvuHjV0rC6Rojfy7lSfyfcG6BZXpAtzH53skAA+ASRuclXog9s/fY/o9wnSV
G6zlu0e4vhJjE99Uv2H+d4aDR6xYtJ9MZCqJ9VG4YD41zPr4HS6uyTJM4FrNMLkhmCvAVSOp6RfP
PbprqhuppQ0yOWQGYpDGemCf9i9JqVu5b99BcbXxCDrmR8B/WrhrfsT/u5OicQPtKOtXJjEgezl+
eKU32ughGTVkpaG9AOehlFanVkShCpLTToZ4LkGfaQgNOO9jWyNgk2HiSsYMw5rdb+s6LUWP7FV9
jBK9Q3VguwFwQXBayFgzIfN2chsvxYR3R5sTJv8ykR9a4hzq1uim1+FuG6JYFJ3jiaM+VMSKwhnH
Q2XSpvDNpTMI8TpIXnHOt+TwHzb1V3OZABS+66fxNY8RxaIarcx0uTgiSEc9E74iKySF2R0FRPYG
5ljTmf8DJS79RCbRBqHa26ZrKkK+zcmhys5SJ2xEsBJSs02Fbs5IAb59UiqtS7CCMljEJg7kFncb
vnyRJSgYHUP/Ehh13GUr/vRsXfPFHi3viZSrYfCl9G3KkgUXnvQ4mpeTLAVj/jP+7Tl9KFZANJQ9
kCblxZqADXC8ddb2jvLU+tlqQk72fps9lxURsZuZkEef/jZAyZMiG0PgJSkF5LJYEFJt+NnN1Pgd
80FiB3jv46ffFZEVQfHB/RZSSa30aOoEuPtR9e8u53WIr4R2IqAPyicNSYhW1tkii0mXBnUZh4HX
3iBlNluraS/DzVRC4/Smz0CPlPDUAUdnJtFxNPVZUbSIJoaCHY1pJWnDTFwtsSZ+VKa5MJJaBpza
XEnCAyJzAcJj76oNGHYxIi3xFejH77p5OOj/424JVCPmifYK5E2IQI7FeMvCtdLFiAo322w3Ipjl
XaBDPAWMHGtev4PTq7D1/MWTup/QOJxXH7Ze603CA3SkwXHj4DpaJuecSv6iL/ncsttRTjqw/k00
L2gl0LHvs8rKUP0dd4COlK0daWAEU6zUVwL/B/Rlp2qvwKrgel7MSn23YdLH2HbeHJVRJwjSkQ4D
aagVSOLHQwBhOmlnrCY9mqvWgsi53cBlRpQqxdSDvO+xDse3igF0bDQ+OnNF9swHH2waiTcbUQS3
HVjApaPyLqiIhR3JEmLiQLPTiW364mlzFcDCM+mmhwiK19PTWJkXDbnH+rMVbEInegCOy/iXxdme
rZehSSepxILVMFI8cH4gRhkwMxeqCQanXXoYIaIb5PETbEUZRzpZd7JgyPcGrKAWGGIEAbIyeIam
r08QSTuDdiizZr1hjjnkgcEF+WGUKYuVIt8CKkKIYGQnZkHDXswIaNDr7OaHcIpF6NcDXtqMqyj2
X/JVcTyfkycCOU/ZSezvm4DMNQ7g5Tz/+x14FbTSlZ7XHXEzrfFa1Wl3H/ldZVRnVIK8vEAvkZm2
AEN29QG2GN+SvFUmCnTNIJBN0LrVSZxqEW0jiAnr3dpNPJEo0cmB8Vta8aIvUxX/TIOwDtSKhBBH
hvqvp9hOT1ZMW9VgKalkRPlZ1nyjG5atDiZwUFGuyrc0ruj3l+INJtzd1xVuYhFGnvfJsqa70NZG
rEsystIldqCRu5c1Rk+Ohd0w61P6fVJU/4n+JDFRD//V6/Z0GpTovSq3ru3mDO9L1vAlOx9gtZS/
I57QO5TZn5ZyYkhgRHB7oFzzuy6Qwqq9iHsOZrGHWYg8TkeoxkGSKf5+WFC0U6xR9POfo3a5zZbZ
8+jWhbojk8q+LoPiqwH4r6+2rBq7gygjTG4KMzO5iX8Ic+9k+uChkJIFLfbeUrJQZpsrAh7p8ssx
k0F6Ms1Q/bpuVRVQsHyniECbWD/EGVnXjp6/ZYP7vr/06WBa2yNqjt7AT7r2fynXQPub5YHeX9v+
xerdbbiUusvqjUQFn82MYnHM4CrtUT1CNnlHaA1E81sBnxkpzNTLBlb7CmUKS4TvrBq///bVqwQt
6TqcKEl30ZSboBi8SqqgHRwGZ1AnM6STLufHTmTrdRzDtMgvX/Zt944XUeansTQHcu6GAxr2st5N
8LxVWrsa83+bhh8DcsDOscBrqRHibfLe8F960Kd4d5KWqx1u5Hs8VRhCe4MWhE6PgA27lGTudZbf
CR6bTLkirU8TD7bMi+wLgc22pwMgTAvxTOHYpwbi7vpM7c/nn+YueV7nAIBB+BKj065soW51UuWN
QftlLMx1Q02NsM6CWoJFYRJwpOBZaqymNTsEM6Xd7CqtKzuCK5oJ7XN8sFINbJGyqmT3ul3wajVc
EhFB1wUr1p1/bztG1nv/ncm8T5jxCVGySAmU2A+ZZ/xxEfJrUayxs4QQ3V5jwk88CHacJmPyUnQL
60q8ZCy77gPz494gDUUNl2mYTrYxxPBt43uCT1ta193vGwigSCagr1OjJKDy6zAghwaOJojd10g8
4XnM4BytzwMa7lpqx5s2AkMq1dcw6EnuuvCStKhqVO6ufV30Hm/gyIuVG1JMDrfA1HvxL2CeGE/e
6nnj79uhDi0yQ3gZMlezZpF1yGC0vxkk7dAU2lon6p5NcZHsXGmOkWLEbvi5hugsRQElc1PVpkor
u3m4sWuJuI9h2GcgJG/jlqg4hzyGxRYxkZXhtHB+WpFlNkr4w1v2fOSy77T+6HKlFrU5teDZsKwb
1QHp1DYtBOfnXuyxJ39Qlunk5GPDp0UX2yWTAvEADNLF9S5yRpUfJ/4ZYw+OwS4mLYtl+jkq4Hj3
SyBnMXTv9mLaODEDoXZP2A5iclxwGWmBqlIfwaOVqXJAd4E818MmgmFBhHn0Xx3XZ2+nz+tS4cLC
yZLa3YOVo57LFhyA423AbjwSQvwVdyej14ULksZTOk/i39NCssGpqgcG4XPMoQVRLKo3bpjs7ozi
rXCFvvYfW6IZtkVyWYUlQyazgcjGUunGihDutVj67QpvRYLpz0U2DGtqqau2mBj4V6gzrGTWCt7j
PGEu7pP+NxGPm4B3kaEvrgjqKh1Lfk6OSW+VkUXK6IzH6RDSXEdvDxN3QcCvd9rGkCHIN9r5d+a5
T6Y29y5dBL1CI780LVNvN/Lp7gF7YAOGlCdo5QM+pl3RUFfgX40jcrxeZTg/NV6dudlQcNEODjch
yooUYGwJ4qIPchxCWKBV4np8RMibj2wrwVdszTZTHkX8WdQMYl4B2gvGmsqNM7N4mzZgnH+2XGs3
F6j3HOdYBh0PLEzlqLTZL9lFYtXw1Ufv6sYHllvSo1pnSDYWSaju4mUMG+b/lbmwELW8WleWtfZB
Y4svJmzjOHEQvy34SqwaGYxkCl0qWgF05y8rUnJyAJeuY5uKdYTg+3weVdZZZVeAi6jcvmlBpAbH
8yfhAE343NqJyLsep68+doUMSGpfRcUjWcdtQ4AvHdcFtEHbepplxkGE0XdHb7/PtZJMESgHxWOe
SV8HATqmLOlWCjOu8ZRnBtM3aGiyTzVTtbFdhnbPDn3/IDQYDxAzWU07vZC1QhP19BI+XG5IJbKY
IGhHeh9IpjayVvj54jeAPxE9L3W/7JMeymXScILOHOkXSsZNAtRdn4YXGqd+iPsAJ32R4X0PgRyJ
Q3ZxpdLKNqmlJQM/tB19ZhsZHLIqkDFu6iU73arA8SSMbfIcO700+fpXbLNODItiBFMqYCV403Wn
xOHQRD0EH3+9XrWwTXobc2lG0offVIIsHSUPQTAHZ4ZZqmmt/WBC8jEZYHzmAcOTMFsUUH2ZOZQm
QL56MczilP8Sp0dFIt0U0T7HYQuzAi8l7pck8FsPw6u+IG6aLowkiHku1P9tR/OsNj79+DH/c8o6
n4ZEyyMYyHn9tx6gCL0vpWMCAzM5c3lCbIaScTMw7+ViBMeZ16KgJWCe/Mn4qPj+G/V7ZEBc00+3
BBVKRDfsKslrAhk0NJTf0QeaduLDkVUdpMDoNMbJ9c8Y9lPZyTY8WsydbEwLLVlCmjtVvuau4Sok
eLoicNPz8Lpvl+HQ2JhIhfkMYbXkpX7XsYI3rWmElO1oXtp7/Sxli7/VLCsAjezMj0FpiVDhcNpG
kq8kmXzwtK7U4VLGRxNNAP8vXREUYR/+OH1HHS1KwTT83cT00JrsGM/WBjLiG1ZT66jo82OkEzMX
h8tC24JEdbiuHIwvWWb13m1YQVSGQIa7oq2Ht4yeWbbhvucMiBaug1V7XqUNeGVvHyHsqnUqktlg
/Pu+Zrsq9YqLbWV0gtemaY5oeFoKm+1S9c0Jh/H9k2tAnPFlnKP5/XdZ8/5pe5y8moynnYgyDNg5
t/PDs9aoKM54wGHDpEtUj14mAV+s7e1phlIMy1kR9YqGAYTtQfiDYygk+4iax9PIQUFvVJi87oot
5Oe9STs4xumiyg2dp/1y5fHOWvcbzWq+JoCK6ztKJIH8MJImQGRDTPDR7jIT0hTNwti4J5tPfyIH
6eYGh4Ga9j5rYFTGzuNrng8Vsdrldzmpstxz2ZbUibaz4s3bq0m/xY6wc4wEQ1niHYw2YD+DMlzb
5cS1A54nxBKfrl3ZrRLG3+kg3CLm910AlGNxGc238czxigZi9PRKjIc2nInt1UBdrmqovg0vxwHh
tXa/qW0r17lTuF/FGDlRHjAdg8oWiXcYLdL6YpHv51JBx9jO6K+5jW+s16wElB0Cw20UMwZ6y1dW
yvlHcm7gDlAknh2ZuLBPb4NhaNmRVMZwgJDg7o40g5tGAWRRwjwWLrHMKuTkTwt2cF01TC0T0sH8
BGF1uTmS1dblNMQh8+tr56GL5uDcQUODUGO+GeaqqT2RZAwoDzfO2zP2TOh1rHDNoNKF5SzNRow4
F4BiM+NR2x4+mB0qnkq9KTzbBxtgrJqh4KFmK4rXebzsDPKrJlEwtudnK2k4xoeuEmXrZ1xFjUqJ
Tm81fTOhHzbcgBY03YFYaNweYeyf5YrPOrynVWYSnwDdMRPCN3R1SfVfaOWpGnuzBXvHdYnfCNgv
sqhIZzWbWavlolbTwsagv19//Xyp+iEYa6JA4ToimI6n79cadaCoNKvVKDU/BJiXQ8CKEHME5bIb
+H8P0luFPiWzCBp8LvFum4lkcokHPRaEdh2IuN48+ers715B4cqhxA4Kefn1aa1RA7EtOapvx9V+
Ym/auubz3fjsWRnAL2txwK6nXQrVqB/P2mF20/067A2M6Eu8XviQqbf0M6YFaM+JiJxfJVQOK+Bm
XcmSWPBQtfbN682qRIaXH8H9eA0LaqZHRbMDQAhz1P4roBQ1UULDLmo4E+LKz/NZhVDiR63xW+Jn
CxQpV/eAn7t52TTX3YE3swglZ/AV/tL9ks5yRx4060SrXd1nBdrvtotQxDzFIrD021LQwTBEL3GN
VDZNQn9ErevuB7W7OKHbZbq5+R7CuwDNaTyr/ICsWU4lHBCmoiyy07vL5iFfy6po6PasNWDoluk5
XKLKY273uc/SC1csOasPddf1Zzcl3QB1gTOVBIrUCGcgSVTLX7GG5qeY5FdrPUzR0XtO3ctN6ZFm
tRfn5XvxGwXC6jkDXyRKIv1mBvONGQH7hRtHpDWPDr8dXWwPZcxErMeEAeMpXiwtjDIeMmJrJkq6
F7DRZQjPWXQaw0j6B7oU3VDIYstXG6OhqEirGVGSkqk1Xito/CUBnRD8+eM5M5Sf8BprGEl4gwV5
fB5k0uKkPuVfRGQCO9iGAdglBOBjxLiKF3LfuDK1gltjOzSNPnrdbBGbJy0tiLuEkugi5MgRUBZS
K216cfy4XoH06AetPgdW66Didtx2WekoGoOM0bNACAO7I6MuLElna+fkExNSF4hLktGyhOBS3U9V
B78Qpe9uIons/Kp8Z6zplM0N/nbzKqJ5gEkrdibVshCGfxG6ajtbxqQAp4TRWrtSSzwLHkdbNyZO
d507f/Q9S0ZJ6Fg0l6dIu+kBjdn8JHMcAXYelkQrdr3bW4N2RcsZTI6fDpSC6iuYDfgE2skslzFK
xbxZICoe02IWYVQ8SusMl88bPImGRVvluEnVv4laplHy8xz3rU08ze11aQBr1uyiCrvnmJYkhaLL
/k4ZZBs4MaTHxunZyYqT3bf4K52bKAo8vNbhzM++47g81Ki1rdKmNRdc9SfMcLtvjh0duL9Ef4qR
iUJv23OV4UvjofwIEy3kNXX2mkl1qe+k8baoclinUJD1ieHuta6loPtAjWSBNdP4vxwops1MnM32
Fy7TPMM57qblmzc4YZnoCtEt4YMFFm9dZm3xNMgjdymPqWLrjnHjxlnSMHeOs0QZ5MOOZSrcilvb
Pe8fVeuKuWwk20OoXA8jPCHJRYp82NwjMP8PHjoBSUPTl10rV25TqcJ/qAFjeFErY1rEgJr5Zoh8
bhAtCteYGcrZCm5U60M1qVcPjfx783HfoAZ40HHBRYI/qmqPcSlnHYMIvUD/j0DE3KgrlQvuKpGW
79S6kxrWKa/qsbGhBzMjeMXGBprspk1xdzJOr9/kBsU07wvGwo1QAOVQY/zrtZxqITiIOwPlDXZW
n8rAW1DwbJps+db3vaFwmGqCJ34QWI4uJuqpVny7vpPB1j0oTm8G77fJ7wTrMUzplBBlVZZPDgpi
felDG4tl3hIr1fFY3PVLICD82h3EOSugGZTWKDs09u7cNAcu6pPTweQrpjTzXhLqMySuoI3f+8aV
9Cjulktvw5zwhHyvt7NtMuM5TLzZ+lma+mqWvM3uoxRsv6Hm8OPq5Q6V3AcD6at420OEaZ5cgihJ
zcZ8LK51llwneDY0jC/WPBcRvNYdmPcnO7U9mrDvB14jYAGrGezCSydUvzHvtjX7Ieql8RWGkrL1
L1Z2cTLDTttLwGs0MvuN9kasEb5xkW9E7sXgZDpPaAcngh220yNkY33ae2iUD0Lge0zmRQjXn4VN
QlgBgbGb2BQnF4TkovOSvxXjVVFA0LdYkTc8whsryWj6c8qP1kbGarVC2m7lw2L++McLSIvsaVQz
BlZdWlf/hYREYk0l2l8qDRt6QZ1Ah8kgbjErmQFqp6+Iwp0hkfNqKKiAZQkvTvHqfxu3KTAyiBE9
TiDMy362No/yzkL0vfwwkpIc3Okwwh3zPVOQJT1yOOBOFuZsIHWBjLYSAV2j6MK+hEDySHcN7vEu
g1VAKD/s4FJ+dZGVDmufNnu90ByLrbB/BjXv1zJgGZLkPrGTSXw2kmxXft4uosptRHrogA4tJJ6F
1KbrP/wy9baJFz+bktG1nup/3TDKyXbGCHtclpRtbu0myFOW7F9VTvXU+E/XNt0Rl78ZMLmJ7Dmh
3zzAIlm59yYYmOoeMNybcFdmtQG59plDtqRcNln5hYAg7IydC6pLCRFF9sBvW6/W6K+16nPNjiLD
wT0tzAPEWbts30wqomKz5Vf6KxHGpoy3uqtOOOLybIpGWrHBrDIDR7/rk8uhVyfQp1Fnp2p0Z+1z
bpSKb6O7son2qxR+em+icp5ej2Nl221umAmYVW0cqTfsikurKmAYc3rJFOoDqpwL1Td76Xi9vA8o
K6d6JymBdWf4VYZRALNgkIYi0btM0DWB96bGGQgKDf72d9jLL+Q05H8kQikL8U0fhidU23mw+mHF
l41UwO+k68MPrVeZpU9zSpgYiCgCFK+On6/QDiR+y9bcnf1tAM6XSJU5OLgnQyQmDy6BwQ9c+qf+
xILI2wxYYEBiORWYrsonMeH7TSzj4w+4XUYHO4D8oy1opwzLtdwZJvEzQXGECEG5HrLb+6IH6hG+
CQfXHyHXa1+fuIh+QK+Ev1Qgeb6o04SgRL8miw/RQO2rmyz5+Nj8M+ehsGBST02+a523Jek6bQEW
K0qmB2TrMnyIFiuvPO9QOvJpQnGIgORx7GKDxXY6vX3r+D8tkWcHZpTJJ0Fbqv2C6fW7lc+y96ci
7i6fhE1f1VWjWX07g2rkq4ELHeKDVBLXHECekNq2OoEttU54K5d8rloQ2AKucCBhsNGDj+HegToS
OMrxnVBCz1TY4mglT7LdJlz5PUcC/6rG069BI6uctkkjYTIrVpRrd+FoAyzmduEUcF00GpltecMG
LYaxZvP/OadnSFNILpLlS5qkoqvLQVGJJi/BJYC4CU+T/UifoJbZckJK1ng4xDVEkW3jX4IrXNeO
LxB681RExBz6n5qs/rSzgk9Mc4POkWmhJRPIefM1H3hEayKwzAPD19tTyd+j/sWpIKrVPk+YABzs
knBuORs8wdu1n/vCGsZMobtcLQB+auSM+tXGsnxOdc1VWA+5RAuZdpiXSpTz3AmQ5oklf1gDJRM2
CuuXh8MzQM/TbN2Ok3ptbNGxKCUF7QOdBsRiPh7MFp2hHhQY7Eg/gaMrButnajPxd1hHCxNbHJz+
k4UHE6Yq4bi2QyZlX+2o4HirlkdVabG65y3BExJkkHuLYmeQRm91TCwE4+n1SH/I2QvTHuNfwho0
8HLmRmz6JOGBe101mi0uWnWI6N2dO6gFXpyjZxNZVRHmj1D8hTvQ79GVkqSSwrfOB45bBZdnAd5d
tJYB/20iD1OBfDYjQ4fEBJfWU0Hdk2w1f6K/vUzw7YLznsgutTip35k9BOOvVlbZNjqzs3NnfCf3
GMSMf0YtePkJn+dvx+vl2u33LYmkj8BI8GvDvT0anFSnTav5kOyCQYmIUc/+yJRupwz9i4vT1F4a
ZP8Hhm0Z31rsL6kqlQzjDfRgvxIsdWZfHxmw6eWS1Jeron7Utw9C9OBZNEBr3yRji38c0wyM/u+Q
TVRPeNdf+KQr3saNtugYHiLn2NeLEnoPodUMbxIsBM3K5SLFQqYvv7mpx9YHlJ0wQdI06p0rccGd
c56zbpwX+udQQ0GOUIMvmF2L94Oucoq1e88KHBJB5RJ48shKaEFZuFMPlGqYr+hOuSe4dy+49gXK
siYsgba6ib6lDInKKvp8fRcne3aoVaWJMdRj9PXVaz0wC9/ga/0zK6ylHW+lK9u2B/6sAU+iZ5yj
b0J8qqntfAErEJXPDVSlSQDbCgQeuUHMes559R3ouZLRrQpqPqGxXfmPL9SBVjmPUu8vY5mkB91i
GQ1GbCmYMBagaqZKQpCDQatmZ/xDhs2wLUz8kNfQqvkbPxdiw4CbTPzV0vXu3fUNZumKzKFjywuK
2mpBBU4RNIE1MweZi3clHvP7Jn4G20JdT207R76Cvs9eeuiwhLK9o2Xz2ddcAoFmQY2Ee/zxsGvn
t8svYK2yx69CQMitldpCeWgHhpyO/Kw12bxGs8elkFVbWRY3col4khcy3PJ2zxnbdRxyRL3mBpgi
pgZSZKpPi1RH04lVJ+aHzaATZp4jhhrYbPQdki0UzpD+YYSTN8devIWVjq13c/NU6/actblM+kfx
0HHj7/GYI3vB0aRMns5DOuY/m82Q+aex6/sWqspZwxAQRJ59Ft6jMNNQ4G0XMwSwY27BUk+LEoxH
RTCfMvQ3N8i91F9W9MrSc9wv+/Vnqy+Yg30Co8QhEOjAeC+k7QKXNxJEScM3VcTVgBFsV2yedHOz
qqTDU+cX/PGIfaTsU38IOGF4D2tln1/6PxugyIpvvVlgcfi6/+zTyLroHHicN2gpqT8atdYhFzIP
cAfWUMVorvtoT7FBki0trkP8MkWab0u8mdx93fvccQJkRY7OewG8OvvSKaLvw6kBwzXangnzz/0n
sYShoqxPYDwB+Dg7FTgQInvD3yg3s5zmSf2V0p2kUFRjXwu1uNxMaMRJycwnvY+nOQIP5c1HOgwy
sjYlKRAWjTcVbCcbFV3/7F/fATkaqKYe/dVxcrt2NZo9nrTtQkl/vVhJZS/twfw98vMQWOz1D8Qu
wqD0ZW/Z/BAXRXEMhBe1RHe2M4zB1QIwIO9fH2s7Ly395z7SPSQXH+cE865Ul1scUTyo+tkceu8n
I4vph5J/EO2lP6Ej0lM7N6XUM6RiEI5ansfggOhaQTw4CHAXZVfVRk/J9iy4IhDSE/RtbAlbVSqV
JHYBB5sRnQclj5b4mtUHt6y6QRXGViH9tCvWwW6WOqx2nSiCnj8Vt5tpcnZDwI4C/dCuc60uS5tz
5dnIxN+ts0LMJ4mOsvkyzmSB2IZannzVqscGCsPycpJu71QchuRr0NaayxuTDiTxPwcd626cSOew
J6ZAq9w9XkTot7uyJVgek99TDHl3d683EXBEgyEbh0GI059/hwQPoe7GMU4M7Qg2nWMp/IIc9ulw
sbuTouVpFnD2xFuWzdE9ViN+x9v0wf3DdaTqpTABZcaxTrwL2Bq5uMxic7SeOEW6xcjtC1VAl4It
hUtDlmjTlRPoS8NnAFw3CvsKNgiG6Na1qU/5r4s2KJ3Dop3WqMcKJCAu59j6gFYU7wNF6tmJ+lsL
PoaOw9RYmWfz4I5ik0GCOCorECRXYy0IuRqYlquJMUYf+b6MFQSJMP9ZzQ0mIt1sjk3AXADtCyq7
F/kxBoLkDfk8o4BKjTDpAFNTx+HONzWF3E7jrYuAsfZ8jYY21GGj2wgpVaYjEYv1K3syMfbxHv+d
R/gYKwhjrYpYn1eAbw8SUhFOZbYPuiV/ZnFAwWvX2RbREVxSnCkXuBmVz29jdbK7yCcF/Imq7Mt9
g8sYua09ARAMLBBvbD787jrkTyEd30KwhIvc4H803Mk9zKmjtmmWjV8dnjL3SOQGahl+o5ZbaTXj
6NpmgSsKQ/kWE5NWS6JpbLlT1L3NhhZ0DoMMbtJXuJrH7CqPi/Oy7fmRf8anqLqW15772Pw4gYSH
6dL1UQZfcwS+lCrvJp+C6c6p2Om9eTT2sHVmPen8nEXNGwzYSDYCmReZnB++wIFm8A2EFdwUh09u
YwzjQ+Lp+vN69qjneKO3sGo/PPHahXlXsKLWBzhDfqLAoFjaB7hsUJhzhfgouwbSswye5vm6BaRQ
KrPo9IrY3qyfJmwN/uKd/w75HGIUMO/+kz36VCueECS8jN/dsl1EASMhWlW/gNg+Ym0UwE8X/0Av
NS2Hjr3dqGtJrrVKiJzznKpLT24KAplV/CbyPhcOqpvj1ZCOsyiygIfonxVC4vLwiTk8p/ihI4Se
yXPpy4+42ue4aVcgmC1p9PeDgy3iXIebSlGvtx2qK0sDDOVwibRWvHcXUZs5jRVyGZfAcUrH0pRR
d7W+VrzAg0MHAIdm/tosMVJYm6XGS8gix8MzOte29MQ/GcGTZzbrK5UiKL2VK5HOQwm+8XdKAPX9
wRlhaOELCM3q8lP6LdT/qwz/zJ3VFPtneQquugCzSJLxuGys13AL17h6OdhGKtqUXqKKh/6nWTlt
WPct+UbvBTyAbvLA2GHLFiUPabedqZWPZ/R7vaFDjP3hU2ttRAcB3zL/0dvbN6Nb+KT+t7AXyGBB
A/Aw5agcjugVohEv37KNREFSkqzk6y5HGJpOotNmND6lOjguBbL4PW02iyMIc/TYB+kn+4Ih69Y0
P0q0nkcsuZ8P7bfiINXSRa+N00fLtyx+MG3iccQ92Qdx9qik7FRWNmomng1J9etO3sdKtNROS4nV
VEMsMKU9cWGWJ/XMZHCX9XgWn6CwZDFwb9cUd1XGb/XzAj821WqPqCvCo8BhkfF1hGLwT4DZxMrd
F/da2sMLJgekUyalW6iukPG8uR7tM51CLhntRs5Cj/OALbxZnC4He6APdtwYqySkMnKlsy3lI661
mbQc7QQ+b7ugOezLDs+lRB8DhbGwKFnEU5qg7wMySfkIPJ13Yta8/CZSBCHqjN55eWsRN1m8q2es
Bx7Cr5ST0MDvHDtcT4jYR0x/cW9Syd/OD8aGUanE80S1sWxL81XQBcX3LV6ySCq6PHb3JSv8TfeU
3w9xtA+/3lI9E/IoREhzogf2+Xzi9UqYmNLzRHnGYoboxtJQfaKwPprIPLgrA4hpdd+cYhfgIjO/
nCSMs9gx/ug9IO8v7YHRFySpi3YTkLLzx+URT3aryILLKestsOcvEGa0hXSvm8T5f7NWRKwwSqi5
9/4cbEMSVXNjOIKmhSBWPyu70KI3ju5epZ3vDR6vP/0IA0vq3+DMrwxQr/onkGYQaQKQrNSES2CE
Czt4LxUqT1bpD2MZPTbImGPURNlMiy+IAuhO0ROcJ2yzzg69Qy7NJy9VoW1VFs0rnECrFtOyhSN3
yL81yzaM1FB86A13e7kdWGmxAExkdWe7mwTCUqKW2frp83E4yeWtpcB+h7Yx1/YNj20MKDmrstJz
rpYUzRvETs7VdQdKak7/0jJToiO9k8NdswyWtAvqg01/2ZjWVp2l8khhaBqoN55HqkRzic434vtl
1r88J34m0C7FWzB4UDt1HUb2ndZwOzktWlQg3VVhCqe6F1ji/YqKrDdYSocHngtuIsPXqfIhQhk3
ka3u+Oqz77jEtdDuDW4jYFhy5TuSaA1Tx8D9VuwcwdjD9R07Dv8h6cQosKRyqbBCOxxjaC5QUBkH
euy8Lhl/gA7hF/SjY1X+Bq/omtb4v5huP8R+EOwn14tQ6s2QHMviZ6C4+0lxM3RGHHFHXuRlF5C5
VoxFhsccXnWdTBHQiSeq6eO7drkOXmLmH4GQ+wI0/iyrBbLvtOWOhFd+acpKUw1hJfsIMWFrvXhh
PlhcDKqxBB9g6238ClbFs68MaqR0sp3W3WUULs7m2KUSYkR7TrVy6FSyEfviq0Y3GenKM5I9clOr
8AQntGk83ZtaWroQlhesWjzHB3Osgiuo3haNUQdQundzvFByn+TKqqbfqGPa7JWWh6UFPncDFdZ3
7hTuYIAvVJhrjIXHT5i+G/Ebt1PxlaDnyKiuvZAPEKfHxgZNgr4f6sTgEuy1Xh+y3meB2Z4wmhzA
mZHK3pv9FRrpEMCUOLnM3norJkO4jNOIAP1QWiDpTfSRcaluezXQcl34p4ojPN3QDiresAEL1u0L
+esHmjideW2gG6oZwI5xw2ReMpImmmN3E362PocrGNYiJ6Ue8fglHn/y1lYFA5qAARYf2i3IAZHr
sV3cfelKkbr8HErSweb7YYq1u1bkuWIfu/T0jKBzmArK6ZTIOuHQz2CFSq4xzYrZWyrNgL1CfSJ8
labQleolFQLk5fb4qqXtLw6KonrlXHHt+X2TfW7O3kBNY4yvs34YnJZnmrJ2vwcEaTVTPeqbxwR0
gBl6jnzJalmtDsv+JKNt8+S2h2+prgSTPKzOmUB442aa8Rvw+sj5tQeZUQcAClmEltbHoQXQ61We
tJ9LqcPVgCT/VoPPW2UBPQrBdzCF+lmEpcbi0/hnTNflC5NnGu7SDD5TY/ae8JAv4F1qTe4NWBYB
BM4XW0c4mJkxA02Tgq3UoqJo9NigTM9FJjelwQFYk0QFg2FQHsPpbsXrn1GfvmqsCsBYYEWWMJgG
g1nhTJ1djPU29c6RiuQngqwBUK+ZTFA6FW+/+WQbf1tTi2U673EqFDsbQ4N2iqyJveqSr3rnBaiW
GtcC/+28/B4/PZVCje3FdFFswIeBl5TXkA1EJ0uXV59EQKX8pqTz8788AisPjaEy97UmW4lf8Vl1
x5qLkpMnzqAp+C3ABrPfFiTIMYvGl/DiN2KyrPK75E1AayRe5Awd6gUzco+4+X9jIJUE6IEcyGYZ
BP6nKVD298oz9bhFdwQnFzcRPu8nbU9W9drUwksXLF1eeDUWfRuQ6zioVOzATWlASkD/D7VDL9gD
EMV5EZlmwnMELKUNwJEpXeqQYNvo6wolhczaIFB523rWx3OD8gxGMo7/2P/Mg2zuY2HAflejjX8e
ghobW5Xfq/Z7Zyyt/2dxOZ4vL162tpIvHdbb/GPGXFMpqr4gqSJ+xvV7vWMD/1YiQKus91H6QLRK
i5SbSHwgyXVJ+dKPgA3S24d6MKBcKy8TdhHAbEHWPj7+iIoXl+fztwfqw8f+HS9rj8m18MPT7HkH
fZk+TMv3u9KC/TtfKAEH64//plYvTKyqj7dlqG7QWrdJF7cHoMgsuT8fZHXDXTKPAHjmCazNouH+
OYomwVvoyHntbRz4R9aNPI8iEsu9TCbM/u4Q2dZxSqc5bhPR4A3R1esuzUYtVoU/qvdJ+sVriypk
dZVSuezk/yG7wNu6dlZazt9EvrDJujeJfoAvvvjIU5yTeuTsO20kr6ABSqzAQ9GN1qRdGwQc26Nd
16lPNXHh5oDEv5zT6NDb0SFTYPk/QnrGolDnmwKwPwDAFsZ2ny1zaS8Naq5UYbXvcaSR0SiKgLAI
IBgF7NflugGRHvlL1/z9t6Jfw2o1MGt7o6OUVkTdp5eZDiDqbkyOzyQzfgolQsMCP4iKCQ50DwMM
a3NMZM6Je7bhJkIn1IBjXg3k0WeY4NjctBqxtBigQPpvzO5tqUXPq9SFS2Y+W0xhNlAI/J4N0b7r
yeqt3gidc/cXMURhWgFsfBc0sAg9nNcqoq5JVJc251EiMUAqb8WGrH8dDrZfF3o2z6K3Fxp6LppV
JS6d7H1qXMLu5G/DkCZzKSO63GF4As/fjupU3WaWoYhDy7pHu+o7b8ZnJunYZo7OCbSO5ongyXuQ
b1TU3MgfcPRzDyJ47U/3yUuRs0BXn9TjEjUhx9qEuIvIZOPAnGDfG5f81ir05v50vTz0WcglVwCZ
AiXZ4CqxNOw/HxwzNjd05hoDgl56SDUQWbATIXJg8jQZdEaFwjs5mwvkltYYa8t6kzd3+B5bDLLu
8rGtynn2GvXDINO5wWMtya2+XI/BgaAYQ9iMxcXKFBU+DbRP73tdCO4GGYEzsJpZyPfQ6Hp6kLO3
8uGshPX+TMN6mqqAylQZCdOepbB+B6NO5Sj555Yt/ye5E9j3f+PQT24Lucp1Yg9v0aflFPUUNjGb
V5XMAHv0D4DHxOlbi2TT1G24iJ6GbvY4jtG3LVGJdFCPiJfYy5lFkUDTLz80Y4R6vbcFppljKP0K
dUlODBykj6Pj82OCvxbX+Ja0bULvrj50e2mx5VT/4XGoh5ybBd3PQ+0nfxtZ9kK2kZn6TxauD63E
zQMqT/4CfjxJHDos4YAh84umam2F+PXC+wZnFrLg9wXGutUMzUlVXRCSfNrc9ypdGqq6jhWinO38
BM3JkXyaOeW+xdpE/y2nkHZTLvj+GJo7NLnna2QrnC7/AUw1A69+0fPhabM1rNDXX9KNnlG0RLMd
dGcUoEKw4A2Xt9lpkx/VWEjmBmbJqdXGBNl28z+ptcP22LK/dzaYasi5VxWvH8f5bQMZptcainjM
vlFHCgDgEkvsjk/oEP/tN83aVOdd9L29b3z6E8/HtJLvwZUTbtgSJUrX6J6YMmfasrGS3KquFW9n
ITf2LUS6ng9Ha4IV9ET6LclHLQ7schMN30cn3mc4kz6fTVHy/R+bgikHezgS2x09N0K65LcRwsdM
nSF4/G5KlZ+2mS51e6EOg6zgX9QlS3NCMzqtMpJ0QXLboRefO/RmmNUA8ohWnGidon3MSzeaeHs8
x6i0FTN319GD+SQ9fKOlTv1ZsUr//RCDi5C3Ozh4CGg3CEyP6gtQoBmTMPgagFA36f5Ii9bR+3eK
pCKd0wO8aNEORsSz3HwBfvNb9tGrlhCuy8sIi6ZqOWext2qbDed/5UmfZsCRG0RZ+eZVIYo8TGLq
RTf6MDHIrdMaB9pmzEAx4Rf+3TeUyu9/6zE5/W+1Wh08yARzPWH2/fTu06yWBHkqCg7m1hMuV6iM
boXAf6ByFw2aBsWQxwZdx+vIJKQNdlkg73Ge9l83cL2SyvOVJzw97XQA/vnDSr0xRIphp9tkv5Po
ClDKJr5XQoZWZ+HKVKEX+CZvwUtQDJKMm6mpia2P4XpPivLzK8ZsMf+FxMTN2ieeigd5gEeRYFsQ
ArRq4mr0JQdcLW4ELwPCAQPGpmDNS+hrwRTR+UXq1ZTKJW1yqiw3wcWu6YdgKgC4YcOJ1TmtbiOM
/2FZCN2DDIH1NLjJsa720J+vXhEtkBfrtJmxyGUD/0rVoFNQhUwYjoKYI/NkAF3O/q5S+NZRqyfY
mTLsHI96STsQEVck/ZsDdnzZiGwpCxcw93BWS/5CUC7mOfRyuchxv51n8mC3RQ7tMcH3MKUSPohB
IMrJQzLRQFo6ZEUA1GaRgE0VxwfIiYkqs9Wkx3zNiCqpuGAtKQ8qtllawBddvBcT8SQRQ3PfTDzy
/bzAk1eMX3lxr0cM2DWnbw6++ERlkJAuYyZjcRxeAQm5Bh9xsfOx/4385O/qGr7U+937oeNTQKAH
mLQTOySV15TJFZ0KTa2bcuI16mgZBT0hQr7iPE3457Eh3FGqSKB2dfK3TasvQnucAbROl0AP7ekt
wVw2Lu9QdQtoH15d/DfDgal9yA3LEL9ScF9gjPfKOoTQFG+yTei37xzUfvsy0wsnyd7hsdo+tJcv
RlFbshdzXCd5nho+WnVepO9ACLF64t/pDqbjGRvLjC4O4dInJghUrp+XduYyhGLMGq2eX+rHWMKh
kVLh8XyKJ9ntxS9zkkvD46UAGncHxTjob6iP5VTJL22dfHZUK9z/xaEvoSSJOQ/KfAT/WFf/wR0T
D+Pf2EV3pHsBE3picyHZoYukLOl7lFxHZw1O13zBytmGjikTBEQB7KeAbrxoFxmB3wx3gYs1gurd
hfWt5ljWKCD2vMjUHgJmx5G5CBJ/o3IE8TMKQelvNCg6W+J8gf33H1XfkStpL7VDDxOYyMNXIGAk
2GGrgeNxgm1Y0wOjM1ykElBfOvG3Wf94L/PLZ9sD9ILEQ0phtSY0wwjuM0gcDmLUWZd9pQ+cP9Gx
7ykii9wS4aNH7wKAlEYCdRUuZMWvL7+8fmtecjcSTclJkYIrzQaFERTDGuq28pbTQY7T3W1yUfUJ
VwOaDY9nazvcJYxQwn4mGjj1CR/4sz6GU0oEuL0GFF/Z4eZ6//2/EbUWDllqmohgnzDsXGymEAiz
JJ0Ro8AZXKFlBQHTldDiYCOnXjGNDo89RozNKYuUVp3O8JQswrgmdOAJHgv/itRLcQEPY/1F8ohX
5g38fR5mML6UMeM85OfZlQSwDAWSXd8nq1f6YxGGHKuXCT+K4NGKy9IOhuy5gFBgz3kJTRJC7RCi
O4DjpBauiMF+uZNxC2q7+1YqsVbb0GxEL0hoNYXPTb2LWoz1fsy41do1EdWBq9FbpsHcr3uZx6sn
ubk5L+06s0gqDi37MSTwya2Tl5GBA8RYSDKMqseowgaXw3rJOYjdAHjpq0yAkgxqEDgcqC++XqeN
IUA9/IHoGDu6FI3xsyMIgV3zxgraQFS2gyIDNhCmHYJwNna5t2lmEbHpww2bIfB2Wh/cBlrpY4Qp
PAOPJt3ZhpbmlJ7iTt4lynacP1w05OAnLoOp9aCxea4h6NHBWB0ohCw8RZYF/s8zxX3r2JSIronU
NpaNeM5RZ0GzK6VaQlnK2I2B5ylbQ400sDkd8ZmBKRwZacISITJxcOIRyTRQxUKQ61DdopDkYISa
P/DYH3npr/7VCqMTvQabwlxpoCzVXKRS+FabJtmpoi/iVlY2AaZKnaWv8A5w5spYey2DsmTAq1k9
j3DxrCkP3tknOsIXXrt4AptGCNzkygaMReOOPXlcrkgac3p7DOwgURrSaJVQu/klGRisR2ga9DvZ
pxekm5tEGo1lwFtJIY3Pf1Xw26cCj6RIcoynTwBuqeKwVYl3JAHkcRc1qcgg00p2X4p+lSeY7klT
irhMTNS1gOsovq+fLHaOwPMIYIEzVqnJMOlKxgIgdSmUoQgf6Mi+KQpXiKxiKqY3Xxmszcf5LDxN
xFMwO/esu46Gf2mFwveu3PAdGrR1plrcLYOEdZfTAqEsqBpG2wbfNM1YM1t9mqGL7ldr0zuaI0k1
PlE7sVEvu1zZ+FX49oeBOkB+zxyAww9zGlXQIK+/Qw3Kn0iCNyc6S73gQ4Lu4qsdNpKgaKbAvKhL
lzlC18GZKNNnc+/G9rYxPT+BDfd6UD1IJjtExeiWEt9cglxwvOYNK7/RnKAh/jouJ3O2EEqEeTI2
1aDlU/TH6bnpKHVEZVCRnQ2nM0THtBqJamy1hU3i9dnhJRDMyTr9Et/O0TiX9NQtw1fLHpYvuztt
gYUYs2+ibBOPSppCHr41bYD+C5zcAjXkqK5s3DfAYcGK3sxgPWGml15sPglS+jtxcZ9qjMa5gPXh
4/SK82MhcfagCxCA95jmhx4pBTi96Gpxr1EV9a7a6bE5/7Iy/wx5Bn/JPJVSmn4AMqLRV8wYS42u
I5PYuNPC1QqsTXhpcOQnHdjOT4y3RcIVzmAKImKdrGlcc16WyhgIKnDc2NvqNUm4V0++jiuTM60P
DR3c5GgZ6QuU/50nHdeemn1eDzXjAFVC+CvSuOYrNHW9GcZypGkKb1dFgzcWePJh/srA4++6jmy3
JGdegXnsCIZNeFwWelIH2S8y58SbV28LwePrLH/Y6xEi/8Lg8Um8YPIC2v/a6KLSFs7UbsCPxy1y
oQ2CSHDi6Vthd19eW61lP3mk57Hx7R8i2sTRaLXniilfANjfEUka2MC3hrraJLmNZQlLcEY2XGzA
zscmN6PDs2rOLwuGh26W4qL3eeGBTpu6mLAA1eslQwo18ARzS53O2GbkQW0yvSQk3P33XxNmPzhq
LBo360kI1bmYn1ePGNRWRo1iTPweDvMWMc510yIw7aPBnIlUdrWJmMaSIhTabkeTdZpS7Bh+58jW
EfRQMcFiD7jNcUzAt5aNzWXJm+YnJtt7qjxKrRVX/9FWJUtGV6KLlYvtZiIWdsrsmBnSw8sWh8WK
c0xA0fWKcBLNSJlBmrgZSoqaVQZ7F4+dQrAdNTjBaWgBtWTkh5CGAXbrd6y9aujPRjotmIBhRbSt
Pz/myEWCEGd9O3LRMCUM0KDXjRVRE1QMuJxXQvNmEcXOtQHsqrn16HoksxDn5xxccbzXHWv16Bh4
1VLhbl2tcZ34Qd87AaUVZkISs3FLx/UD6JpAPDmksGfFuJCba9mxxWfvax7dQK4rcgKc7BG4XTNo
CqN/V5lSHhMbStoZIlNc7g2PfUWUo/kROhjnsX19NavAlhQ7QeGtex79rtPt7IjcTytJY3I2gG3g
6M/t7N1gxQ0/5dsqFEosFpQTAda6qemSdqglrXBXVTl/s4ikpnmXFT05mpjDnXVrfnKsOXgYkT8i
KKTVL7WkAOh0TGoiNPZyOK2BQXhYK982NRc4FJPYN5QQZgOLYDKLisTp3/1f+tQEA8ZykjUzrXGq
fyVJNyr/7VZ2D47D4CAWZAlgxxqqk//sQiAdrVnpp/NvE7/Ldmwtk8/wBIRz5LvMoKoIE6o4tJf5
iJJutFznto0tiWQgd0Bnl9KiheM2rEQzS6fTLg+fy3x3ibLbUY69cwr0t4+oYC+nmTBBq15dU/8V
Yiy7hIAxKXUti1KUZ++0JOWUZ046YwHO1q2AXEJ7R4sCXQizP+mt5PnZLzmGa/vSH6Y8e5QKJRk0
gu/onYTxEA9O+GFQc/zgrvciO0+cPpEA1rIyqd6Qzn4qodDZqZwxvET60SvNPpYeeCTyoiPf6Ue0
/+3rJNfksbs/3+HVfZCaInFIf8dGKuTUrZwXMVNBh5pv6J4NW7+3OG1WSVkWaIMZYpMEbtAs/MKj
S32djHQ0GkrZhsnDu4chwosIFYFOfoZ7KxERw6hdA/6bsb5R6fswOCSMbN070m35WRc0xLXPwMoA
8pps5nScsFbttx9njPiJzUR/zrtqKuQ3LKwOifjVs/JxwVxXoxb9wGHRvMilCvkl94xP4ntplEfN
CBfRb5JMoFe27SuiibteQqBF4bOilIeCh+TnzcaSDbaIplfpVUSdzTmBrUva3+rIVTvsZzf/Cubo
OxFMgclmnAbSEQB07JQsvq/P0rAt+PuJ14/BoSFnZzVFJOdBbtn/wbBFsTZVa5Lq/I5eRciItvCi
qfVx8VV9a2WJ5f+sLA82i3ziXIXCBmp9Bq+zVAzrtUnexSSzwJV+wQITACSK6+GFEl9oNuH7siu0
SeBLgjazZLerhWjZsuGBRlxn5hRnqpcxZcVvKkJA86SOkV4NqNDR93df4ZXe1kwnzz8zPVK2mfEs
plv+2Fmt5txj3kt67TC9iDYhwxMDlIcU/1uE7T9IOr/pfXM//wdlBmJogjqJpuKV17hL68yPp4Gk
ugcW7pFQAm9Zi6LKN5/6F/B5vecaWco9e50uY3w913HJ7SH3LgoMNNKkx+OA5xybXq2IWgjUzsUz
ZeMlfgCBRrtl1IrAcuYaEvE674qPwsyDWLcsLvZXILE+EhFaL6Liv9fwrpFFYKwPIklcy/Lay8UN
vRK+lMcKdGnCl9kfrpxNDimeIS3LRwV0pOGxzSLj2F1QAlH+6AkgX5wTQmOtZaO7xh1P1Lz/Jjkx
CQS0abNvlVj/cliHY6gbHKRcL03O4iUDzoKVliQiXQYBciz5AutB+OVEYbuBlrH+7qS6YPzt5tSI
bXoy7/ogywquSB5dZjiopZBhrYnn/iTBNacC+TvSTKpmPF5Xb5rJEbCFI9n5AMGYUqA6zFI6mK/Z
92mBAz7hFSJ+rGllRzLw9riZadO20n8u9I/tCmdP5O6gWkEtSR4DS8j72Vp4oKuR8w1Sm/WQO6wT
S8nOByg5xIOv6jbwzQKXKO5rvo7jkKzt7mRwnEtS1zOmuk1JVGtwVCWV7KVeuNdHlSVlmsjTZxjB
AG+Y7SDSTukTb/MlZ5SD62ZziL0IQ6Oo9pXYHkcBqxJnV9XYPGHGuCrE9Y2e9N9pgK+9mRoBvl0D
hBV4Fgl4FOficGJHKXKVRC3u+1ba2IZA1J4g27GJF6tw466X/iBTiiOrtJZLKhvAYBxksLroPwJN
iYQ7Kyu3WswhYjqjYfHzPcOW2OMrsFS5T1IQCn8V9JV6Y+HAmJyIugZOFvaeEsYLCH/mbkud+xm1
3R0K0sOB2fl1rfAq5Jr6XBlmYdDkumsLiXz81wGkwcmi6xQ0TQL7LbSBD+KMSvbvs3eFjks7bx1r
ymDz3fwSWWo6C+fy7Q+kr/LXmoRsDDAPi41JCbtxcgbrDObEqjp5kziJvMvLPsTGqr9BV4Hlyg0m
1Zb5hL4uX5EYStPyzzG9+zJW9d1PkslediizcY/l10RZE1g8+RaEr6goFTjVvIDx8snn+O9bSq0A
TYncNnWtiORT/jN1tVjtKYbvQCP3d2hHbtYDUxIpx7tIhA9Ni4vRGdZK92yCsjnNIFNT0IVK7nCp
Irm0PlHO9MTQdZLhpGaUjABu2EaWFhpEdJwRAqgnpfQt/2VTs9q1mkdNC6alV3RWoCsSB9sCrvqn
CgXcTdhEIkwVW8LpDSQ8xQ4JUJtbwtwIy/5wTFOP6DKNDtFp468FQ4paMOjDizahgo40pT/iX+fX
pAxY34+arzQqAdDXbtO1IF4Eeyt5qvpx+7QzEay1ZbYJiaWBf6pHzHoTU3W5NpnMBnsr8yLeb9tQ
1IsmwYSrRDUFfQ+M5NjX22uZ/b4LFNViuxu/YSAnGl/Uz//UrQ5UyhcuOMwHKQLnwRCGbKZvi8Ek
IOc69JxFtr1OOQYdvBheaGj6VGou8aidh5F0LtKi592UZsGVZM/a8YLfFhWDpVZbrKhaHkMqqShv
G9cYwJnvCjDJ3ADNkpVXMJ1Cc4r2qnYw2/oUQ5tKk+GFm0VezmjTYSPjkLqpI4zj1btSmXNYme7r
qAg611WhZh9wWUydxrxF/W0oUrqBgisPetC70QBZ12+BE4xCLfF9KzkHUW7h/HJ2vqOGALJNZtm0
Bxg92vYxCw2FW9uDRwcyc51mkc665pAOhIi0nBEB6z1iKMyw/99q6GsYIRMX/Lg8J2iAEkf8NYLQ
jJShDhL8bY97WV9xU0a4rk9YLgcTYTCrLsfq4lN5G+ZDG4vHIpmHl9tjFdr9StED68WlKxaJ1BhY
kxqEekgeiadI0uSWXJ/HTAwWhN2f5YSJX0NLsckFA9iIICwPSUJthw5Aq1klnREEXfFt7iv95LfE
tD85wqvhV7Wf5ZQ5wWNH+gLi+DJyjwTefAtJHTnvLmUWDHdatvRgDjTufSdCuz5QUfvSYEJYXhIh
NnKJQsBZFQMk9nTQ5AHam4Amdg/wmrpgaWX9QCNHCuRvcamIqXjs3PQwpZ7U82R71grQvaGdnSw+
3j/hb5UyzGe+qTQmNTJS5SQbgU3WDH5gP+r3v4e7HACWUAI3/Bg58Jgx1VZen2CQUXlpDp/RE5N3
KaRl+4CEB6T5/HtxWZ3yiUT948SnkcCcqxuYw0OGTlFKAzb4n4L5JSAcXAqUNdxJ2UIPIkhD2+UY
A/3jQGnKL7s0I/yyVF1e+Z5cjJ62i1/kN5mWGpNjvjvoTKhuV8fkp27FENUL8oXSlAu2w1lY0Zza
xSSXHKDBV4VYXPmvC0Wrqhy637Q/onTZhOQPTyksRNFo/F8iVD4EFX2YYyH1tCsGSPjcW7/j3u1H
8KI54RIX3YYgtiEwl3UuD5dDwbnsHY1keJDRKkDAoOq1kqShBhaF0nlIyo7YNXOZcwNfZtC4oJUT
6W78hmEqj/Arvw/uOCaj9l2fHLmCnvCEFDiTMqOa2KUlJd51kYLFZErxrKspy1mNLGIUFod5Z55N
3avLhbQvxje7gm7gvO/+7Mi0S+HcRT6mx4aqjwROuUSVbvxN2d+iOlYkd+OEuOIUkcI6r6Hq0qSd
hHAP8R6d0DpTgXOx+2zFHKQ+1ihJiqUKL/IU0AzKrPYEEWdX3bwogmOwDAHiHeSs3uNCBbEU3IEV
9CGQdT5lB+mZfWNas2zuL8pducvMC3//BuuP8H7lyMDmu7IPQi3SMP8ZWYUxkE7TfIiXuclE6YpU
pMQkTRanbIVnv+m+ukO2Q4Tx3xfDUuMb+RbtOqqX2pnXrsHS9czAkcLe2kUmgIJzcV4oeTfdGHhJ
wB55z6zzmsV5LYh5Y5kuItgBzIC34CxUbiqa4n8B0occBHla1eEG9E7KbOQXUNQKpHHRP7u7zDrw
U+ZsXCMU0D3KCF3KialXlO/Kl4cRLIdvfsl1WwWXevw+i5RSx+fkTybZLrdCoCCmoBNeYWoYE4uW
oko13R2V0AKizQOSCHP47ai3u5X+NW3B3B8tzvvV+yoX7N/s5O1EaLgdFMEQojfqd4BCUR3ethBH
aHNcfC2wHBWWHpcfueaPMlD2qCdghBkXNTk2B9oSO3c5fi/A4tQuORC3P3olCasur5BSPf34N07l
0y8r46F+7Cy9eVysLkBHveFBpb3EyyiEtbd46f/lE+cxcT3PkedDbG+IsT5Id64+31+IyEvvvrrh
R6PGCkerjyzD0GuJZ6/wCbNxhikh4ByseIoADSaWslIH3nU3bJLLHzio1BhRu7Vo+T7NIKvgIF68
KEzKNSPM5dVIAdyHHWH3gnUdKtOGwKGTtn3B/7mAQTv14ZnXy9VKsQwFxpDRJnRZrbak7bhTLVdf
cWN4Td1fyinmpJMcp5+uJqRoyJuY9HiBAyLLNCxyesfqQJuQajqZ9DqiFx0VXPeQvB2Qay82vU2t
Oo67uRqy6+TpoOOzF7HdZKgHCpFrfBqln3AbLnYOP7AcK5u/GYREFTaln/vAnVRtD6YoBjlMugch
J6fe13NWclY1cw2YdJefgJ8sIfGSh5d75tQFMTk25rP5SooN3U103GmVq5NfHfnseSvpM1E54DtR
MDF93JeaMeRgvwTvgU8jLMfk13+hOQRV1qR0nrawrGF7o3wKij204qNfjfIrrvEW3NoT6NJpsdVa
no7OR82o3Nc7r/CDpbNlN/QsYySbJb5ho9CUWKiOB9aj1yANgz3T9AnGozZBaDJ6M12DGvegTkGc
8fL/ACSoL/t6ozsACHMZO4TZoGwPXn3pF8lQoLjs3mPaHHFogq7iAC/xWLLTmgF5ZsSXvYegR2H8
ABczqG9qDlAQgJG7GskLtvW8kFkyeZwc7CcQyaSzm6nntZ8Ra2yw3+hjizi4RAdNjcxNh5Ec7Cgv
X9HKOh4edPUo5LNSu3sR1/c1T4wupuyx/gsp2mR343FyBYcFpBBNsKBCnbJdYwVHPgSeam/fRb8X
g7ozZiScXXsKOZlDfKuIw7eTg9nSxoswBEn7fbv75F71I59l7Hzh8gOrUFeH1em5WEpYpkCB5MAZ
e0dA9dV6MKHvp6pPLwCovLc4N3kfJyy6CcMUSDg1MAbLhlB+lHOHzGYpkK+v+l9HXTK5pk3DCiv/
zR839dSWImCSTWC13Fn3+0IP2GWtG38GYVdOCfNCiT30PzQhAOeJqz8QC43rpxo+CTEFDKMw+Og6
rxG4y6I0LxwQE39TGiktk6/EGpLkQotYACzQwf/Uqexq0UdGHlHTfkUcGHqDL3dWLmiv76B0I+h2
g/eWzPeiwrmPy+siDqVLdjIcKX0erkVCqy/eXHV6a2GHTFXHZ1kbD/YP9YsLbKOTaa5pmNGaWSVh
SjdWalvWjXqsZ7IgUe1qlmUud6B71Uk/aPb4Jx4rOUbofFlGYkCN9AdMK+BRzEXa6oCtsIRibHWr
KBn8FmiIS/nHLfk3bQMVnae4oROmzNcVRD3qg59ua6l2wj0PAzQiu3NqMVxoOXLbjiC8yFpvGRiJ
UHS87mdZtGGkGJ1pgZh05YHhQEuSyv2Xe1wRzVnu0NumtZXlNWI3FsLjxrZyGlq4sp/KrhrWSTeN
7dkbw0ROl0M0/fpk6cClcUNjGIpPgasO2gBpFai2u8xjeeQ/qUZzXZAWGXyMIgVsqmRCx64DRsFi
FL+l7z5UxM39SYCe5TIZMDkvdDdZJS9evt7hgNDX7WbLy29MfJ//PaJgIczeOP91HPmrjubm80po
eMEstzRqBtFlOFY4QlltIAHqwdybOQDJEwHszubXL/k0gW+0QURFn4dA9DYmKxfnVwuKqr4M/Wfd
SnXxa0fcf5whV1qxE/0MU163cHjs1zP429Z2/mDNHFZu+T4y+ABWwHH/rMZQWCZ0v/EBcCNX1grM
pfvThpSJkCO/EEyrIcpdykkzFyavuRt9BMDdictmD47f61p8RCWl0FkDHZdoRLWseyZAFE9IwVUC
aku8zwfnoKCVMvY/b7q8phOlqP3a+dDZVWQwR3cDusHmVkV6KTYWKCYUVQ0z8t6vF6AHEJpCyvLY
SBOYlS+/+gmRxYArSdiK0mY1OrnpAK+m8o/6haMcaC/8v18Q6kUaaGFbtZ/rETTIjvA30+ZwyIXv
kMe3HLM+YA3G8F90aP+TcVnSeKP3xf9tC6SCuym/glu7hAokbP82nDXPwYVmcAHG5XVVGkdjDWNI
5my9tw5Vyyw9PFKIfxRsqAarxgDQZIEggSbx6XyHNpO/zcsPYPBi7cBXD+oqIc5qEIPoywZu6tBx
3Vk7R5b08ztUO0g6LFP9CVDFx7KtMHdoJXf5Vl9Di0aLEf1memrufKtrvM/kPGXVXA5q4oTHQz9Q
3hckejDSN/CV4i40UetdWUHpBqRoNTBgUZxj6Bsao5qM9LfTaP+TRaZnlU8xTMSWdDBMdBjcR58b
ipxbPuEOsVI8n33k3prTOCiep8lAo2pNEVsTeloH9O06yRcO68iBiViR93zoyGMHrKABIsqJF3Rz
tUAxnzxMD3PgHBFxB9iq3ZDdEo7f4NZNfGbmRA4Wncm86usBW3w5amHFMSSZKS4DePTr8OSWpOXX
9DNMfnhnWniB7XnrIXr57b40fRKsjk/AUv8e/tQQxYzWClWt49oEAmgvjV/Jnfnz/eQVR6W9qdjI
ZVAMpXVcLDvmy9rJ23sjHAMYAKzH1ulZ0xhz7NLdJn8+O167Hic4VKKSvrLqv8lf2kDoxDSkgP2F
Lmcd6gpCi1SmMXPTxX7xufYJQGqjSz+MGRfCeeOq+89U5lW3dQKvm+vmtocSQ4chpzcS2EvGqz9V
3c6TX6njZgmEKM9xqMkK9274kGtJpxcObM9qXPND4jV/vt+kdu/qbu/BwE766h4qZMhz5gGb/ulW
sy8IMICO6nj85qiM/oCXf9+yL03Vwnb4qAJQ3r+wOshVQfUsiN0VwrIpdpDbYzwvN6BZ6HiuDBJV
nDTZIuveDYjDTmxP3/uCyR3AEs30PjESLVCzxfaXazlSONQ5ZENvfdxiLBXFnbJezQ9pO/wvOvfr
1wgZBTU1z2bRFemCVxx/JiePjoZMk5ZLM6THOke/+CHipRGozOFj+zGFw20HFn5z5j5Y1JmWNdH8
Dg3UEyIgrKn8+zhfAczVUpd08UrFs572bjgXtgzajGuWA4O2HIfhEe1U8aeiWe8F+ujjo+zM7Pm9
kaKt0L3lo3nG9hmQQbrh5OVrh9sLufY6iu3+RfFzoNHANBegZVv9ROlWt2WvMVTnK0RYIYQzRmHj
5yyeWnZsaIgrsu6cHOELBLjv1JjaO3RLcHfmybUXjiikcClSMreJ6cFUhoQ3bvKC9y12p/BMzLm6
dZx0zDleMv6aZr0xrpGbPh2pacWMLfCaaMfkD1Li8ELiYfO8a+PrUq2v3dMldjZszowq31389dqq
ZtcY5doNrdApbLkTR3OyGrIz/pYLXSid4es3+f6TSaJIUtC2hXR8XtsQTxr4y0nvBZvKbuo8DGOI
fXmvnljujh1pzzIYPNpzP1ar6VUno2bboOFkC20aa+J2s7S4OfDBW/rUrrfA7hiiiol+O9InkZGS
C+LR2AuAlqsqnS+9bd0jdHxLF5/dkrbmeaOZBFS6J5GxckXBZkr/t4UNl5e8eVyXPCcCbD1H6BHN
CO5SSb+DhQMtuTWJ45Me8P/DfXWH6PF9wf9Y/8dMCDE9Uooojm/Cqk6HAw34O82UInxG+yAdT8bI
VZuX+d0b5QAIQGYqdS4QTGB+9msZnmks9dWjiyIw6dma7/N7kWx2pUL14kBnJuooh3oe5Fr0bTFC
CRZERIQZR0ingL2mIKow3LiL9wrzPnn9fqFjStpFvT6VOQDprF1VxhadDnWs5Bap76KyYlGuXzzC
KeC4M4eQyv5dZQlIvcvktvmb3g4SgosITIUNPLs3DWXLr4Sm1DF5jc8dYNkbs9U909xZXisZMobI
XAjaxLQmGcLFEbOjzEXdqUgutALDbh3iW9ooUdmlY7Sv4G5Gnm/G8zRlaeL1dGR/CqWgHEuwWqzf
fB2Xg1LURhGh30RE88Zlz20pAbmrJAYAk6fSHlEcOWeS990BgSxB8IaG3iMnNqIrJvzFDtcPM6hN
nQrjpuDc9upv6E92f87sFayz6haa1lPXR1cEtXN9nqISH3/VYPPD6kIGFYJbyghbJZgMN8h6VHiL
oPOFfte9Bqsz+TAlcdhHgKUEvNgmUvuOP68ueO5FXpIA1sE8p/P3TO9aIRREXDW240WyVDcpogn8
bzgkC7ETdTxeh1LFxCkbRI/i7GDE/CWtaocqErs/UGl79d1zB7MQQYLyokENRu+/DFVjnW/2pzOI
TI+54XARcKFF2B7ozbzTS3cd3qL2WuqkIUW8kDUrUq8epshXbOUVpV/11jih5yyyxODODVg4/36N
VRRUGPy/I8U8UZfBl5rtLoCvpLBD87t8mwUAZ8uBs2eByrTBFf6V6sBGz1ATeza58YiQ2QOZz7Ox
tdcGZrriETDzrIta/wKSyLD29P0Yw5X2RWOF6//lEWlOjBVPhJtz4SyuB6v0qYFgEzOom8cS+2rZ
/NQ/aw1fpKtfi3kYSlfasNSdA5SRjNeSTQKXOaLaeI/E+B+Nc1vd8orAyqVtaZuUfRfgKl9k2tbD
f0u6hRMR7DgVDsr5fgm9qRE3UzslI0GxDdasYlyODGL61EH4KpAsD8pbYm5+Fo/McnX23ogJVIUf
74PFpNGp/qw6i/deFwI9g84DCYgoK03RO3buRRJ8vFGpkL7NFBDgddbeZaiGmX87+vQPAA0yrjSK
YqFYwYc46cE/UByWZzknjJ9pcecLBBTTGOvrNOHtUr8kM1PZtuNjtbIdOk7XcLHBhkyThErYQ4ER
zmWGzgcKbE4Pa9h+g1+NkKiKhR92xzD1qEds3XQTDHI40OfLt4SF5KJd6v0CVTGo4enMAEWnRh2X
9DtT7I+Dh1nwOpdEwcN1IweMzNQin0JDbXbfMc6lInKfAv6Rav6UzNf0kN0kdLvXX66+PsUdaKy0
Fs8Pa2ku7AKA0dZngbvhOLwWI1ivxNJAy21uf93jbRR4nTkbTZezBE0XN16ijb8VOjgAZhb9lXip
O+VBR8mBy5DDkrTp0Zbe1vh3Q50PDlvMWPL1lcDvhjYsrPUtzB8p+4N/yZdqE2KbAvfNkvjRhdN1
DQecjRJnArW3Pkh5JMPZbAbRax1l6mz8oZldqOUqzoruX7D4i32ZkEGxIzBf3+Z6uYZ5O2e+pp+5
N0SSz5HGFkne71Z/SHpgqFHhfbRhWWPC0kPGt9Ib2WmKlULMSEUbXaEEVuc7qUnmwLXSFqdPBA0a
B8oO1xNw3U5v5C2PLVgGLCH0qPOPPlk95QrCuOpS5aJkXoV+BY35tdgaj+8bL1IrtOhTRtkNHnQ6
YFED4FXcfd3YTqgREaccmjHKdpv1XjHaMkjzz6zB1zXmePxOQifs5FDLbeDg6ODmnBU7U95gGIHH
sPSzqYQ0LMcTvqPx+xFiClPXA8uac19I/rdxP+kpiC5ee/6DjrBXTC2HfTrTtsD//blV0G/Ntgag
t7ezXuAeGFcqVaI46u1tOAncDk0W5vbYFLQHYKMQbjmJDHhSz1PvDYp8+KVz2gKBioumRqJ9K3rW
kUeQwqImu4NmD1Kk6/4vq98w/DRJFRzAH7MEno5xvjq94AjhWOJLKZXy17jHb2TgCKQ9bw3HzzLk
AwpoYYNnfmTJ5dmqd4mAEa9vMwSVkz6n4WYvJY/styfy/xH3Y5HdZF9dFtZ5nU6owFadfqU5eVc+
K5QzkEXLGjX0tPUyJgo45NArl0fZk1Pb5sBc0qd1MpGIol9oeTVXR7qKM1gKaxB5zjYVTpfLdiKi
jTgkHuck5cFj5GxuYqF0VAr/mljd5zicFx1CgYPp0PIJdrG5i48jDmtp1pRRkjH27eNmuWnvlM6a
1v/K527Ar+DuAL0Zy0KshwCifeawu5dxPwZvbAm9pQMGRQIAKflgOANU5EZV8+Xbyo09r3daWb4U
FRoTBcNUhyWgIf0nlLecw2AMf+1FbXdshgvsL/owmCKGKXfgpekT74PzUjUh1HNsf/zekv3Ar1FT
qQ2uupX/3RZdFJJvmziXjQrPPYgLW8n7oqnwuv90/s7ZJ4QdL0QNOnqDLqsVPewCzr7O62QokGcK
cAtHf4S2HxEbn/f1XOqesEeIsdfrm1vZJQXwViPbbWBpdxP3vvBlYdyAU09WXG8S5jBvnbTxc2j9
ATDVxa0Oay12al7j7E61es2ZiNikjUFRKgJ7i3jSxDKOJ+FC0JqK8snkt0MoC/UM1ZTE2gPq4rJT
QNN1gT6cqtpReWlXMbYnbqDBYJtUf8dluNhNTMqHiQ+t9gYyJfudSgUcHIrs/LpEZsVB1ktg6Web
L2Ik6xL4z1xEVWnXrh9b4BpSPWeFXjwzZtXwQMDHR3SKkPzCuXVQfZqWGHYncjl779abHerNtOLn
udIWKs3QXFOkcQFYayHEhrmlTEIR05JEJM496avcGfIT5PgY59hglAK79hpHGUZ/YaiywfEScTKR
pvBDlJ3h6EaWmBEzHmykICzpoeCWp3GcLAnqqGalO+h6gS1lfw5Jbk2g8EWX69w4DxTZsh2+nBxJ
ny2z6b0GuNERSyz2LgcCRc+yje5LVPvd38KfB90xp77aFm8hU8c0/agpyITgFTSf+VzPtftAQJxc
J4p0CZ/oBWQ7oxgY+5vRTaIXl6U1gin6N2z+JADCLQw1L3Ah903CuDESlf6yXDAkutyk/eqlkqzj
mbzTrl1hcunXmsiMUGzf+BzQvFdZAebxuAogPH3YNWxbz1AsUCxgBPhiW298tkNH4VFzj+LuZQP/
5N09bO9faSOG1GGUWYjqcN60JrGUFppOjziravn0qLiwf8z+KCHHJ8s7f/4Q5609ZCISQLYSvF6p
MYVFPX6kovpnwnUMQFs54qTQesW8frcCKsm1HjzdWGwlzsfUnidsFdbABmpo6asDQoa9pvfwbx+/
kgu/ULbH8WlBbM/5toLF6sictDj6tLIwzUE31RYVvFni9FSqOhZVIWNXth9bVBinNB79XJFdonXP
d1lM6uCZxhD7rLGwG09IU8Pr4eBvQSzIaWOAcBEFgWymEOFEkU1Xt7Hre3NSA8+yi1Ve49hJoRC+
USh22t5UhXRUpVvzKGw5kHf2ijxAknVgWSLKZe9T4CRQfrB5WEOi8FUXAmpVaoexSCWYhTZb0GGx
RZ690jRdRnd8oc9V1ygxJmeYlZ8/RiNYEYGzc9rj8+D/YVr7Bkmeu2gop0EzdaJSkA8GTlezQk6Y
ZH4hV0fPFZL+5971bYkPuMI/OPgVu31temdCPBthDBtwOOHdBA5jsO6iMEihCj4DWDAAf1YRH6bZ
kfrZPJn6t12+UOsHEbUqxU+6jqrvT4rJg0kT4aSHIOE54tKEgqOWcnkgkEyP0WLzHxl/2MV1MgE2
iu6uvWH/JhI+Kxgb5MKxOQ9ufBSefKU5VzZ+DsftiuW3rVOSPU6F+HcG3qnFZsiI73q1PQ0GONr3
2DYDjyC6fyYMtDG0vtVL4w2+mCk1qw7ThwisFf6zkop/d2CoIs6U50fLP4iQ/vbKxqmAbv95Wdxt
af8FsS1lFOlSR8XaI2IGZK1jlBk0BE51frk4+tD+sVS6mI00R0RX56Z5kCcFrp9SWLbRTNHvzy/S
FswbpJ3BGt38A3JBXbTGo2Od1+mHmje4cXtZASdd5KJ80YcRRACCPmfDGbB7CvIhnwwjk4lK9T/b
JR6l9/9IEsxR7DYS5vcCg3aS8hC4Y+WmaDQ5l4UyUc69AxEThrfNF2Hjipjrc9Ln3a3Jv7b8w0x+
EboDtvz/8QJhuw3oVqrairzb8SwJga5W/YgMp2IqsYO+JGi8tFEXefQ3DK+f7aoV09trdjkezhRh
XqIJbrVop8p6irUL6hL8dQfpSZF5Y5s2cFZdBKU07iFhIeUjAa4JDhIU3eiz9tJRNHR8vOzpro3N
xA527Hw+9O8kBfObWTJ+rikZk/2vsc6VJbM3WL+LxKhWaa6Z0Me7gyLZZGuOb8fKHvUao70t61Nz
4elTjxbnfVLWyGn9o/58k6u6Y5ELLsuiPA/OqUOUnQGrQjsDBGj/kOb3vAE6IqiiHzf7vLAC9o9u
0+IaDUlxIQ1Mhzf9tGG3NfxKhdBN36giEhb6236vJG4sT8S3GCcUpCxnX+SM3FHayCniJ2guZuK/
TbqI/gC+7yaVppJkYC1U7r50o3BsKUSluw/RLlehDuFjZTcekCNcFPIJsjtJycUK2Ql4+XTadPU0
c65NOVTQsIXAf+tx7CeShT/dARgwImyc3b4y0BgqYRU4yM4PsKHtwqI4Z/nDBnqjE1It3EO2oiA2
GbkeB1i4UBdBYY2rnbT8UU1WOwKdgAsmtcb1YHSd1tm88LKzXYeV/+6cFskQxoLP5sR8s5iENDcv
rfwXgmnXRppmUor5Hll1491ghIEn8LyJfZfGrnEfaUIg2wVwevRvM2/risu5+RsWmqXf7XrqSUpO
cYzxRm0/BiqZ8KCtrXeZVeUS7MgWRRVUU24WxCdDsQ+pX6DOj6ajr3ud3AomLYHy+A/3ErVq0Jle
TWS1iEIEHvwV7t5+OZpcbI8v2xzudUI/rN9j6gNlibMX7O4dK0AHf1TyqAiaUbW9/JjISXX3j339
zQIzjpV6N88gYiSpR0XfZRkirRs1K2HENRkGKrqIazuLSwsL9xX1EuuqP89ewcUXn2/Q8y7AB/mp
uJtGf72x8vNSHIXBefxKFMPFN2plYH5FSAzVVurZE3rOZ668/gIbM3SGoZkIXZW568YB3kKE2SfM
OnNfAOvP6DDZzkVVoXrSY/LgmBE358xiug5+TQWtvpNUw9U7fwNBxk5+iua3klXV7kB5Qyaf7Gvs
VF/ejlQSz6HxhNxpBDcbtsTign3RePcW9Huvz9ioACpRP8FIdotn5noMP447954jBoI2mFOBcCr5
vZXYgsrE8GtNaE6m9W0KFQ0Uq4dH73UgaspRgcqSJXoJZ7Xii21L4mIqckpnw+gV0IsNg3DnMjUk
+LOUciKXrvAVcxyQsfJ+Bur7Q7UNvFG2pUEK5Cnee5R4ZZxhDssTH/FvpR4EzAv1m/2oorrLRqw6
OkeV9rjvEvXd3Ok4CZlLDf4iNkP7V6bjacOGYeXY2ooWdWcgKxv7LaUgkAXtJpISxtjyjUB5vviY
cii1/nRzpiYO1Zl65rnkqwREYJVGZbBn664szqXQu5Oilf3wYP7J/gKN9pq74zrdniGF+hdXKiTP
NScyvrFY6jFn86plHvzdDZlQ80D6PKiC+yOjve/Wri5aHzcPsqCaiy9UOoSROsg4Vc/Q/eluAAlY
CGLb3GDgTcaeVXsomTbK9q5C3KekP/AG4MGYqBInh5FKGZPaDsA+8sTpWdYQWUugQwsFw6A5cnbG
rQ/qO2j+mwRUTFi1B/iE8u6/tTZS1rMAgIaPQ9QaomGycwC5GYUnJXx9N/j68eqwmhI134mmNtaT
HtV9dZ4OB4ztrRbpOuvUXYY+e26RC60tRmsnzXI1y5RQXQidAVN9+LLcJrTDkYcatQq73skgYlvF
XRtFVKQTfIRlXOBzmb1yXEG4u1gZERibH/dTzSKVPAA+bBwRYrPCspK0yYXw0WIfTNnB7vMIjP1J
krYb7dp5Pjw2hylDvedBY8fO2WHcOBD1Gjd88VOAxcSMaxrbVxSkmm+PHO0Ft8cg2HQbJJ499vJt
dN9qr631nCghpP2pmNogZISWtRPulfFICTR58c6TujlljFqvFfaBDu399YPigle0bgCkyLbtqFKj
XgdTVziFkJhyfviU0QuwOG67R+Mp2SEFRJoBI4nwrJkC/bzjmmVT9bVBdg3QMwhdaMuIfqOtElNa
GCA6tgFf/cyKpocmZ6eKUd+ppYrJtoc4Uh/lzVwPd8BzqX1VPDMbLC71fQib3ySibP3NKW4xdPoa
BiTC+Sm7F06CybIRYnE79a6mNmpEG4Z61Pa35fJ4UEYwHtzZwzd6gvgWiFSsPe0c3gwdg/qXcE3s
q5aRd1eohHyQmoB2eK+l/LLVeYVm3xe/ALIWYKcwmyOkVPl6JPgLIKsjc4Tz/W6aKb5K00w4b7Ju
9hCyATNWujoCS68CBoDVwfSKsGCpgQyyRMmlLBjFlp17VD3zg3VMDR+/ZB8BX5woLmD2zZCWwmU2
hwE2Uxpdhd4L11oAovKW7RoAYejd0OhLtdjhjtIOI1GmqPq6T3JxsCXJTZd5js8vIXpMOx/BOWtr
4u/W0ukQsOt4w8gbPfcKKIUEbjbK28+wKsIpHjMFk9i3ERe858p6Ijuhl3WGkvaS/EBe4M6hSBpo
Lwy//ZImJuyq005KLSpr8Rjq+oA91ihqlguyFAwCh3L5EpOV99n/D5PSZo58M306SV228rReIqNZ
ZQxKOogQtM5o0dfJEcGMcjOlJYhaT3TujVDJNZZKLPCUUT8M2aI0D0GdpVyK2ZH1Z841n9qyua4e
eAH8FDMfiSzFl3YhmA36JZmgFcGRXldbqgcbEFIGtW29MiezgmLUBIoJUH8WKTUB8pl+NItDJoUv
Gi/hW9vEQAKoyLjJhrZJmnzyVli/XnAvMnNU1jMt2GQXo5WYRZGrmwXZB9/qmrrwzZu+k1ypEy/f
5lWaLP3ag9/mgvLAhGdxL8wmIo+uxvQvJG1Xdu/08nihl5fNbvmwEWkRxKmu8CzNWo6hHk4Aw81V
qQKuKQjJ7gehNLRCy/GfmjsZtHonShTt8zT53QXsPbqHRFRHxWCJdBf7aF9A3x+Ycqa0R0FFnRH+
uPXTnVuHrorjTeiqRTpbkcK7XlaXIDo39uz0SCd3MbEAAdteYteoHdsgvnQaJogmB27ZXUVag01/
VdC0dncQNWSZ16v+Fci6VlUiCdfJSdht78dkDE5Jdne0MxhinS9sO1XRi2UWByLldiu0roQRoPMg
y2B2W04Fvw9M4x3jl2HduHjrKsHptyLv36oM7+5uncPpCNB51Wx3IB0APvJGGWROMwocUc9o5Bcr
au1yJQ8hxN/ptedBag1PuDHhMJiwYGDgugWP2OP9tr5Tz3jTVFGeogqxozuNKt7tEBkvJ9VZCYia
WTgius9yPugP0iHJeeISEZIeo0Ipc/UHy7YJUNgZrmtv8JnyT3KV6jF+7AkrkBDi1aXkIf2ghp39
wRRKN4DNO9mbkUh4YIK2cEMmG2+dwegHM72YoutQCFe/bu6sO9qQtVPPPWnONdlLTjGngzjToNwT
VOEexlFI9gA2UB1wz/PUOns/q8VZduP+e5YhagK2uNVCQrwmWxy4RvYdveEgGl7+y0pTro3cATFF
zCuGLA11jnHMwBOTicPLSrWSkYb9sCPMe3mhaQwHvqZ8mKrv5FKeNYbxXKTFi+sUyhQvR5IMFyuI
fKV0NowzcfvzRaYBoTndItU1bktbw8BkMxjqd1WaN37/Q7a2AR/oa/oZhmkjeyUzWiHIOAUianQu
xsKKQd5+tlKWQ3wBIcc6sQJKhbAT3QS3FjB8phRU2mmJo4L2MrzIuD4Ke2BiFlpXxVZaE+PzLnmt
zQI7sV0pPqPWnGw9eIGW5YT2jYwzqYKur8N9fraNCmrv3JPVXpVVnfq7PAQEtGuNsV1MyHOS/gTu
eURunibNcFo1zWjtvxxtNql/Q2kykkRse9qDVnI8Q6lA7wIQH0bfkolXlHogev4C+fSPOTcxiIFu
aqQ9TnEGGhRbBHVXeJ2Hz5nEDQpWnXPIqwy+PlEn48NcqDJZerB0aFCOd8S/wGTmRyiRVsrI7Xg8
OnWQd/3/1SiRZW+Bo4SJT7pDza986pVwjHR8TY1CdY6omPn2YE/w4smezluFqMd6DEEKOY3BB855
57mBFI4HYmppSHi+fXM2Kn0UpPSVT3Z2CWNJa9o7Mu6EYXl/yPjEt7S+AZjq8oEzObcdsHQmTz0k
t6QJpo98grhpMd9dSewfuDf8201+GzEOwMo+r0pKuTT0MaSQcY1BUkhmrSl5VHy3caqETUwgRMEq
BF2lV//9ZtIgMdzT0hsOcong1lFA5HgWXXyYv/KU4LYyL9max4dM0H002U39TmYfjzjB/LGRnohY
OMrqPHLNcQ4lNtMY6aO9z1Lq9KKpANJ15oxT9jYoqoTHGS7+/DZ7B7twrS2+BfHsVkws+xN9tJDC
O4ZYbAGEWlFtomVC0C4nV0NVXLD7ski6Iaxdkm+Che1Q/J5t7JlFVPKcRY5qHhSyZA7Hz8jxSIZe
Lu6FSQpJ4Tv8ulDOqr3UIE/9CEPgRQrMREUonchEjGy7yB7XQon7XpJHMmzA5H5VJynScnzdnPR7
s3Ud2+GAs0TZ9hXBx6OsTcdd9PiyBiuq+w9MYOnRmFevI5NvxZBWOhXEaHfcWx632Z4lIxy8jahh
jiyQmlmn2UGq22+6pTBwFlX+GFtBjNN681XOcNFwWaOExjpe91oOHgZuLR+Swqyndfr9sn7qEmvb
HDAhR47BfvkhIjo68K1mI7RZHqI9l4Pq3qa2aWVD/hyLVQCmWMk3zs4ts1z1ITlKLpUxAAWGv0aV
Sv6P2h4pAhobu9xzlWrtDthyBFVq95L0QZWkkmK4yGoWJaVGaTYM0eFDe63K9zw6O/jx94Q5Xwrg
W6XR59aSYgc3v/Tdz857EwLgY36bVDzyvU/rc+lAytQ4ak2NQ4t5DhdrTe7R8yEA9isBOk6dMuc+
aYP5HMYGfL1Oy4p9Ry9uu3nL6FJZEitua1VusV+lh1Ig5gGVt3LXXM1ZSQs+PCh2AdYgEjK5LCJI
2WU72MairgtcVNxj5jN401NguAdpkujJx6nuSr4eZDsQBp7lywnXFTwHMDrc7ndMIICt7JUTsbrk
YygifOf61v4zE6osSMlvYsHCcemwlOKJNfs6/T+e68XDLx8PdtSSzsyBgkiYntYo+cL47YTjGzIO
eAvn00esz7tmRwcBTkw8wk/ESEsrzu1b7JtIZ7ACUXlSqksYrg1jrxzSHRK46nL/w/ZnbpRJHT+w
/4v0q5H0kUarYHy0YsCOin+3Jww0OhqfuRmhYcN9wr2Sf262g0H9FgBd8GzOME70C3l7OZXg1qZr
5Xv+vFJA+QWyq1bZz9Wfe5ENiS76xhvdwVX9BVxeYNBRdBczcqNVa0lvi0n+Be8bD6kbK5mb2v53
aoy8uliCCQHL+wzIfRGlPi1rM/HeqlS05qLX1Zn0P7mMELXYNUgSdPu8gZP7j6DDVIeWy0KlvbmE
W4X1u7tG1FyDhPn5DlBgSF43nfgjClxzpId7OdwbJeTNWLrpa3HFTDfNjXi2/FdZaRYl6WW5l0NN
liEYVwFMEMIL691o3GJuUpMVU0D9kRILGiS4PmemOwTwCnm3lcWs7v1WPREIG9VGA9pVY6+EfgTF
zFg7v+H6XULj8gNXTiXKtIFfvxIfJScOnOFD+v05yjBtqn3K9uf+Kdp4RoGYmh3oon7hBmVIW25z
EvMVbJ7jkgxGZye6j5zvFR5AsdlG6+DjT6r35JfR7ZAs6p/OQUEEb51loTSYeugEviUWbBXD3r9T
RYR6A4yN2dSgDElEui33JHvpVds8gvw6lplWHFb9iGlUt0gh6dJpoKbtcl/DjoIK8aADBffhAFTg
p/xlSDB1SISesWAaSdr+yboxFXK83pk6XEEKCCN3bs/pn+uawBdyF5FyYJxlygYNugkETvSlxLSa
VyjFMV+Selsuhknf0IKVAQ3Rgir1zjx/PL1UXPaSIE90VoH2bNP6TGRtYoDpG8BGhjL9RquVr414
2t6xdxZbeuTt2CSXXJJfTb93OOlUsEJkFgAnTWZeiS0MF7RfZvdoFXd05wTQAEKcZcJP+ALQzUtl
A0P+93zbWNHLDyR9pGG+Fvcv3CBWTw75/3sPFPrArg9C90i3bgpY2OaamdklJXJlOCu+wPFFdwPv
EVRLXwDxjzRu+xp++DDIQd1ndEu6AszDn+XzdQ/Qw2KuuRi4ylv395SKByxXSgS8WhnXKLzf8VC4
x5jcGu+qvFmBSHSuvMEKUucvENZMEBvYKFp24iJUCm6CiP1QGMPGW1Vh4wdE7n7NKPZS3iQmknMn
EZla8eiK4kD/qTAk8BFpFYrN2oTvYd8dh7a7Qdk7EELf52ctjdg2FfJiHuYimpJi4rzJ0jJSwO6V
cYGmIo4eeHAXAr68ov74WUxFs1+fgDdMuoZt0x3nWb094L7wm1O4a5IppBRQY/wM9xzF1RlrBc6B
hery2Gcocod5Esg/Ycb9f7w2Eex9uh9c8l9f5VHAQgeHk7dY+jrWIDR2I0I3L1hMGAYWJw3+CZQj
jC9ZXQ0knc/1rj7ej+vwXdYHL8pVM9KBPouEwl+waidOs4Fx3W+DE+F2EdAO3tFxDEmhLCVLOb8h
tiyVoGfWhWvvMIzM71AhjanFu/hUMI5oaSeLm7dVaOLd8x5YGHuKvAzaHZcyqsFK5xhdanAuN42l
iYdpanc5K+/IpSrXUWsRX2KliMxZKRqj7Xw6frgE0gxho4aU0YSE6tZjwHXotyVOJkXLRhgS1XM6
bfozkqWCDoymSIKkjjVEeMufwwpUPmaViE8DDtRENlEAPjqBGvpuIOiIV8wJSoX6QDPWRJtDklmz
oQ1/tYNwKqvel4iKx9DFIZqTM+aAg9Uv7ZS9E/yipteM6fJVigWMcXWIkSwhBkxt6/C5Zi4dFs63
2k8E5Yz0JWTgKsbT9Hercvk9Ss9v7RBKpvqEBpk/0pOFh6WgINnyW6OvQ5g/BRjEqrsqTs+2Nd+E
jujTQPDe/iINNzQ8M/3H+ZEdA7tT1gqEOAkG1thmetZfLS3OWORwenLOLhk/4FM59CFEkP7yU4Od
pM2yBDoZH65DEy1+ksxCx/25J47xnpSBnqw60NJbauaJA/Ky+FexH9UHNONIhgGA8NKGLENYqwNL
ZlKkRw7NXNq1+kyJiSrK4u3Azun95+tSqm65cvp/EldaGV04V8GxNy8hxl8LMDB2vlFnlgyD/XTR
SI2aTlteOikE5Thy344xcDZp5MkfC6kZ0sM/9yWVu6PvUE+BqLnz0syva3ysRS0efCxS7RjmlVQO
cKX+7zv7nXaeeAQy+zijneKQeJTcTVa4CvHNGFA2+/YmObj9qgRGI+JzomUhPg7A+mSjJqpkUScB
4kMIj7E0KhIwEcU0IJkD0DYuGPnZ5UsT7ip85dDghFZQucnsttdbMeRfR2pO/2IbMnCLIpLx6gK+
I1PuQ9V4afM1CP4qzwOcfUmD0CaqpfNFv5drTl35QMBeqN3qG5ubl0itArBFmKWfkZhRcC5RQ5XQ
B39MYZGoJgJf1GC+5nxMiaboGctdy1egwr+vfzY7DR+m4DOYqZS61L0OY8QQiZ7Rubaxw+HCiOto
I9Cnyl+C6pQd5b61DZgQIlw0mr8S97J3yadOS5I/6PS/pVeBJMYIsasB0U1GV+/Owy0B4LTfjr9w
qimMYtu3AR0USZaTg5DXW8GG1WcIT1OlcNE2XggQ3D95CevlLDa6NAzHtGoxLdLKlM5nGbk7zM24
QIVQG73QpoRIOBT+Ik15hdpiNKqiFpIlcIwh8N7jv6ltqkuEJDhpUHVERYwJeFNhRNJI+nguJNit
9VH9W7W4KreND52Ple2yOLjwlLMsG4I1bgSa5x/Q73nlBssNcldY/XGjyo0g/Bx/1tfXaPfF6pQh
IqKIuMcSxTXrpk9kogYiAol+GH7r7vVFIIY46X8F6XaQYMks9NpqTQwD39N0T6EgTKwAdqEYzDD0
NWe7N64tl9rpjCDw+usSa5eWPXf/C+xXKnTRh4I0COFbI3Eez2Zu8N/gdltHstdFSlQSKd6tDCL5
OiqEfgdiLchkH4/x+kkcH1vvZ6LyBQLLJyOVxlAPQJRYCIIRz/PT10IZd2fvrerzXlQwwk1f00ks
q3gz1Ps4usqOvzUMqlbjhOqi4gPanCF0qKWQzMGHahs/uHNVUFQYRiT3VOvCHNX6aw6IhH126N7x
4M5nc4fWqm6WRHfUCky1Dyca6Uj8yBgeQz3VGBJrUOLuDVkIjctJB7Xfom577+kvjk7Z9iAfuHAC
DjNiX71dKhggGspx76JiFsrVkG5eoHRCXfifWJSCP6j7JOtoBbTOhoHzQ3sHOCAlhkS6BMJxG5NZ
KFy5GQG2iFYqkGMdzrfxtJEU9f+dC43FnFVa1DhEr/27JDaevihCmlQhJ/TqhwsVx1qOPlG7neLn
sBRr5ruXDqsBZ6YzqyLEuaiP4SVc5HVmeTOO18b2rR7n0ZrvuwGajBd1btnh8qQ+2/+vksAWbuZ2
swIEj/QaoWPD+dnuTmLzlllKCyd/bjvpvjxOvp8RvLnMqW6LrboZZNg+7Sz9LkWUOaaJiS1Nqgn/
fzjyZ6z1/Of6ixD4L5xSJEVwlwF7Kj2eCmy2yvTCXr3SAQUaaj/LhrsvuVZQTl0T+8UjnS4RvpUy
60Yw2MIU4qq1it33TQ5nmP3n+gtMx07w6E7q/wTFyp8T120gbyBNxxkKNuUQzwXWU9xPq4GTESya
IIIK+ZOyFw70MVzYlxVfcyivSa9gPSJ3uez9EJiE2JUDuG/y0r/78LJ4p7bd7a+LIVTY3d6HOQa5
o6fYPzKnloI4Eyd8/uvx7RjWx+MQoxjAT+7msn5A5dMkZiDafIFlzzjBvWSiVL/z/K8SKbtFyi36
hMVL7WVKtREXdtNt/xtLlVF6i7jgtEfKC4/OmTfPF9j2wIyYDNU+MFP7DXc5Hcl0pXBlMfnWSY4/
yh5HqxQ69rrRt2VE2F2kWBH5qUq/BnaNCdr37XPDDIJRkJcToLqrm2GMgYYEicoCHkY0sgWXt09l
OXYrkwRVb/o8swO+T2ziXFozDnIzVGXEGkEwrOWsQR0PZi9jGbItoly/dyjAyypzoQ2SLf2+Bvt9
rhGPGPSIBIup89nuAV7YsIxF4EDj/LkihS4md+kwTPNgxTqReQIrKk3LPLsnP7Pp5YirKeZnarzs
wg3qMXoauvypFrgtPnsNM4o6ZeuCnUhY6CPl6UWBl0oeHyBFziYImbltaGq1Urd3CiN7uLXQZYR1
THv76lH67T0/3T47IZ/qwc0KZL2jdXyQ6OakzjzUp/2+TzuxLhbFhMYgnuPHnlrTrjTewxP7+T5O
QDy8cq4pyyVOsdzKfiYZI3qWRgiTHjhTHkbGQvG1+g5Mokt6FK2AQ2cEBtmyKbXHXJL/z42LaC0x
xt4LgtkRG1IU8yxUmZHUl2KlPiymw+i5QCiwdpF9BRn65j6UifFynLTEDNoxWPsgTSNCjZCG+/0D
m3N7VoObXqA9vEeKBvtIv7hKSYogqfsL9FdC9NJ/KAbns4v0KJVmeVgYS6vRw3AOq4H4P4be2cim
YOK262vjN4lo50LweZn+sXUFzgM8AEqizqsfzqJYF/88V+iX4UlXuQxvIiU1xoy5a7vqcTINwTG+
+aLuKPIaZYGPatIWv/zI9zmoNX3TayezIsRW9MJcttDh78dg+u6+NS50yB10VoZ3YY2+1ab642mH
KnU3IgiBK7ukDmdYzoaMcv9Fq4FDdgYFzDONfMcEmLMXcJ41DkNKnfHSO8oMkaKs3gMVGi6neTLI
bYEhCHHKIT3ox3cld4wOUkn3AXgpeSE2LMSgsLns5UTVacLqzxzfLH3PRMDqKqRPpvdae3zruhYR
njEfftZeNiAqt898+6H1NoWx6qZuaqaGzSGXPvW2+S+UR7TkkMfzSzwR+ytiYAn+hJh/vlf5A/i/
5Ff3yK3M2UhMG0GAV1rXwAOUggk1f741ih5InFjRujpkDjZu1Z2HGDuh9g0A+wx/EeFFZKayV7Vy
UF60mY/Y8FSuM79yaI3s/dfDmj88jDTGlaDJN3bGcp6P8/w15by+0gMw+cuh6nmGuIBzXf7dyx4Z
hvv9YVYrZvF5N3Hk5r4mpPlyrhd+b2mk3xBOFfwTAU4wVK5gEDHTwAuilrYuX95TBWO1SuF9v5s5
u2BqFaa/qx/a5VUEShV+liv591t2Mly6ova5DJNgp7U8Ojs0IfvQMZ9LITrEO/qiHYLS7bkII1Q2
pRc9Hnn4k7Y9E0jqbHLx2S+6IyfN0ptJk/Q2uaWs3UNYJivSikVHoXUrrwlyD5bIhvENzzM6IUfu
W3EP9MHNIEnGAABXvz1Rw/ol1GzsZ15OSHjITRXRrOT4yCWrVUAWfXm/NokjFLhbgOaSpxClDOfJ
D1KD4tDfOoNW/4n2aOkF/2y2d4MYRLdIxX9Oi//Ay7BK2VFBdwtp+KCoT44TfdffkMLLxGrUDc65
zSOw+3PRVZkLZQdloBuhdtDlhcvypS/bFRtORjQWYXnWqYnm9CfC1qXloHBnpqhj6BA6wDzInMU/
suMnOwaqBxLPenVa0VNytJca6EFUM58hVwlhwNsIPEFxVZ6ZfOPYNFgYB2nYFxQnNkIGYsyNpf1+
xWoLhEUxBogJz3RKdij7iFcvWWaZoWtbqlG6GakHL2r80ueuz1LcAFDbtrBOOvpWdtUMGU3GOMPf
4WLXPKBCq+FhfzBLJJaH4xB6yvZHt/Lc86rRi76GrEeT2t9vndo831JeeL0GHDmXnYELofhOaayo
KWctwMQQOdtizwXK8lgCn3Pd0ip+gTjKMn2JG5DR2t9vCmRnDIP2awD87O0IdcExuRFRMlBGRrQp
xVgI6CEnfOB/NxDp9mHvhxpQql5eR8kSrsmRTZi6SVDM8TmEY8MrZYWlkaxgi30pw/oOk7rCwg3/
iWYW8KcQ4T/afsJL9nuTYKhlU30Adq3967+HgnqqxP/2X2m2Cl4+mLeA0IgaG8hH23ptSHgP56M5
8q3jyDgab5HaSkOFrJY5OnhVWgYY1lSPrk/AgExayJd4IoXcnHtq9N34OaQDu92hJJVYhFnhDH/s
30ZSBs0y6oW/EoZrjgPhLLa9D/fawU5wFNDtP/cLYRlgjv7z5qxEXi9Yazlo1gMbyef4FKNLkFLK
kKwZu5OlKKXrOq7Cd+kEqvBR357tjMnunBcxXID4BSIKRVGSrps8RCcd91By0VafieAFoodLRm2O
rE4FFdtttFDLU56E+bnwxHND69o6zkJMmgryD7Nkob0Kr5I2MrPhhBdDhPX4XGT63X9ZCIIBu+U3
AxnVJD9a935tuclQMPiETul3s3+L+bwaD1qHDtojtcFaP6FAD+2o76Zzh19PlPo11vN366sYrFhl
ag387KzzibhWTxQAydAiX9a0noijuOloXUVEhWiU/Mg9kI1g0/kAMbEMpdhtD8F1easNTn/7Odcp
ZUuX6v/CV60m9I4dWHMwFbtkQjq5QnfwHTfNcPo6FC6RMzYl/dmuUsutHFaLKQc8pMj242sEc/nt
rYB9/SHr4DCiKis7rsGuy+YsytMDDhowjxkrlKrBeM80HJwGccQCSdpZDrILVTHwHiHRWjlM1QTT
Cc0XTi0X7a8zPklenVLxPS6RThnDsjfHXJ0V0kCxEd3ieLenMbh75vuR3sJjuWAWV8930LAEWtqh
0eGasdFZ7yv3PnwnPGnmOyUKe7AJh5acKq54LNDixGCLzCSU9RMw29xROYVkHK/P8smBTJ13L29g
Ux87BDC8HfHMG0WFpKS83w+B4Y0otLenivWqW93TOJ2UWdz8fbNFDnTiOuS3EqfPVK9aSDXczhlS
ILfyH2Nd2KOJc+K562Ri1PT1Zuf8cDBsiZNfSFKR4DoQxoErD84pLWmgz1x5lRUPbkfkQUe+GuKz
8LYbEdvuTp8D2J4NozzwoDuHnREv/xWrHCnYgCy6aDgpFnoEHodz7ApSqS+jnYCc1exZBiD34js9
APVujgGnSnVFm7dhyDe2vGJLC5wFRAmT6atGKS8Pj/poWBWk+ffQ7OBRk+jq6GKw4lyEj0gBfh8j
HoC5igAAAI+1GUngMXTxTvEJVM9zcuv/17GiYj1Mfy5Mz8l8fMPbpgxXj8YMnOaaHPOphEhNzXyq
O9v+D649IRhmfzpAkgjsqwDVgXcH5uny4OijHwxvz7LUazE/pf0ZgYKzMIbnG8+SkTWzKYfYjGH8
zh9eUEGwIRvbLxFEwPyWN4quurev4ZPOMS1lR37iVPsd2BV/ocHM6bKUuFILBnS+gXtZTo/hR0N4
V38eamZf7uAYRl0zDpBi08dwAcmsBET22CF2t+vCU0dOZ8ifgLZaSFuwEuxrHgZbLDxjlqgN/vRP
4xUH+rL1Bw/0cz7U/ZpuORJ2Y9ZLHZ7pcyIxnZR/H0KB/nCJJ6AeOXGd4LdHv5yAbS9lPSKkoIu4
U1zN3fD4mD/o0fDy5Be2KnzAr0f6188mVci+Sq25Dn/rrQyAf3hXu9H61UwWCXel+n5F4UVn0guZ
dbq6Tk+4FNyPHHr05/y9ItCR+JNDppCZoM1eTUChAbrNx5uUbTL8NM9fjo4EnujJR1iFvOykUG5R
Mf0xagAa0hYXPSBM4vn5DLaNeAHYcJuFrrIQN1sPAztZyObzWHMWgZjimYMUMhEXB50K6WoN6Vcp
r0TMmwga9o/fkdzPEF5cuAK9DxZaRLHVtuK4+WUZz1qVv8eLegQil33/QZHjgwilS3gqLnCL6qJj
1A+QyStFUew7+ErOaRdtLR3vT+yVYIrJuhZXXKe4D2ED/rLvR70wV3AI8w7kslfD3lC8my3ingg9
MJJW9mZSLosP8qREbAxZ7hKS7X4iVODVZLdyT6LSEZnDBWbKX6Ls8gKlJBEraow2DhqEL9d4xiXW
Ih27XLVJxmQRi2r0xs7mqF5v2cLKYeCcDsBY2plbzAKTW4saQagTXO1/aU6QxBzJQ1aI6E/3WqJk
E43UGJ36SMzEx8MdYxEdUY0TO+IMe42zMdZW/6k1L9XrDoya296J3Epf8hcSCLW5zpii9ToNlGvp
rBmOIGxE+y48xTELbSLNWq/RK/otRBkOmXt/oogoQFTDM1Id2EXldAaU2VS8SBNVtmeRMxNiA33p
azwTmEa7Y/28WYFqpGBLmvzEFCjnwN8X2zlycgDAD8aSr/d+7GLZTx3W3+fU0apVztY5TJ04VWjw
NUigbeEV/C2JUWiuX34yPHgbTUPJkSEDGpbgvlxbMoEPRKxDE6aLVpefAiNC75J3pOUJdd6cqbOV
7ygB2MU0KsGlQO98J3v9hwZsveNuCgzDpCZQm5Gq03Wadj0FyUprck6pfR3pVdfVByZ8DwiLHCoT
VQil6JaJS4Loenl6zmHhKQBCq/etHa3J5ILpM3SSyOAbF4dislOnr91G200zeMGZezE7LlWwq2gx
bL91M7b0j6q4ms9e8noCRIUlEiIzdrVqR1bIYY6TAiUtfqSz5Y1sij9DE1Odx5imcpDCCEtMpK2G
2kfYcF+lsacBb+dwMmAcJELS6GO32SXCyF9XonG+3y22FLJlphUUUxH2eYhMuTOXmmR3cTJvG008
YUTamDiIrWJni4TPzttaPlLNFG7+7VwxNticg8Ywv8r6hFhkF5tLe8X+cDOZKB9GzuDT+/M00M3c
CgNL9ZQU3bDVgFjBakmEjyOAcm+5Am3Za51jGhVoQdbZnZXiqM/CtSeTsJJmXGzRvqR/Q7qdUh7i
d06Q8EUwA4Cjtr2dYrvkLjLKCmC4CKl6rBjrkt01STgTOX21H7DV1jtNfPCUVBQLFRHhPMMyWIL3
ky6oq732VC6j9kTU7dg3jzpJ9evUyjTImQdWOg+M58oB81NPGlm3dEr2FfHv8qO5E9CvosZ+lXR3
mOLZY0d/xIbPI2nXD1UB1M4rSEo5FzYjpNL9ag2FLncoh4ndJLtf74SREsiKbwlSw+CCjFXzK5FY
w7xy4J4KUI4UoiCxf8nqefks3irslUQmRsTSszqJLo3cA3hhVPdaU5fgrKmohWuCh5v5mTXdIyMa
EOpGVl0wKKUWNgyl+Zk8tJZGO+pirvBmrSo7AND4MVgE59BzmDJuT0mORZRYugtgcdWA5LlolmWK
G7shOlmfjGhXrHWLD080rvb4/Tni96aGpudpege5MAeyaH3iVHq67pSoJZULDryH0RVUV4oiDu6L
D9zv+lcMRn9hD3cO2V0A+kWFMDmQ0vp0oOx5Uah9OHOAlFeYhpHEP4XnNKpb9jx3fj9+LJMnbqVu
pAZ8UCohaqs3M+Fhk8uLuj5nX/aa5UU2I2oL3cY7W7mTUL81km6DlRrCA40GTYN3fbmUTkCGZLRF
asmavfMOOwjtk8vUE92kSz7agdfne2w/FrGaD0dTsAbU13ieb3/MARn2Callgh4Y41FkyXPPYhFB
/hSrmhTADJg7BIo5pyhsKvyPZzNzXQn2xQmZOrzuju8sG+QbWYnNxlBwPZ/I0qYjBbEZSuaTGI3K
0D6ASEmBumbE9nJdWb4wOjPVZcXI01Y/5At5QOQj4HC2ru68BCUmJ7KI8FrthoUl0+a71DYL06Wz
hcd/MqB8/GdUCMYxprl7WWCcJS8Ly8zkeYE09olW/5y6JaYFoiC9RV/osyr0GLdNNJ1CxlqYe1++
ty+omj21CQ92T2BSlZLLbKf7OBvWsvCogFLjQS5zf9VHfF9SMecj/ZVskM6BlmP2VyoGyct6net5
3BtY91fE0fkzsUp6yAFR6bsurUT4tOpiL/k/q4X3LpMLCphi6Opz4/ExntFJdHf6WhblfnJYhNSe
BVsa57dHYa2sNZMvF7PhMwxNJRv6VSzNQckCe4wzVRS9x6VQiyv8b44rdfg/zq6nD32aPIxY2hXA
P9ydmvx/FwXQHY/1483sN6dF4UjwK0OUmYVt5IFCMfhLUH9ZvbX9EwopdGfH9bCaCHyB17pdHgCl
ihLEDvfrX6+8E+bwOnU5LDPb6aFrzvXkPJhV0i21c85biK2Tqs4VncZZT1pRKUzSU5Mk+BdejtIA
Wkey9VPV9nif06AfQgnD8qeE8jKmGpSSjR3m1FH9B/b4+SokpDh+EvE8XqSvFAhdIrCP2HKPRVpq
EKOEHTIzRCIbbIYLgsjG7+xckHgq3fWkRus+POzYo5YzsD1XAh4ICQy7yKpHLR9ldi5+OMiM/Xdk
gpAtS74yu5Nn91KsbejKL+uR4s1yNmGhhlr9AP+XX6LV2/savnuksRZFqR9fX0eTYcE0Rn11GntS
pWUXx6PpaQrJ1+gRfLHyXQd8sAAiJj6s4yapUhIyAFiI96DAD9FxVevYopw8VhwqFFmmfURHQIkf
5JKt+3Igo/pdX6BUnMrrm8e634vQLRCtTv+44nk/4oHmQgmvUP2k71My+MtUav2DDpaDPwGjrzKu
FWNKCzbmbCYBrJAOhS4lTHeOWuHRsVRzuVIOfyDIkX2W4qXmSnBshiVge7MHICsm+B2pIH6MBYIv
A2rXThqDgMRI9FChMu/bOoUa3QhbM0bsPIW1NpFx9tJDMCp5cgkh5mpqOe91r2/xxrkZLQbCKR6r
h+h2Sensw9UeF6eYNwRg+XQoOVGPQG+Vm7BXQR5K1c6Zsui5ULJmdfblLCuAnmM92dkWKsXviY93
7BNUK7g2qnSDoWZm5V3OkrWv7Fmj5cZltaYydvyejcLe98BIK8Mdf84gXJDDWoRiMeBcOu51VuOb
I2S/iFizABOL7yqCi+lgv/XW4W+RrTJsSPG30N8sQ/9sCsXo1RkOcOE5JIdqR9yu5Cq89gFRjYPT
qlxv1++vqGkCdCI1oAO8nBc02a28pdgnuzG58Lzaty4Ybe8pR6fZwtpjw0BpJ6jo4yuoq3tF4Vzo
wfcNvwMf9aGk/wWn86kT5pwDMwbldXpWaFhX/CyP+XE0/xj09UmgN0wnXlk/KcbjEZ8T1vCwesHJ
nTCHj5g6K9X14/ZWdC4OzIzvT7gAUedn/rWjrvcZIeycU38WOSXJHi5Wqr0TiB00G8FEQ28qYLrb
iAhp4dmpa27H3YOl1RpsrfK9I7/fglzBhdEfTPqLDe08UU5cdnobpw70EHZKJURiWGin5fKZUxcc
mhmNAk2NesB2guhg9OfN5O6H7bA+FuZelU7p1fVU5tTz//+7PTmPVznP5/Y2FR+nZNobDvPlPtPV
iwSeog5QJrcZ54fcZszvJwtmieiWblM/Dje0LH/C8pFqcJBwLcVC6TgASgOPkp3bFxpPxp5OKfm6
3Qw/CvqQtpJNxdmBjOLks7ylfDAWjOHilj/dSEXx/6EYvDNffIVlGMkmmb6nLrDy2XdJi7LpJ1kO
4UfQL8SNNxlcyoh5+4MA7BSGnr8kSNpCTzfBu3/N+wIlKSRGAQUrA4iP910NOu33QxOKxZeC3Bi2
W483b1xBz9NNSbEOFkRva8EMm4J75RNJexKqcrZK+XZyAXRYOkX7wYVlgs/o1WkijW5Z3Sv/BjSL
CpYGIuhvoaXLwxwbsgYQrocKu5ShNcBwbmxQrWjoyIczg4v7KjzFAzVLfn0eQlIbQ7mhHLvNJVHL
HusdlRaLqldnwxpMoa4Hv3414uPfittazpfyWMfie6WKek5gdLSNaP4wnLQAky8waI/9ATP6dIN2
qJ1hvU8OiQMZ165C5N51diCeqf3zk2H0xYT99S1dMBlt+3eZcIqstYUDmxmF64nyXMLcx0deXwtw
XKsp6MbVU1uwymk1iJVWEgfaFKZYxIiV7XenIYfxB/uR+1EhVEXSkQHcGs9TGQFWrs9wYR7ipdN8
o5yx7LVsGlZyoOBPY6ta7Ybg9ZI2WR55fOEvdFJTjNwJqMiiN7DjuJr1MSztCcTOc9Op3llw7rUd
s2/PqxS9m05IA3j94dKCjWRc89H3xmZBUWq9Z7KZMJFc6OEYrK9+NpdDZLSW2Iq/DKJ6CLsW8NRG
eVDTpqhna3k2XPFWRd9CO4m4uI/KTxH7bM7EnuBVFDGbtmsdkUAe3kqSSplqtO7IdbMvQyA0uL3M
W3iDrcSfdBlOmQ+4VwHsrnpD7uBUSIYvFrc2agfUa7nrK1hyS7QwJ0cAc71fISKLQGglwnY+upnp
YyRsOiWk6w4jyW/VKIlwkmSe5PD9FqXDnA7cUscO+ENoaHSBYAkOqUKY3qe9xtGQM/zgvZHwtzLg
pJXv1+Sl96sYtrc/stlTVUa7h/+RI7GV0exDeFscwcMcrnZox1r9X9cO28sCNEAlF4vwyCxO9JyG
zfEA06RIsair0A7Mhj9/wleXGzVyzuimUKeNXeZYJXuTs5iyR94rQlr7g8c2clRzKOCffeQUEFIA
mTl33b0EraqCoB2dMqITSLw87ro0VXH2RaJU30++1bB2SH/qtC7Imf9xPVPX+2Cm62d6t0AnU6K0
8WFHBUAyfzi7fOYSBQfodNLdMn7A+6Z/hmxW56gnBctMg+qXPUMq242ZnMRFeEiBZ9nR0qWkH8QP
NQZNJ5gVBnMyfBZdklm886zxdw43uciNYEC25EizUGpq9cwy5at/viWLcqGXcdSYU7z481V4aDgY
NfLLx17hnIpicCJBhiC+srO5kfmSwlHP4IegJ5l9cBZDbeAzf3NjphXsLT2hLRH59CaOnk0ikCfK
B/W6nQnO3bfgYjP+1GNbwFPAR41JPitUSQ2hf/IpkGoHIoC9APywitTp+hMYQc1kaNkG7vErn1dG
GCUWt/N23jfFkFsBHlAImXd/JikMQEMhms6kTc747bL7uWHsAkQltGAQDCA8lhsOyy2zBc/jNBkv
bgRsoVUpGVMOeHFri//iXVJ42Qf4crRueJXQHKYa3VYSxMdCsgw2/ecvQc6ZtH1dzkh3U764REdn
uba7pp+3iSqqwnX1RBx00QsyFsqcmll2UqMLhAFD2hgDWIk5Vvl1t1Aq9I9QbWCq/R50XOVDHGL4
wrwZ3Zf5YcWjFwbAmF2PPtxc/gEFJSZ0l3tKJzBZ+ZjHV3pssBpnO6n9E9FNU+JqA6Z1qS3pPdTT
OYTh5Pt8cceKWVZy5sENMjcWA9yBNfpiFJNYklb/lyBbI1VPVxsgu4wOoAoJgqKoXnGXchhTCOnv
DyF2LOUNzI0wcYsK9UDUiiA1EGricd/HGQkATOzPODN3nIZN7+uywBEiYtY6gw1HpZp1V2KcPINN
PbTLpJVkTwswYwRjVKhN5i0xiS8mbkSfztFVeUQbIN+8FDseAIweb8b6A49+oAizhgWpurNEySHF
kyGsS/rsphwuuvS+eIc0bDJ7/zUlDGzJ86CfCAD7dIeJI95BcQX/WspbjFOc7RByEXQwjUMomOCt
j5J+Ma/qPNRgkrs/fCPjQLZizt90fV/vN3Kg1DVBI1tyNbDYj7VSS/QK6kjgiRSbhJmHXJqJEXHU
mypuw96X5Tl73Gq2O1+nshb+pdFahAxwFt8vHWBzIVwXrft/eEiMB+//ohpGBlegmxYRYFs/ki0X
XbxgQA+i6WfhWClz7PphzBwiSyFBYgnVSl+fLzczxXJxDHsnzy78J11yeRXczZH9rvJwGCRomfQt
XtAQhry4ju1GALqblQb+B6LgnD3z+MpMcku56SvX1U+yeY8mtOSHYjVtgq5wYm+NMfmE6i0C6JDj
ZQJJESy70plEL9F03UXV5tx6pba+eLiYyo1FSjQH5xXgN8sQdoDU8QiIx/iWTMZKrPznvzJwDuUu
ixKK/1JuG2yX11fQ2mUloRZsoSSSYbqeLnJdCuk/jAxfqZBqIKE/HeuOG63R+9e8NFJ5sULH440q
WSopWut2NzGhFChvnbSVk/Xuf3V8CYe1aDUIu2sVBUL988P26ewzHYAL4KXobuM8WxCQj1BhDhKq
SSJ1MuOpPpF/KF9VVSdVl2qhrmuJXSpz6TjJDmRtry7xMlD4ALQcS8ykZpDMG1NAozIIA4YoYWM1
CzHAX9wX4zH00u3mFhD4oyNAb3ocTxiPQLQ2ioj+3eb+6aXVU7SztpRx9kpyYw8v16lx24rsP3Um
SJ4d+xEQruceiXc/DcXaDjpVBV4Xva6TtAt3MsBKuyS/tV2CAa9KLP+PX+PRW3F5fgK4Wwqc27Uo
XVYmwuprokw5RsDfCH0fr6Avp4wSEeHNlJrwgTb+u3a86oTrwDzFgZKPmmQmgqbEIHbkG0W6lI0f
e2//c2fI2bnZBuKGyKtHr8rUvrJmXQVUe/ZS/Y8fEo0exx//JiDyLUWQp41u3wt0m6igs77w9viF
KhFbbHErHUd9IYEBATXovlFJ3ggKxaSqM4YfY1deu8pG2LDoYCVbIbRPB122/MzNid6HJ8LtnxwY
tUoLZXm6OVmgUNUxZ1fUGd94H/loqJTQARnKRw8FZokzLp6yvtVayRW3Jbg5tlNb45XAvGbD3TVU
05wCqI1tJ4rLl/ga7lmaEzuPO2FP0uJh6XaIg+1asoFLsHzQVynC3xnciU7vSEiQ7H7jeQ7BfKIY
Q+KHXAnBqeXjwkrAblkT3wwvF9gpnmYxEwS5Rc6o0XKP6aP3jTlvwpmClNwGQWK+V929XKPMv1MM
e1LIsRdsBb8kgZegrthr12y2105oaDEZFnMUbzV1F1P5G7IozbWZSl8CcMwKdZyDiLvL3zxemmD2
xh8ZsP2/NOWI7XSa40hT11V3s1SeTduxyPE9WtuTD2OD2wh/uFBhwl2gecYu/Ior8x8wHuU212pQ
hO/9xvrVdm5DfekOPbVDexc49H7VwjSfXVVI4iLOExJmpk/pioYvPiCfu0zQ/W78sye0xju06M/0
jNXQ8UuEODCTdYFOQDotsA/rRIug7v7tBcTRsRV0Odg9uVJebgIZ/6G71n56A30XhWE+dk+LKe3R
IU5VouXMUMKBtGm9J/FSWjxJp5RlXRHUEqPsCj/od1PG0hqX5P97tq4Jgvlejz/Yap+yEmFWV+Ri
IsfCUt+7yXzS9U0KRoiIrPZ+FKTgejjVpIj5DxT3nQd7NMArZtTQW8L5KQeutjirjskws3+yyOUa
Lxtq/tNu4MFKNKqRIhRkxNMpIFFPCGNHgdPOpR9qHT66+WkxV8ZW1u994yLqSgk+fG2e4ogzKKGX
R7TP6JM/alSERUDpF/q5OZ62dCSwu+Dz3/kq67Rzz4kraoX82a4chUs1LnGjQfcwcj7ETDuj2EEm
sPS+guY+KOv1rQSdLAHe4gqodKmVg4q+7FR7jdjUVJYcdJT0/oD1e9dB1W6xihEunvFOptVZ779l
nI47L5g6tIJVboCvTKn6laf+ln8Jf54Zzid8ZoLwQPL2nQCixBvl83QPlxhWzjstP/aL/5Sl2ega
2AY/A6nY4Buf/FfHW7aPZaxzsj2RnLiUYJ57Hy+h48ed2SkdxkjDA9E5GeqN3Lo6vgbd9ZXbYf7t
mHQUvX9CmsURpLMqEbyz8FLpycGeeRGi1xtlBD6j3MUg9Mk5aiBNBQsaPC8xjk65EVf/+19YEmJJ
2aRWx9d29s/8OIDWnkzy6eC9XYi0Y5ZkRXlDhMnIAAv2Zn+FUQKbMq32LLNhPYPFELlouXiJy2SN
QeBSY462W6tN9GKMJ+CG2lB5Dts7cfG2bqkAM2Cw1WBKGsP5fwd+K3XuiTVYf4+cI+xNaeT85CDB
KIu6L9jeiXM1rxwc0/PqdtigdlhVUT1PCSDtvUB6LSXmPcKj06xWdr3JmAIL1N4RDZmy0Uy05bms
oWbMJ86S/wRSjwuu5kyvjaHmV32HWlVwvM8NlmALnAY+BcmPNT5gJu1DYaE3Lr0f/xCKGdOE6zLx
hCEAKIVPtmyAxvzP72H221gImAXzghoWdv3l8WQNNpx2xM1QSzMgcJE+9Un+Vj+ruzCpw4ucwDKY
GPjtl8zvzGHNo9o15aSUDHiOpKrYmORZFML8yVNK6r3jauwfR4hHASXYBt1cVBE/xKknoKDX4U23
0BM3SPCX5tOl9UYc//VeVwUpg7DviJeGiIgD2C6dErhifIcdKofhej0bfM0kpW/OjCBSzg3OXOfX
VjaPQbI7P2V79EZVr/eLjtB8et2Drq2lQTP2ZltvoD6WGu0Q1PPYgbcISJSoE0Dr+wh2luf2e1hF
NbQiJMjjfkkohFTSr8n0/2lCfAaRx5YbgaHm1oPCeWFObT10KqFq0oRyGpdabGHI4jtHYemv6bc3
PTCGc2ZtUXjZatTJjYTehuwmnmayHoUjL7uW0oIxckn2oxcYQu8SL6FoOunIUyZ2fOPJWXMvQ6j5
58BLQ8EZ+TreS6Vm/Wd5gsGFIkYIVcxWhjF8nS2hBGFdrdPA44oPF9I2zMNDeMtoQPO00sbd6T0F
HvICMy7+67Nqg24g2ZpVbr/LFomJ5+FxamyocdzwhOxEKlnzZoJSgsAD3OW9SobLwqmw+K/tS9zM
dHyW8oMqyQeiLgAQ1vNfkzbf5HMiuonbGmnc/KefZP+T0TBNTQhAbGEy3Hw46bcVgEPVKRH59AAd
0v1rQyQwPfIcoGdKgDSdH7Yw+WLmjOjMAVWc1i9zAb52+jIehi6iyEgWxFjgOL0P8nFUpzJHXC0a
7u6NGSddkdVeB9NzE4OGPPk+szAs9L23Fbi9pwI1r/UT0w1jiAmVzMFNrWL6hXsGZvt2hk3NLQjE
4fX2cGRRCl5/q7MB/PZANXr/QLru8A4nkOrw0WNGMc9sdNn8OGum3gU+lw/gTKhn0dBG+vCmDH1y
rm1o2i5x1hnT+icuJaCMqrSmnaZdoePHSn+2rUe2lW+ydHidXG1njtZBjocktJarX3BZapPtPa6e
5qgOhTpRNwF+Y0BWYr9WAJ7+WryghwLkWjnF2KonSHtvRxfk2dl6ZI7/PLygcYNrk24uACnpoRVy
xlX/Vu4JiHjBLY+vB9PYrG29eLkLLwLS2GpllwU9W3qFBfBB23hHwhDY0oOo5Cz7vea+KFOs/OTA
ojyJvnQ0P6c7IqWA6U6cLzCWfwQVW/QF2o2TnfonBrIO++DGn48WDa9/w7zZNtECmSYUQ7oTpAP5
KxzOpvWq8C5QAWLAWcHFG75ZiYbPWeboN4P6HXkZFKM1xltqE9p+q9wrEJ8Xxk2V+taBnlG9qBk5
q3t/mkPzTUB1eI/JQVXEWXi25VmbP0QfGUAs2v27fRI3OjIN7P3P6uH0upRWsJMC9073V9NZ5i5h
Po5oFiMAeahNJAjMMow7F5X5bnGnSVcc/CzPMtB4Rl4nXUtLPDYEikFjFRTJMIwBrD5/q7AGNo5Y
8wzPMv8w/CMgPrQHjAbR0xnvIf/2PK4c/f0evnx84z961qevR18El4XhiWCa/t4cPUUs7QtLY1sG
k1EBIfui7qLyTU8PBgpCj2uQF6UTpCc5CuKInMr2Z7+230IWSu0wBpaqMwaWLjS9xmsMkank5KzM
dvNmrJ1BtlgJlXCxYRIbqJGw54g/mwQXsy6hm5RHB1mkOMGXd6rMrt4iPTLZa/0DTc9B4Aae/atu
UQIXzoHOxJkXT4lYMae1qCH2+H/5H4YP48jRVkGeEox3qQVzzs3M4yEmwCCwug8S2lu8BWSBgbRO
+IhMecClhjeD1sjwJtFlQiKQ8UzOwJpbTRki2KvIgcjtj4cnmlwiZD4stfMB15+bSa7pGLlIE5gg
MOJclEkB/qSZMbTc7RqnaUjOvgpTj1we6Igy4ZChMVFaDHqNWJtx9BqqgVdCMA114Rg4q8hexEC2
eRwvv9K5Os5mPxEXDLzdrlMBsjpO9g8fD/03uphI/XTPUfG9VZMIW9e5aAfr9YZgcbsPkHKUq4yV
0QCJtMqaPJqsWKrck1I5p6Cm0txZtpQI/dfSFGEbn8ucVXutWJNK2oHR1KCO9cSLldco5NLyGn8m
nLbt9CrIyI9lU7618tjAcSUXtIBvKrm4oAjeWDQ57DIJ4qFb7iSsaTTHfquKLq+iFExU5mderidR
2bbGzV29tl2etDwV3EphtU5EH1kMpjO7tKl6X+JuMqWmOYOeInDLJGlISUQ3ivbsAht4MUUVlWlP
4UoNY7ZNLQv3TF+Tg6VOYSM/ZkfDG9S+A89+lC0xkZCmICDdLcfWnGu4c1v/SnVDGlPAsAHnn0qw
OhBkoP4IEXI6rV6G239JXyyM/R/lG3oprPW/Yz9ZwnDUoofMG6V0mrPqNj+03vMfe8a7pMhL/m53
EoNZSnpulNpvO4zi75RnB4LXeuV0LXK6jo4gto7GElKSWHvoHD21bk7c3qAQ0wiLMdTCFu7upXMx
IKNZ/6KQSNSbjDbcY+n5OMqINkjm+n1AcWUPeNTwyQMw6hRot7TdNTBr81iavJTiuc+0jHL4nIzY
y5EPcNV6rVTpGuaEA9OYFAgMg6cs4ZCjX4fC3rUy3HzlBV0fd20ZFgbs++a6dcF+B9Lv6MRrYh+/
VsXQjyr8GlevmUh4x2T0dQQ2htiCvtcLIaZv64bjsFj4ro0Cl3syJ2kJo6I5+bWjG4K+EK/lReg3
z9SqRiRkUFi1G9VbpZhFRZhHoX38A8LrVg4X//o1tL8wOpYxi5ZKigqC+DkK0JJQFqxbsRn4EDcP
soEDuWOpU63vkKJw5cN5vkVaAbGng6yXlkZFYY04cfCXx5Z1tEqq9U7QllT4WaUvD8pHH6c66TOy
JMjSTl2rbAL5YFUidcdnB9ltMw5njDRFUCh3TzBzyoes0v7az+0Sbyty88geGSU+6zRgdaXx7RJx
zJzoRrEV3BuA9KbaL/jnfxfEZSO//W6yWpx8PScAsfpUDtddfZSRkGKAmU+Fgr0K+HwdsU49gAcb
N/LHd9Dtk5JJaEalf0tsYXOPRmpzchOoX7ebSpWbxcpnsBSzzZ+VeVuIwzgUnROwjVUw/4Sjand0
ALMd+wWBxcbzMtp8Pl1LJ0F4Lagk5gIlrsDOcvKzg/0XcSB2jkbRQT227p18sG6HnDD7jCIKbfbz
+BcKdi+E+1Jq1TxEu83tn9M7/zchHcuQ/+nauMsTrzvTdU2OtSEnNP7mLwQqjqyLtnalFpO9+3/c
kXPysKEj3Pp5VRl4ThMEpn4tOcvZoQP6URGkY8TGc2wdXXrfjLznXySVM6A4q8dHu0dV5a0S9v6F
0C9rRLOe5+wtaZLmvdrPH/wMby0Q+E1WypDvtLRMJzuf5QWgvNcbk977MgiFYCmc6oIytK4SyYWc
2pu42Y7NUxkydaBHwZh3/BUP648iMXHdG6fsr3+x6/OKcN1A7A8H8c8emDqbi84L1dvIbRuNg2kj
0PJDGs8B+VfA3Pe8Kp/DWEutoDK72R/X6EnP2EGSc8Kr9N7GK8vhhFLdPKEJ3nop3Klu7HVvZGbt
cPW+J+L2goNEOTvXDIqQfj3XmlSBjxe8AF67RKMSbQENmi77CMxbGDU4v21CgYgsiZTLnOEgoosf
EFhaNvxJ6T/sUr/pNIWfUtKo7wORMJ+Pzi25TedKDDy2vw35iDwwoPSFHAgZRGN/kwNLLZbt8rTT
2LqjtT4gE06ezKRIcBQVzRxCGrlxU5b2KcK8HFr+YS1OjW1RyM7gTE9NgSverO3ctZCuM1iiFZ+r
GfCtClE4qp7PcT9fB5RLkRJSpe/01wQi+bO6Mh1EBwQz3Zgnnl4FWgalb3lce3RSbgBVW13VT1+u
FI3AIZmZVucB2PyJ8CHjynZcgcPPCoYO4Rz+NJIbALfXBjTQhs/SPaq0tJl1agoyfBCXs57tPoEe
G65t8j1+zriD69t75hvjMczDjuXbxHcTPTSvwkND0AS1zA7HAlQ78r52X3hd0/ciXSavWOYhWLDD
fRv6OpGM0hOZOlmxEuTw9/IHkAGrGnXaqZFF5urFbszEIuEBoCb3PQp7SDnhwXPL8VAWo112i+rQ
X7SbYYgSDn/n4jKwUkh120B5s9KgwhO7Zkm0sTnV1O8rfI6X6yhalf7DC2lyx730MhQRqaqBoTdq
7T5azlrk/vRz8MFM5H5u0UVsa2y+kkG6BILieciJSkReK9msE5whadbMrCMBnKvW2M4d3EEgxlGl
W+/O1SWX1XHQf/rTs7jM3TvMsu5lkGmnJ2Jb/snEMVMMWUIuQcerPpPhTsbgt8Dl6XrdmftChjas
m1j+rY4CPs28ilipLImmYsYGSDFWDSRwQ/VE8MDOtpK4fF4fNUQ69aUjtcaXCAIZKQUJdnSMyiLU
Ng1Obhyk1hhdLbqtm4qT6RH7t9DBm6eWNsfbaZMp1de5Ew7vdpbZ1aELuh2Tu1hC+5Crqq4HLJQn
wBMdy4ETz9ZOEpLFViKpf7vasnZaZqUoniUAWcDMrCGEKbwAC05v2KgdJvjnkk2bN3hDSnNijWYb
zcseloaov/QiRzRrsWZz4ESGn8K6XDnJglEz6xwyQ9RwH0EMKWbB1HfN2hXAKXbzFCkCUMQwWtA2
GBrAS5ximp34dT5YV6eBhYYBuirOFF0TEc97xaD58w1veu5uK13TAYEk/fWmWGx/gxUksMuDEZYT
IUh3iAAxM4apQe0bFiL8rmsbdXrp9zaO/gvMe8stj9us8dqBjccycPlExrf36b3AE73+iYnADtfJ
dZh7Iukji0f6w/msT9btwJcPeam+e55re0JNORTBGL3vfeOClrgVpZHsHQEvIistRWun1SIwh7NZ
bbq1h5OuDKuBAHmPJ/kqqTMFgn7pP5NaZtjcL3Wg2LDPuqVeYcUkgjFIdn0fO0YUKMlq8ao7ydEO
YtTQ+fKZ1iQFH+HiGW+Hp+DZjoJjJtNJE1+jDjAoAa2vCJG3HASehnp0UWYUWxVGnNxe699n23bW
UBzevdrTRzWGV21YYZMhFMNYeqU6+toXrkzxLn2nDlzEOSMMVysglmV9rZl+s34EfH+K2k6I3lmh
lrSfdDmntti3+gcdxDfj/05b0sQQUcRizbCypVJCnfDHbEd2OXe3iqpPm9IyOHFEMYZm0AEaiPX7
vCrekKQo/K9whIAxSx1VPj8sFdYTqQ68T6qn3OcK+5ss5IdhcIcXjpX2Kcb9nTVERf8Cp9mvvldJ
BwA5/77AYswNJOr6Custcr4QngasTOcTPzhyWLzRmTPj9ISDY1ZBKOsHmHroHrZFzB0JTGL+PGd4
TioGbmbL7UUd49PxfVmD+GN73oCv/WwD0IZC1XOSQEf6AzBqQB8tb+4wPJmlDG5/zmQ/TU66WL73
hMPOzc4hr96G/PUMpzfX/3poVIvqCbgmTNLIl5XzuLy1YLWoZW/3lUBbC3zfcjRAw6JXsRtBDkoY
hAIOWEUzR65EbE5NCmxJfa23IddxMYsnlMACk5WBhX8HJrD4+/OJZKwpHPywjzJbAUm1eEgsBfZt
xj8pojNpD6bfN5sbj9DT+FATA8P+dkMZ9Mm/DnvlnyGMCGP9B7H4kdB/6dyqjM8RaBfEwZ+MaIkI
/m5X6xCI+mbwCB9Se9tK1jpZnEa7bkZhxrFh9GgdUCrgnYJyTA8CpXdPEuO0LibL2hZTFfRQFMxy
5Oc5pM1nlvKv6wJYkQ5SfOaqnU8gXP9j0thkX54H8g4uydV7Yfx7sSXlZQ8CcOiWBc25ElX0EZlO
Y0Is9ualUB5x5HG7OybbSVsstjy4iRA0sgAZ3KRQZPVbkWsWICuAex0XhCHsGcXWeQku/FfkLFNg
xUkQSI1w2tfQnH5VNKDy44qELqCqvMeQDE3upIY43gIa4I/khtiNfD0/s3o3kkHtboDbArEdcyc+
WdbYQiKo8z+9GaAhA0jW9qZk6Jlmozpx2pN8H/TlGtnIh23A0rqtUpJTEfK5f7BqxAlq1bAJ7muE
z8gHdnhj6zugoHs17pdx92IslCCBWKiLLZVgL3/lHX+N5c/WiHRxrRouFfQZbm6T4cOLwmF0Fyqs
9YvVYPbGEmnXm34vzcn+/vV0qd7+BUGPowhavcmyz57aV9/LUet4LrPA6ZcchWKGJtYxQppan0yK
/pqhB3d0xRMhV6zTw1P7h0PKEk7Vl04H42hYnEqsQoXNSpJw18/icg2/lUMtLdGyHhgujyx3N6Sc
LQY01XXx6Bs4v0ZDZSJm3TFkU3oBhZdzTHWxiBr3NjFoCEOiqAnucqNuNaBagfuZvn68z7DvvIAH
oyBdo4yPtesok4uvq64mn7aVN1UJouHxq1LelGmBwdFnKaMwDRQTBC9HZODDXcbaVHFNIRYRV7Af
yQog7PVp3UVXFzThjpiVoqvkVPApkUMlDJZmkJ0jmluAA1edAm5dYcTkN4g8VlymRxv9wb1VEaQt
OGBi7GF85v3LHYIP6dhw65ylXoGfsDEzpCCLXzWZI99/ADVEkJESfo8FAeHsDf9cuo6cTW6HukEg
9E5yqKJFVFv/TcZly9Qas3G+XTLUBlcxzS6udoE7j52hYWJSQ+SYbUFLHcFzTgujYVQujq5TXSIY
cf/C9SviGR2TYnAnFJLzoWMA6AXtFW3Tg2G2aR9HwVM7/VBzlWTZCmmgAW0T7eRbA/fOFGcGFKYx
RD1Ic7AcelttQwKHrLxo78DqgiP5vVdvNmRdk6DfU1JShvcQgBWpf7AJzcbCFAkvDqYDR/ZU7roQ
GFkjkVQ+cQ1Nu63k7u6D59yvQptYCA841feybITbs00PStfdlcdl/3ndHm51ougS+/7UnvTyX77Y
Duy3oTg/CwRwOHJmyFSZZjgN1XX/pJUGROUMyJoCtzxwizkRZ4mL5IRS2Paa/JI0av+/SnVeZvvq
x8wtY++LQ4Orlalm6bBFkGLzSfikOOcXRhKr70YB6Ik3WG7SK+wXgP7l++WVHix8adUVY6cD0/mH
iCZ83wGp76KqQuKdPZrFodQjHQwEvm+FjRux2DNng8/K6nFQBa1HaDxDSZd/MKf11WNMVQTpFj4i
/fN+fj/DTYYqrIhSnXhxiJpaQXE/BWJTdO3GlfDwmyzz4iJprAc1vVzhHCiPHKg5cg5JsBVrwIb3
7Jpj0VWccgDsJIL1QRxf7Dn+XAgConPeKwTBDDmZNYXYeFq1/HregBndlzFNHhegLH7Q1xMXjAV/
vNQ2bgLsDu7rsifBh/ocPfgxQ7m6xQj6e0nLl8jLfed5mNKCWr1W5Uzm3RCa5T7GRx9tmTVfIl0k
FI579ERsB7wwdogzsq8GSsM/GDmOBST7c3eQQXX5XvC2Hpiw4lkktMEmyP/P5YLnO/qfzjLHy6Hd
40Hf2ox6b5YgJqBeoycjTqpdjykdLKEXGAw5kQEGVosiHpo2l6nlRQeQJ8XlTMQajYciFIDAd2eN
R800HmWjhr9Cx/rkSDb/Uy17mERTjrpYehKVkawHDGNCNf3tXNLu8yLproZZNa8zxDXLp0Zqrpyu
F4j5OGsDlScrs6bz/zwhh+vwjShGygB+kUYKn7HRoMBMXGTQ3kn28pOdrSxX9wH36o5mMecK8GUZ
6DVHfmeB6v8YlzPmJAdnMX7wNzzsirVBMqigAgaRFy1LpC3AugvL4ii0Mjt8MoYYdMcFAgxeTcOF
SE1HcCkm6yVov88LkRJ11tXEaiYyoUjBV3mFbZlpbY0LXB0QJQURq8Gb2/mzK9lpTOuykVHmHhzz
uoLbhh2JCLb6e48nrtA626wqU00A57bcZW1SUzZy9mh4IxMFQj+Y9+xTpeIQHpTPnlhpUsXHQDJq
Xjc6tI2rqDQ7Cl6j8TzPuI0ZvCBKPrY+spOZMjK/edRu/DnsQ26palO+AvDSjk06omkDS5tIEnHI
YwESHB5yDyUapAL5Lb/LoXWI8EN9bpR0Y5mtElPfTVD0CBjwyCmuc6f3yzCNlL9VqJYF1nx0eTNR
ECdVb7kt5egLYBkeJR/W2jVG6uQR1wYs0RPUyT4AaAZlsSCgmYEwB8BVlTpgI4MiQ4aTAdTSofoH
EKtW7ZSLYKISP3i9gfED9fx5mJ64HXCvvyBsyIASkDfCfu8SU2rI7wD2WMca7N+sPoHrcQG7solV
3tUEf+BQ44TJ1ZP8pDTfYnn7YfA4KeZXyXyTYTfXHU0Y4Pc0jOdMABy9YjDG3vkxHfB10JfOqLHx
RnSoTDGTmxNVq8FXZx6SLjAEed/GUPSasoynAv2Su13ATEKjdcZoQQky3Esuq2cSX6l8SGMirQ5j
b8LFz+Qme5iwR3tVhol7ULnid6G7uGH3VasaXYmP0k0gdGrSr9jw8w7vxReG3MxrGPuNKzHiiCxM
wEfP+HhjdSLkrj/HVksjYNfKnrtxdqoGQolMh1MoIK4MTMlm/D4SqwRHvBKj9ncc2yAAWTqfFGV6
mexx+9b1JwEAmDSJ9ys0ij0vU56FzPHofftlBXkeGcmmroZ9OCz4CyjVb6bKT2svpXcKKSq2kn97
g3iRk8tcq21RPwfnMZ82yWc3WEI91+L/kA+i9bfn6JLuvj3vOUn5JSkPUnA/TELvUxlXcFoiy34v
DyrCkcqSweBw3ovBSGu2MSMCaOiu++f/JgnGedLJH1eQWmM09p/0pvan87f91lRZS6za6nfpXyFR
oBBBKZJV9qoZ99FOJTCfA1yC+mHF9m+5vTjBuV0KffWvgZl9L+2YVubr89+z1Mkb7+0U4X2wVXLL
q6FliMENhFDTZF+IIdPkVuh1gYPQrmFp4ZS5Ik4UJU5+uoZ0VIa7xm6+NuobfjYhiAFNsoB8YG+V
sylS7TbeLUEcaWQd+gqreSZusQn5XkelES8Uz3BHgZTgo47F/XhLkx5UuKs7ECUEqsNYyKI+yBBS
2avUaiXADwku6JU8Ey8s5Wh4GArG4GcVoYcFc5fzfkyFV6l621SywIAU0DhIgPJXYZTyHVWgzaQV
DkM2y1+gTB5ste5a33SGpK2SNK2iUGwma0B8qOmLOI63bnRjlAL0x0J9/zsAKX8ee0W2ZgJAxpow
X6T6ulC23YXRu3QfkflXtmEjxe2WvFPFkgN4pPCkT4/2Dx7YkbMfTgn6QqQjSSfTXykK2aKX9cwr
B6vbBXDFQWJcf3niEzfiqvzUNHbpzWVxX8JqLv8K/awFI7q8sfVTedj2amRz/oha5k0QDTdhjlDG
5JXjHAsOdgwmx83QYFeY58MNQydjRSntq+jjmjlWCUfX5NfBeeMjeys95ZQBmro57oJVAgtima8Z
+qF9CxNQpZ+xWsj+4jQxUelCZt4KPFewo0ZY+uhQVURyDinBBIZ/DWaX1f43zYZTd4oZFS2sAeuX
LRSxaK5x3CRvVeqBos3jkKnjahRccv10q0/ZQA1lcitGEuxDHn7rEU7nxdclYYhtLHKHTQ6S6+2w
zcx3bQpUkwXXt/6KVSnQdHR8++nLqa8Pk/N5c3NgDeUyS8pAtM8mJyfcUcDC27NYMOfDVOiqJx2E
Wa+Mz/97aVW7lmi/yL2w+90ifaf4GqMG2DT5XIYnT8sXQeY2Eam4cimdkvrs1uF14aVDTZ6TyGuz
k7KVHqi1Ih9C0wB9H7dVklNgtiRbWSFZPzRepwkKtpwt+M1pxHAKCFUDwbqHD1/tK/II3tJBr09A
kv6wk4/9WmvxlFSO9PtYOiD4infuwWzMCyIAHSoBAi7tiBNcVnX65k9M2y8cmZZByrNfAv0MHmMV
yy2ig779YCXkYFFq0xpWBPpX9KaVhXUHY5MqMHJyfuugFBuPzbyIsm2H15lCaQ9k3XLAsNLer1mY
R/cq7CktScNPV6jL1sRQffCky43r04N776RZZmpoe6B+zVs1I8mhhger3EH5tjYhUnYkvXDJwalo
Fwl2+WrFjF/+7LQyXcjXGA2jZ9RBmnjZJGw5L0mIV1oYoSzGciIRh9Es9Nwg1xslJ26IRRq7Y7ht
f4hv4KWvYUQKbSfoVrNTjISx9IPfiytQBd94cQ9s8frtvp2UdDKxMMcGLhpJJfFSY0SAruspah5f
p5BUZxhUbGSCdWbZcAAbA61YpQ9z85LV2DDNe+7PjskhcPpN+5sHmMSmU50i2L/fz0gMiZ1mgOz3
AyDQodryiM8ZyjX3b6wNd07K48q6IBWt3+qWYm9wY12fTsNCTl0/26wuh/PzB3bagybIO82lDJdA
E8cPPfTnz116CVp9Aulz3q7qOR3XZ8UUKDAZe4e8nOKDbImvlGZT6/RX+tfh5OcWo4MVyVBAD0Ku
sWkMg+S0Gej5Alb0GxCDZyUgk4FbFB+NliMiN85SkdHCcZGDL9AkOTFXa5chz4sPon53gKdSPzmt
n4AXL/1aG/I7q2FNm1YU6sObC1JtBzN2H4CbwhuekJzrwgcat9Ed5lqRvh5teh133TJkR968Uimr
d5V6/9ealdqEDt2yg9IsDRwxw8+PkKUmGnH/NZYMtd26/ZfeqMB2tLPfHYbmuyRoXsK3h1EBwTeU
JeWotDvs1Kp6M+hV0/4C34DN8rQkJsOuy/zrbTgqVzZeIGMxIqxGUd34BFbgIbx1MugB32DNudZr
rU+c04d7zFSMf+DOFhy0J+Sa3ufNwlKVzFRLnn/qDwDJwg7KB206XizWPc7ybnJq98ar0jKNsWA4
PfCAtFKWCJI1me4R25TEtu44QopP2/p4PhcPqqVJj2CjItLctUy50xLCwFIDGoqasx8KMybehOAi
5zbqlHMsiZkScw/9AGCidk9OXxHZnv+DbvhH7CSn3XZ/HgbTbp6TLBi13R40Dvvp6eB4WedDCijr
w6Q/sO+BIsb+J2UdywBxH/iOor9uVMHee7tLBcA5YfsZ3U0bn6MtgxlSekuBhrq9otbuRitLXSAd
oBp3/zTwBcA5girSlBU+uFgU/lZ/XY1u9Uhh768YgN2oj/fea3zQfbf3SzXAp1NMy/yHp446eLjI
ia+OznukZGT18n55LZwn9VCMsNLBhw8Id2avbSE48yjeoUcxbST5VZdZCk/db7Ar1P9VIBkiecsd
GZAcgynjWRDWEpFbNiwrOkReHJtQ8sury+mn8DKUg18G7g0utwT+kHuUg3/E5hVrutlGsd5uWYd1
Om0Zd2hJZV8Ps7sRZoFoe5gBwv+xAJ6jdFMAc3ciKtu0R44B21kW4GIRCDNNyz/u7lj2kS8sVENN
hMduku4cWP8Bj923OJ/5hklDRvQ+wEsME2gmwwYpRt1pgiPdFdIgB7qVDoL404sq3K8DRAfQO98n
3goDa5faETMcdy4QXkxM8dVsXodOX/6goP2NNdRCeDAWQBX5l+Ljg9Hdgj9QVy1FAGhB2g63EptA
8ic0O+jai9vYSVryPDRUwtdM7KR8SCdAwJe2gOuGpzd6ucIXF57LdS0MvsZU6PQjQS0S66U/TIYn
zTBGzPW2bhvtww1p+11MmI1wrV4TlnQcmTZfE7Vb4X7RnGifmu2IWlS3ublZVJxbBkaogQa2GsB9
hyF8USaC4Sjbptu4+n/pZMUdXwcwrxoLB+76bBpWXM0hQlwXYyupYJP/F6jK8TsjuYRSPLgsPajA
2XzqNRW7SbIiPKnQoa61e355tospPEMcepMdft7iTXLlpWK0NmUgUqjnFWKEWW8FV/wCjonQ9AGI
7BpfZcSgCdRR2Nih6IWp/6QHwGMk5T8IqakDrjuFQk1QvMmCNeu88bGpqk7pBiA2YF98h+Yacd6z
OKls9TKv4QCyuB4Dof0Bn1NhOXfcc/n2iFdFQvkSR1icioJwDsirxEIMkNhqbBG1vKyxRm8zfg3k
oTREixma1D+8hqlE6rLUFGrnTyaBLDDoFwg5SjZW3GwphPMZJZl5/rG5Pu0ohCSywmy+KjtOTRWI
JJn0JYXXmpqu5yMokWF+LcjdDkOom9tjO6pIq0VetVQdhsb4Qd22Xr4SsYUDDvQ1s5Nt07H9QFin
bEN7eEdPYdVmm3YpHg/YltIzvqyNl9USZ3kYy6LycCObiVlcRZUU0FaTYfsbfmIX/yQoX8wLtwQp
XcZ/3DmJWvkUn6TSZpmRONBhQpBoy/qDQqkWeHZAovwljhGMt4BBm5DHAurMkjjemTX/d0HylWbk
gG19cvbMoXFe/EgL96lB4aVRlxqDouAJ1VvVgCGLF1FNjnT41ZpTWyIbGnYvdSlJGm8yvZE2q8QP
56iX1AXT4L2E8eN37lOCerFJK2MVaXJAB6ygTjYANDmqBXmA0uJ8t1OvpHzreFK7yAeYrsG7JckH
7pxzpaJGMw0pPaTq7OrIZrzNKzF4tij/rK/4jGs4ZqteweUF0dpkx8h+ENOm1Y+kIEtKYC+SlOvp
WND3s9DZOcj1DxCnf9xLgseTonpVn5jawGZhTq4z1cRt3aIcU9O+uI7vN7cEHNp4YLw1yMSOqSaQ
LOnDFZyJ0nqhaR4fezpmyjrBOD6GR57VBwduoeIpj091jc3cFjRk5tBbg/yZeCbU+TPucbivEnUN
blZsfMpve2iqFOvsf49CuDEi7+wrQBcj0JZUsdytcti2kOshlYuO2agPs1PSjmRPn2Jstz8SaXin
Vsftr6We7OrCzpApDzflls/avlalpCHY9VleGIFrco9xldPsMH/hHeXCbw48x9IGHDbvRXl5k9gb
SYfcMUuucNamMZf1I2fWh5lL24KC17RVKHzNSu6EK1APD59an4cXWHlGlsRoLiPkDS1V4bEnKLXj
0iw9SBK2ks3MQMcVGFJIMikdqU9k20iZVPre7m/19ZqSPLMvTeALcDR+xaW3MkwJpUDbMcWk2pIF
MSKm853b2KP6J+BLSdvmzG2Z66pZCgp7w2p+Xt5wX6XpjLDirwnFo3GbOc3ynZPuSBpSDsWgwAey
37V6oHjKZ7ZD6Fd9Lu1JSB+RaPprRYhUdVWaGnttF8gVeRtBMdm020B3irdq1+1km9TQFNGO3jjD
PUjgN4g/m1JrzGpVAqxa0fYkVthI4WYvgsigNceqCWw9eGIXcHmqqIa/sNzuT0ncuGSYTh+GTvMJ
lrta4YLULTwC925oWnPztXphUMUBgV2uyOVxtbSb95VAgRO4tm/n9LzOJ4u0FkAJKussZAJ1Iaie
rg0piftybbhmi9b9jlOzFN6Q5mMjRnojoj3c3/VpKeCNcDno12j9hMSbazof9Um4zDwbLhU7CM+2
EncTxIDw3rqd6Ojieo7sA4TFBPsgBaXg/H1fLTOhlODo0La8dlQKCjJtBdF+t2oWwAbraRtNyVrR
HfiU+AYFiPQgg8iDnMCteFlmDkpznthywkNItVEPgcTlDrqr3liwXLOgJdd1XY/arDnqvnePCuq+
FkngtBctbQHxvLSnjkrGi7Lr/VhHwKTXoL+xACWdVb9QwaPSE3RGYZW4iCylJ1RhJxFlRl5wbg2o
+iRAquBEAFNagDSdR6BbqfjvYipI+cjmZr1n3YTYfYMolbWgVVRrBRnhHhntZ5fAvwecQ0si2s6d
noEjaKQjZyfF6noxcJldOyJ5Z1whPqPcVjYBIkH07ua9B8RIgIQBxcHX4FWv+p63jy201gc9l9KH
8rWlM+aMRTOS6/FxTb4F7S7zy1iX/LT1eMjtcjeFwPcHIjYkn5X3vVF5IQLD1Ka0J8Wzjyy+E7be
2IhZxM20rYrqaKZEuNrAQ0CNe7XBB/i99vDvBChulQWZfhWPSDog1XUZlr1/CKDBG9VelvWLcqSi
ATLqalRwrygpLAmj/OlQJGF960l/oIwZhA++b1H5o9CMmmqQesZHuZGopMG5YKO9Kf7ljC6tAqNT
fJsWI171VNGAME58CVXToLjTiOVluRWgcepzHvHGMphrDq+xf6b5Hwz2njSVzohFFELg/aPaoKQ0
735H/qvb59w8QNb3MwSPVQpC6gMQOX+2VtPgr4kdulWLeKgDxzJFv0BvYyCMTK0amJ2Xy8zit13d
qKUuoIaYtNF6CaWoeWUCqM1zW9P/qq5x9H+bIhpS+icBPQVdXa8+gca2QixK++Exyl+tswxL11v3
dRS+E1REqsFEB06+Rvi+a9CmpgXQQY/mA4TWAwNqIwH1wCoxWJc5KgrN+kFoLEajx6m8WFPsiuti
q2j0/q3LFAFeWe6cAkEKVgL1Wp1o4HJI7FxPqeCz3mf09AqnweoszSsmoqXCtYfRBA6FpwrWpD/1
gZUc6IB6G0DLwG+H8VrpcJ14Zze/U81aHlAIsK3u3TmGTW8Hkz5L17jzPbJbD03+tVQMBSwOIE80
OrYRM90OD19uTW0I/wUCspgA9SYSbFxi75RYlnbKWAluPr8ZgoSF0B6KjQh598Rl0XDo4M6GNEMm
rhkYLEi25ikxMOGwEULyqftHNVPnN1hbuh738QSjbHP4JI1aoNwbRG92NGR4QzUofzlzoyv08iw3
ADa2zhtvLe1XTh2ISDKcl0vzd3zCAe4f705KiXIz86xDAPf4oEFoeuiidx5GyqT8W7J5i8iEMDbO
7suw513upoqojGyApJtHnDZgEIdEkplTNwvpFOfS6eQEqCHSR4Cmuo/0GNP6VCSeZzuBGwt9lbRZ
ZUEtD9VdB7sp96GDmeSTEDL9ISAsSrFtuI+u+UXRw38AVwpS1Tt3Pl69vsdhrRHQoXAmII/XKL/I
S6k2dgLOHUpn0pLJZ+S5nlg6QrbcX5Ov+6gez/C0gIwYC2l+VCTtV/0zK/ZSYFoVnR6gt/qQQky+
Cb/EaX3ODxSD0NZrzdVzR4J3KCotUSCk990Zb1dgBnSINTklzepJfHlIuycxh19Sx2vvAi4x7pFU
+QqUCwX10v0oIxTRfbq0iK4Fhd1ZNf0x9089+DgwLachrVcC/0gIbZqLr1eEcUKvNCLlfhlDHHMD
rtkYj0myLTY0ne6SHdAKATKf52MaqSNdiYARBZ8ePJ/7mzgCdwBtmIykt4MUKeDROaYyaxa+Hu3k
CQ2SuIIFPMkTCUjhWtFbbPMADEPX1Rf1BHqOKphpM1aDL4U/54yVKA8aRZij1U1rUne9GWe6Kfvv
6hM1c+edyL7BLRHMAOarsrgRhlYZ3oHLbIWPCLQcuPOxZZPZp3U5FWBr6Tfv9g2uoc/1vlvqIRAc
do/5Pvi/p+T9kxaedP5NE3kRes98+WU8h24sSOCYnRAWsZw4kxQCQ9pg2ib/+mhSagjWDOa2BTtM
Xf6AyjKsPf/e2OJ23loTlfWqZkU637jekk2yITU571D0xqHWfZWcUcqsGL5VwWKX+ezf/bUU4xr3
FS35PSiP724L+l5Az7zCvivIldOCOLwrC7Y7kYqyOhVLRDQAyDlBexn5ygiPc16Afiqswz9V24/m
/kfKe7qleBntxx9TCPnmLvM6NeDYTyQTkvCEKxCwGUB8OIjr4YVTt8DpibevEyYkORat61qsBjkO
y9ElwQGWHVt7Rco08+BMPMJ0q2mhimLQjU6NHJNzfer7PAT7qAHtVEc6hbVwawqQ+4WiWnITU7yM
qpHDQHcB9thFIbAPcfQJ7tyPq68in7ckqPfNS0CWsFqGqGNlLtQwnhGWIH8ACjQDjyqoaSwtAR/N
NgxQC6hSdqlfNIKwRmzuIZ0h8O7Lk2FLGWPFTK4w02KlqERkTc5ZeZds7yBNII4e0Hqfrwb3fG9B
LmnNwNhnpflxtYSTUC+EWv/4rEUUaE+22Pl2YMN2UsoOLW131hk9Gzlvf6/UrueeAL2ZpdEq7wEl
LJIj2B1ygk2Ll2jzySErqMdKTy2FnWmJlohHBzPSjfw6IzZUCoSooAaPwcN4sD6S7t6O/of7nQN5
3omLE98G3el9Dw5bApidyKlCAk+kFML72VmBxuYhIuypAGcgVYL//zgDMyuMS+pq74XyXG5pBima
BQZzlx1gDsgZc1Foet3XY+5WARtdUCa+fqRSivHD4giBz821bLq9lik5Iox3W0Bp0aoyxG9C1nkw
WUdSTjaAPDHAWL1uXGu5yByECoYY4YkQVr9if3bPqgERiBDmsoLmowPmOSwdkMtsSYsVtufuNbOb
xJBSCw7WhvdAr4oiyAR3XPx+SrJ/YzDU9aTnHfbGxWLw9AZfQMDWZWfxSnGKJPgvq5dNGArntb7O
mFUyZGWUP/E4mjtRAjkdAv5LoDgt+lz3cJTQkxRyB/yUYXHu700kEYk9THyBNSQ39mgsIMS+W18E
0Xg96gGCwG07FIwrRfp4rVfh44+r2xIRgnxAD/0YfUyjx1xSFsH9ZeGafx8YOlKMH1mk23QdeYf1
otxwa6+/yueGMIKYptFXV+qe+/R44ZinxJaYwUKz5fYBS2AkwESOaBpWX6ndvCNYaQIWiY6nApkO
go6ZU6IG8dSR46PlLym5VHssVUSehoLamJAROrEuPqHSOIgDqltXFIpuG60egBbj1sFnLJoNRHJW
9bcqY0Qfeg4gMFOTeF+PKswLQ3yvxLjDbpHpYgbdJ4cDUqfLI4qXrkoQil73vhN3Es3cJ1SZyD+R
wdD8jiEr4v9mhaF7POceU3mUKimPoKGjdySRMwmSVKm7/d9ZpSoHBZZbTwZflJxdrSmw6/IOOfg6
9GB5Fzd5qUd05K8zaCeH3CfCwapz+EsbFnSlSjcsMxUZaR8NzZ4aahRaRYHQ4zm20UL2knhbVSkR
LSKdcUf2IhuafHXzdnRq4ZWE2nmT36OdTdmyZCC1OG0wZkdtZ2fbi3f5cb5817EkOhQiv+3EBGn2
OJ+4kc6IDXE2EYcwQgTuRMm8jXSGjDy3/XImLoB+5uQTS/McKjXjps0uyHpFnQgJSWIycBBZqH3x
khpBeMVwPowe8YMvIkAseWuDxkgAP2V5d0DUcUZQReqvQWN6J4NC7jGs7T+tV6fEgh7gnV0W8xuN
w2KAWyQWCrSDIBB0n330EvbW3gDeYffrUTzA8vDktsbzrp4IcjVsdqrkMVrMdRYy9yC9qljqb8JX
eWWb3LCW/RozhIaqAz2nq93CSKLdaBB1XsO4xox1pQVOd0V8m6pfwjOdIkHpr83ZKOLnkdH6vnIy
M9uGxZRwq2pNePOPuAWXF58Lnvr+1J7kCuVvSOPZUwTrfcjllLD2jI1FH9C1P8zpReScoH7zOW+3
7GvUsd+dBFYtTKxxOg/VVagfLhb4j1zdrpAFfRwS+4Y7Dn3bYc1d7+H0/X2urCWpSpOqmXJRl22+
ios99EHiycMJPes3jQFztCzyYKhN8/BMSPPGnSLv524poH3cCuYjNOGGceCgofsHUQzbFFTJf0s3
zLhmlY4REmvAu2PQtI+JnwrnjRIcVQBJVB5JH0mHSURv5LT78DJYcNnn73MGxjRF7V4lny4oCNJ1
NpDxOFcTsLxFS/ZsbZ9J9Zl+/OJBOaybQz5BA7dYt7Cts3En+Sndedn9MOd98184wN82dQpCDp1m
L1e6OG3oz/eVB7ROhdD4oppWIFZsz6e/eiqvVFkmpS1ibKbR19Qb+3mFdBenay3sh+ZEDb0yOlp2
xrne36GdqQztLCg6425y7Al4rcSXuaanVYzzk/JyluzL9DbuGPi05OdV9FT2tiDMC0ff/brz2qlh
gWymIEn/PRlbq1KfkopqmlhtKsCRYopCybS+ldXkmYaDXVESI4FFQm1ano8bWG0wn5cCCJNfF7iG
Fm0Gj4HBR9jEZ1dD3/qxSlkYhyJy5L4lsubXsvivr1O9yQmsoxW8fCur0PLsQ4VmYPXJa4sovwjE
K2Wi1uiUYwS+fSgIJbViVhkWjcaCy5cjA4fczgoNgyKHQlrSZasIkqjosN4gPYm57ZjKp039tzH9
f92B43GlR56dgsuHn8fm2g0LDGlcxJIVFIkP9lyhMgtvnhLArKvaHdDubxZgZI/QW43vXCGcHDs2
lUbDna8omzAJVchVrexgmnbAlKkscSe1wy5OZmkK9izrwxNuqXUx/E5HXD+WdSyN56CKWttW3FuY
CRM4dmOARfag3yEnGpomMwAzBi0hSqXayokZWaASc1slEgLlJO5aE0kVHmS3lRF45+xEBhLBcatv
EboeNpoynVHAnkh68kInM+AnNafdwFcwGNYkx/LQwrirgOlHEqL/u4q1UleqRsdiRllE0dWQX6xs
LijXqQQxIBQ+Q1FfDwIsTAuE7W8ULCoGISGyOY3zRgiDcNYtiGqEZs4TWqIqDJrvnQD1qKovockk
SgwZv36NP4+NTqxvRR9bmd1VjxTTDc1cICoek0LUNT+3L4RFLLnvA+81+ggmcYdFWkYA8ajQY0IW
DUk1DXocc2xcrM0Qxz3/hbuVkvKERquAgXInLrwTdc7DpuM83NUnUD3K4FpfPEdXOq1p+fDhol4e
7s7n6vJuK/gK83R+eomDvGvTviMVWuP75VjqUiOxY2aw/NytS0DfaeN/7UOrGIiEq2Pow9bKMp73
vT1+qUdlnLA4FeVgen7yjAZ6wnjsz378U1udvcxqPHBE8CMoTp+H4XKQscAyAGn6Hxo1+Al20tit
/z20b3pNdRFmJYCzcX3o7uaRnp1W7cpzaH0bZOO3AMYzQ7EPx21kmiVdxOSIW7u59GbYFfcEo+a+
M5gtOEh533ALNyj+oDCcVEcSVzvr1/tnlKb5l1qZ8dwnLSudZIJSNpNjkRfw2bL9BgtNiYbmRL1O
ZFh7qCBVTgaWr44m6lg1d4daxOGpznlsNnriIn3jBkF/8TmkwjGJcwRQT2CvfU2YqqIEaxseTilS
+alJ1xHq1+i39C6se1BgHjl+/mYeyxPMsKiXWVocQiFxv5hqflTFE4S6Erodzm0VGjhMAZo0IZ52
ENyugvtwkP042XNDh3hvOjjg1lVAJRVe0Rmtm6KyvG4xfq4PobTEcnR+EWsjwR53jvTET+KekzH4
W+BrLtuDXpxxmUP5Xgry96fRbCGdysLGrC08O2tB3mTPS2NBnHgp6awwisKmxbuIzedQGSFmWmKi
LGRZx8R5+4HXd8DjOR0OcFz7v3mDNBlovSfFnBNUX43H+gPXdpyyB0x9BIyb71MGeurMIe2WCuF2
KDuO12Cbgcrd9suls9JyxaVz87k6u/qOntXKEWfLpKVHwICqtDcdOhh2uNdI1pv29n1sLDpk+q0L
aruULPurrhUEZjhdVCOnejW1lOD1ow/tE15tTMXuPS9W1AoWuADaUouO/pYnZ785p77IFLG8rOzW
Th2qz4+n9SVQ0W/tU1357kqILp7ySmMK3iOPWCsib2nPkRvchb1kRJxjvZo2hLIJkNjoQtS8ByM5
t/pckxRax2rDj2nrRvrPDJ/1FwzlixO9YiRf05OVIvviHVPub1HlXI3xG8g3ce7kRKeQW23VMDlT
6XoR5CCT0qNuGS9q2c4x6brOQ8wzq0/ubwLJDhh+FuNbqPaoTxmE4hK0BvslbrpgRPqJzXxbOv9s
cpH9JwzPDbnaIRwrcpYOhHfe50yKBjvM9HAV3CzCdeiyc5FcrDBsqMhTP9YecMjNpL/GmOIuOmJ+
L/ldGhj5PoVE/0Y9TYSpJx4wNXpMwqNbAzXyJx2meFi/kz439Bz6YyM/RaCn1HqFi7mhU0eV0j4P
GnEnVwovQAeIN90LF9iR/dEIiel3P5oCmZc/U6R7juBj1fHn2zarG0Tr9sJPUdk+KJbqyUWg0Fim
Y22wep6TEH/B1ibPeH6pSiR0R7C7B23SI/zN3aJm/ZHzMLr/S3i4HiKwtLJiuAaem1eTbejmMMcV
THz1mVwxosh4uxtR/VQXIZkEfMiMON4wDfXUjdBka3Yx/hbMhc17hTo4fsqBJ4pmMl+ImTd/ciM6
Q6UoDQQ+sbmbTlCSCVU2cZK+wAWaWPq/6ENHVgbR1gtYDda/nedBsOUkptZmo9kcO7GV2rbk3Xrx
VaGXO/EQErEIY83ARoQ94lanWDe+fg2tCtaD3O5hS/4TpAN7sVGfeSMOUyioiqBAPOa4BQ2n8z9q
2K2lV/z7+XFtNGIkseIoAKwka1iPOaAW9oBKptE9+e5zyxTjYPUGWAppBx3aRAfFCh5BymTNy1np
+iqOrzXpPR2RsihCmXdIXYtCgXj7NhBo4go6hGFnZToyTtSZ46ZcekRCQGgjKeJjwT5Sp9NFgs6q
BbtQ/JuY07S/jSxXtsIhDk3IfWsiGRQ02BtwH8URXBu2h5KPl6zX5dw9VDuTGtlMLzTyWRzJxYPG
Q52dNIjIl8LY+fB4sJV+hsudVm+yK42xssOPY9FWUypderYE3NIzQ1K40Oi/gTLG9u2qAQNxPE8r
jzXM7S7V0mHDPL0L+8z8jCrznMSPRJBRk0oVQG3yzwXWz5/eEOsljfz02jxfxj2aQu1zPJffKMpG
jCGRQN+HXAkVuVKvb3oVPOBnQ/cSB67keFENcZ0dcFib8WTl2jtth0BpzkKMgz4WyFWCYDmSm3mF
vR+L5GUlHncNeBA3wsdZcBNGdS5dKAzLYX73sAIrLjiEW/w4oTK5QuZRluyQn+At4cKXnnpahzMr
v3kN3IKXYCF08Jr06qXcA55uSHs+uhDm2AQHMre8xQz4oI/SQ53l2y0m1YpQWNKFB9ux63ixBFTN
G45ymHHTaFXKldMcnyzWMw8IJpy27VA7dEqKB42oGQ8DrZQtVodRbXC5DL19AGSxSfThVn9h61sy
57dVIi8Xjz2HE6QbeFOrAzAgN7HmM96DRaEsHusZb8v/si0sQ6GmcqLGRn3EzuZZ7yCkm9jg/VsW
Gw5WSrO2d8B2WvltdSWJlb2Ig9svDT+bmZ678Be5hWmKgotYmgFsShesJECHb22ib8BpWEEI9Nh0
MiPxF6+Zi613i5L6zHnKt0TTGYhFQ3Lx+WfmUHZB/HW87E0n66YxCJijX8K9jpi6REBpIk1UlEI5
qquvENTBJ5/qyguqLEovd64GQG5cXYvGZFpzqeDco12GC96xWgFh26vnrslp/Uk3Z1LHJXka/Edk
dDMY6FgI+NeQP2v+2qwQ8UrUZewnp/mO2l+Fa0jjQpqnOqJ74Brg43Foc4V9AsoRY0H+ALwMwhLD
DfBTYw1rWzdpeBbI14xIV7hj7kSb3hSQd1+XFhBWzxszYrwfvwCBapnZ1xmQVKaAgxApd+DlvI8a
KnZUL+Gp1IWl7jaSjb3+VpZEJCBAtcKpN8UW72rqK618Nw4iRkBZnefzdTW56cNXGBpm0+1sL2Ga
6/Yp2cK8jx/kzkYLV+q021cw7reFqa5OmCGsoiOvkOsPkUOYKgFfskL0NycrHhNQ2WHEZc7eEVvY
Y1T8E0TmVG13sfn7Si8PoSk0yrTFwSZha4NRy757zl/haMqylnnijajkQ5L/4LF7Vzf0hhRe6IDU
hWuzu5/oQK4/SOa+W2OLDXPulkd84k/6B3Bjc3M3jBSSVjSLHDxxWODCtHoIWoWNwmezaoECOUXj
liFWi5690JJ7JA2B/8wZd5vrQ7yBHA37bYoi2gbiVgRzwLe1hB//qQWiVYQ1+Wm91GC3sEbnFMjN
TGXc6m4b/CWTwH6yfNE1JNiKQ4E4C5aDc84BTkBsOlOkW5/zXRK98Pciv4pPt7pdIM2pNI4pA90J
VfFwrNd2zVUD6oyaK/T1MDj4Kc4M1S13jDjr/PTxVJUwBOOis35kuwknDIifFOtYw31mmqjKZj08
bibjPpmu0FMy+oILQljii7I95nopwGuLVFk8bMaHJiGWFZxCWShpN2rOLwcLqERBp2TwO668VDSC
BwXOtrRMy+qtOfB/dZPq6umROLnU3LjaWmzwqbu4RmmadGboo/SGCwxrVjlxUcv241ZOAqazvSAD
+Ie0ihm/dpg7W9n5Z+rbUUM2mf/A7HZvQqSaIha7lz+am+tbOK6EOCxDdHK4vf2C1/lvQkvhFuMi
yn2WpuAfKLqxMryQKFabgLmKz1J026d1tmHVHaAe5K28JKKD5dqXrnaLh70//9ese1zmlz6OooJW
SxXqk/EhlppDMTjuRH2HbNWPRlYsrrjYRsMVFLvWoD7QuEpn2UWeeUDkHxg5ZR2A47pS20d9aOCE
5EMvhpfxcftHw2BXQ8axoW/ivI/QyY9uE8EQ/I1ANhFK1wsTHYcniCYu8yh2wWcTTNJqGoU/BHuq
6+CFoSSDw7JZMCY1ZW2sdTrSwNiRwrkagZNPN0KpKDiwBxpiNA7hSd41WDgaWCYG3V4tGfDsZYds
TpXj6uQFWcwbN9aDF9Op9yI83kp3lGpK86B7C7ewEEcXCsTudKNDCtlXjGwh7ijaYBmLrey3juG5
PKxm1JtXE8Wm/WsJ3pRoXQQqc1FUKn17PhkOoE1zVpHoiUFOMukXvBQTbDZCVNdQypSqtOn1O+pL
oR8WfiNGXUC4y1PmX0Sg0XP5X3Ni9qSb2Md3bhRNWJJG7J7Qc7Jri4fc7NSnR4G8vmwkvVroZzjF
2sJNrPkKuM4SJZp+sqj5axOmYPmTLhGvYIuzPX6B5ERZNOFxhGffLeX7Hd/1cpZxK8/Ww/vFhkmP
Pf6f9vy/FADUMWzB7nmz6y5p8vv3AYajM2KfY0Y8HJDOFl8mTxzpYBW4HtZo7jeUYWViBhrLUVXP
+IT9IoMfdJlGJqdqtdp5DorhuJbUiOYohra7H70b0z007RTB1F3lFBzGhcujEBhqmem3GfsECKUL
p9xPswZeSAKBq+E3ed860ep/SNq0usGorFJUM0viMBYciJ9A+1iH8v/aV0+RwQZipw1xbJ8DXDqm
u6vEm0aD7lhiQIm+jTuYdOn4XMjLoUDnVvcc2v0c80Kxza2ZBVD6E9mohMPON2jVBfsY8b6GYXAK
h2K+/X4UDrJg38tqTS4CGrISnhncUEbs671peEXPWJbzNybYN3uKyR6JHGzrPZ6d3H53O0v9hsxi
fjP3OJK6OhWmxrNlyurL6TC7ElytpidIIPUj511MIRhFK5BSnli6bQnhuWDgd2D4bdYGESd0C4xP
6JUt+PLqvyM1Gxh5Gxn2CPQ53wICdx8bFUZ21bdHAZlogufblb63rzPgLvuhOJA4RdzHauDbFhri
ml+hAzCSzT+l1mT7Sgd3QaEmriDY9QO//kWd6mUPOyjjkYXmZQwXzkW0a97vydYh3MQAIzChdETX
5nmAgRm0/WZjcHwMstnyKZAlAaNaSLXMi7mtbOmftuyUICdkJJAVLvBupOI74lFYLsdSCHzeBxGY
k1s/pnwa/1BKN8PNfrb0Oa6T9qBxhw+A+TYNgH0LJOinPIiLrwCuMN7bhvXz24BYytH2RHQ04rsa
nPumDVJTyznygcNbVmbt5GPfEaa3d68PSx6Szye+vcq3xOFczugdCVYprPdhxq1iDNfa25UCAuct
hGiXjtTDqDfuYnC8et59kpM6155POn0TPr4/2bwfK9/NttZ78IgRABo25bxfL0wfsWFEW4IxLk6v
YqzB+v5eh2QgBVQikLGkupwxrzXuXsR5kfIgMFbst4caXgxavoGEpuFtts1coSZ50d9QVS5dPD9s
wZ1PpYh1k29yNKwlR5Uap3JtFraMnnnLmWOCxchQWGFwQfX3wu06xApjoT5+G9cl1gPjNqaOiIWY
QTiisp8mp2VKeiiidZiQB3ThHDabLZWtanQS4j15RsF8qJhFBi4a39mvQgHXOf9h0RdwQZ/Sg2bo
EM46zPYJ0VoXtke3ohC0TszqjN6iS/WTC45m2g6AL4APoFoMgWANhxaSSgN0cA8UvvOB5NuQXM1k
PVi8cjw8torz+MRx+wlnnAA0O5Lodkd5Prhi6L5sE6dqnhVL8zUNHHRsAsvZoPJc8MYQIis0aLqM
lCHw3x3nfp5WrvhfIAdImrGip34E0ItewPZUHl2cIt6OlGils2Jfed/dka+AibTJexZ1S5pWimYn
uQ8ephNeWHOsVStC6ryLSubWrGNmEuDjNuRJKN1LpEWGqSTE7NYcpw5yccdJmPe4lRU3RVcFs36C
s7KtDQvakA3C50A76TF4yl7uC9jAgYPwRx4LN1Ar2qujrp05II1EVzwxlHXPL1+NM4WyspnNTUYD
BmlMibdIBUE02CP8iyxNlGNbGaoHaJirVwwQsxhAkBEK2fAzuLq3H0RH5CsG8iUsTMS8jS2WTTI9
WrmEivTUrX37Xs7FSnIqJ/7k8/8eaHOT85+rMMsB/bYg3pPbBbiIkMS2I9xs6hMwQNM/nkZtsANb
AWSfdTriC0LJYCpwx1jly2WvqRX9DijxYeA8H2jsZBpLvCWMHqoRk7WdfHvcVcSMpXHBpmiIZ8PH
eCMyAoROv+1wH5AhPLyKfbxygZWPYeaETCPMdZEIgjHRWypJua7DC45BGBSjDmlE7c5Uh/iMRjLD
IQ5WNgDlwzE+Nc6U4cdMIGRTC681u/GJkUmqmJMy/A37G3t9TC9LG7otX4AhwHMkc77M0h5Z0L5q
olN0/At48bi9clUMiYPUi89U1aoOmhaQoeuwp5+Kh8s6t3XO25AtaxHKfRGCF1WC4z9TR2DZBA6L
DRRWoOiRBht2oewqXiQlaRU9Ir7DsEygipOu6tMlPbVk9HBjHGPMcPwyi/TVF08XCKaQErc4PVup
9acy2YQbdfW2IBIrwMLKyRNOgDbbCMNnCpqdDEfWR4wLXYqENeVsDgYXiSX5uLHihCGFlgPMddGY
sY6uO1u3gz81raSFhojagWp9+HIRuLNcDb2GfyHXcExC80aRJG5Wjwh1EerN1K0/QfQxXCRAShg4
TGm7soIpZakpWC/t02kMNlr48IVXhTgAJGkC1I7qxUEGnXsTujNYtVCZfFiJjuFJY1ca6+7MtoYN
FbmULSEEwe/rbK0n1oEf+8JhQT6eMmPP5S/2EChMspMfCDHQvrn0JY9uNdSPw8Vxt27yKijY8RQ9
38+SHKKrRDZx+9pN/iE2g+2jeq9qB83rfIKByWFpmHqrmHsOcl3LmfFJbnqrEh2OubD1tIz5Pzxm
BB+QasE3HNrZMTeOG16N955cxtV0XS69g/i3XluvpHRS/Iwg4vP5igNdy6qKWUWbELiX6ocdj2ZL
TVSQnvWdrWCKsXWs0NLrg947r0l21yxDhnAQxkq1ycWjYqKs+0OxPo0JwKGiGEePoyaoFo1MW6d0
Ha+pZ3T80FJmGODLt+11NDU4ryPKhXKc09mzcOIQ2QQyTa/9X/ivR5bpPBu11QP6wGk3TI4gtyGv
meiejBl8i6QlSnoI4VozNejmxlc+d1jWV4p1Rr0NLhYY7ONlDukVijcnfdMrT9LpWYtxOSwvWnP7
rFXBmuOKwkuhzdmLtRDNeAT7prg1RPlagR39crSuofcNTiGl4exbi63gOZDaZNEJD62ZgQHXZKMH
i+XKAerTz0TDZvjJuHW7LQFsds51UsbUBBuYSKhomd9kVB3JWL6zWXThbvcI2EAFtIFPQ1vQWofM
M9kY5h6BIXCG9J+dyiPGWb6NuLliVHbQ9Bza+pIOuVEc3JJy4CvGx17B+FxNIfHyq6bKJuyNUAn8
ZEEjmL4YETMOU2iCblibjcxP7mCNn58a2gapfqOBPsCGaSwDGAEZIRfHKjfhyliDzARxaLX2bVMs
FP0Ko2aOtccz+I4meBqqsxMzivlA7oTOhflof20RV6HAF7kGcJyhmazQFqBXKTJipvrOqjG3vuIQ
euxbGVAYB7FF4c3tiGejugKSDHHPfJyBlRgZNyaTSPkLYNOSmwIeDYotBnsIltOl3rwwoumgOoKT
9ye7ruUzRyp7xbQVjJbKPGUkVkbBuPU03iiSO8+t31qAl63crSRjm81Vfo3qwUxRIi0Xwx0xwSrm
EcZ6/M7thS7ufd+i8rhVncYDooHR1EPJiQXG966+jugMC7h8GrbnC3EQrjxaV32Qf2PxGDuKzYOi
XphxdftaRTVjpN3mf2/A5BLXFcIDmjJPb75yPiEMn6N0EGBW2I7u5t/R5rFcFVq9XVZKyjgZEGIj
V35tlLJniOiw6jgjd2NV+BYp7/wm9KEo2ryYUxstsCk1Jdh9o99LU5keAJOswSyUAEQhm15TkTVv
fP1Xe72SLhfPyBYJr7oBDn5CIZ6VQg1MPpcvmpBjxunOzyTGlllmkxpr8kZrksVXET/6iX/z7dso
p3oEzCbAM6vi4jmLbmL7+xn/jMZST37JvgLNZ1r7/AvemEzbr3zFgDniPI9jrgSji388/16bR/Vi
FaWsUVQIXaIbDTF9M6X8UiF91DoH1Agd9Qn3OMvzd0watjydl85mwjDuPgt8BSz2ephiKejtjs9k
iX6BtLHRThHKnl2I9TXd8RLdzOK0de2f13EfWg1v9Imi+blHdBGQxvvAjMp65MFy7GH8/wLQOaFI
Opj5f/3/dP54/b0plnliE09xjSUimSBrcDqj4e0qUAOTH2LZtmU4banNg8iUXJj/5+ZL/N1VhCWn
5g4Y1WJ0NvOTUcbUx2GOUag5luacgyFacTA9dnqg1OCevAjejFyRC6c1HEbD96G137eo+DIAmT3V
fX540duYNJZ2zYQuoUWVc7KuYapPNQPw/AoaG0yleIUTXYXExU8EFq8/GrQQ3BNP+j/wDrPeyVqV
M96fohWCWHCRWzPFNKaqBJEXEqK1WBCn8n/hornzSLVd/Oott7M2IuPQ+nBzmZ/Mrqk2YW6qeNpW
UDOUpWBbkffxxQfjYbL7outWJ/WRaALMzs63XzC5BEelxR2mWnUh8iWMdCLo6Iciw/Hqmzo8iIGV
KUxBOktS5jsNrnwdaup9Kl4rjR4Buer0nY7seL+XkZ7WzOYDt+rZDa7nE+9hRH2HWKxRcNkHfIhK
4Xw9aLEFVr1c2yS8ul8EYJ0ep61vpfcUXpe7wiUac2XG+DuNT82R7u8GYxSIxmZIGNfgNcdtDCs8
1YSuQhhrUmA7ocgt+4jxACscx3bIDLnTcZYs3c2DULNA04RP64LMz+VDKFMpk7t5wa+l1J0rmgLy
vQ24bOGakLhIuro+FG1FjGQhUlYVnz0RgIZmlZBVXg4cS5iDM6lXuikaTMlH0MhFMl8hzZZ3c5eb
ykn8I2QJgeddtv+D1NJ7fxz4U2ZDR3yKA9yf7NsAkhFl0ISgqQLjSgF95tDby7aMKGYI7CzLMLi2
oxQn8WBNOAd90xTWeeJOeMxMYLoXPl6+dPZgBVgtW4mGY9dpPQ/ERHfWdeappgfhPTwlDsP6N/At
fxB1iNWsqm/747V5yyRi84HGLOWRkTjerGQ84sC31dmyePJgZWxwfGXlp0uVoazjQwTeTjwvzT8T
/mWaM+oV0fQ9dedzNloNb6wiRwdtteCI3E6n3j4X9IRbEHScGQEvRhZu0BgglLaO68OJ1nov9Otr
INtCVEyDa1B9c96gcmvJ68KB2GPr1Y/1TcV1zBpaDJsI799uCaO7KB666YjB5zXeg1AGc3YJgltT
VyJz11tmB9Nw9CmaZL+Qx+x9hPwnFkVEZfaKQb0xoGnlceNQAm66u4noLTX3eEVfPoGnrMOxWdhL
zxZVkyRilJyMxIuqWvB1BJaHY46WC8K2QVBd9uvhG5zkSsFsrYTgcr/R72FkYK+W2RKkSxxy2qRR
SoA7rGKjGRofqhhzgyDnmDDuq5v+feAVGoVvs2iELicvM1Xhw4CTUreWJ30Y6zXiefL9EybR/dAe
wiMnLCRagoIibchm0l12h1xXusUrsDvYmSXAvQHqj1XhI8jrKt2YEklfH8+Is7I2I2VV5Tnse1GU
dSptDMSrqtWJAdTEc6+DmjEngNjtwwRAC2rTl0NiPlVU9h13pYbpn4iDm2nbyDIsMvffm68mkMbM
FNjQKH1ijV1GyDYB6o4lpW9pVD2J2WV42jcq10aUXXDOJ9vmaCqH8SqtSSvtwGGSjFaQcW9dKvzZ
rZqaF6gFSM7vOfyD7RRSjctfbPtKSySxw98Y5y4gB1Sy0LQkBSg8kXEGwYUn7DTibjpUmlpbSZaj
MXE/eH/KsighH9Gf+S82xA8o4vgQ7xSVSFFbPfESVuWKw90Mg/Ese7bJ50O1dzKVICRpTeS20OS2
Zc8mX3VZJjqzE/jHgIqnpuc1bFedT2czDyY/AtYav4165tlzPc74BSTNZ35FJ59koqC8IU/OX9IV
o/t6Kh55FhgTF8r+40YccuBAXCHWIeARHeXjFIFrp8IphchIOuvW3/qLs/0o0AZwsDtaVIs2mcXO
kcet3KntSsAnTYUspD9bB2U0XtJgl9/eqc59BqSmbpaFRXkopyF+6pOE6L7gnVCmpOJpTPMq0LI7
AxZLKWb5IHIBFzRoDEFoncPdCoWWoQR2hpRCjXk5qTLADhGKJkoptLSngJW40ib4j9SopYjKWluH
ChlDWFefdaR3E4v8D8R7pADPNhIKZ/+30MzDkCk0bbVlI+d3iqH9WY5Pfjbk+YSVo1+kawOdwr8s
R+bWBIaj9vEXeCQIANik5ATvOdPqAg5RMppICvMTaUPhu3c9N8JLRmzkQhCGKh1zD0cjh1ZaHAzs
Aq+OnjTu8e7GM2HVMK073owLpYSBnQ60iPnbC8EKlHmgx3gHJCQqg1puhq+vavkkrlW7SQdFX+TQ
Prsd2uoIIYM3gGQhMeyX99Z5zYbyjF34W7R349pjGkNLEDCAvQwEsLdvj8CIVjbdW+93OpaBeLWf
YrEqZfbAacaxgVcs5Uopmf+nkpxTJ8G6iOUEqkYPxZQfTJgmtFdve8kQYQpUTTUHZayaqF54iu/O
LyhplONzCYuIeo2Ts2mZEaEKatAV09BX+nIxnGPO5462k6hwGGIH9310ITqihiuWMxNgFarwbzMO
JadS1Ks8rnoariewbdrykZZEt2DQKwusSJnk7+lZ85pSuln9a9JaGcKvmgZGiJQyf+PqJ96WNer3
PlKewiCE2Nbqd2+iOoVdfGmwr/m/vgXjsafjbiORjRrQvX9z09OTba7gCsFAZhNqOHwsYa7hopnj
RV/+ebVM1bmfi0Iq/VjJwsc+pSMm0AqbWY3tbRrLsPJs1flm+/kDMXjgeGuzVmlGXVSSzvTIl7TX
+OUhFEMHETcOW+jQw+wBUVrs31NWkNl6VHA0Xty7mF3mwtCQMolLP0i0uGoMqvYvBMZKObqcigrQ
LBlucX6pEP1Zgm6heKioJwAo3+tq8+8eDcix3X9H3EOdPaxu7QGttJDgNfMdXZZHV9IzxpT7ghuy
mONeaLWmV2KEg3MAZs3UgWwTut27vj639bz266RtHvThX2B9pPanuNpOw+w8ThSOYUpffMwsRhKf
U9i8/pjTyM7VRfXcfEzpwEZSkS8mk3so/FE6HZzaaSc0P00AI/oU5FJrY8p1jlFv/wifPWyIIxUk
S+MfhxR6LSwsQJhFP/eF5bLoFmZrWIubuoXSXcDzKbxQLbShGmlGz4hdIlHOIfQ08MCOaf0mJqck
iIgXB9jk2cMU76PJgye+dcwaoLyQaZ3SSa7kPRZSpY/6repbLoxyxDbCSvUw+5+rzqrm2VJTyID7
tqMRZCOPeqYgnBo5/8q6d+q4+9uu4CD/fJHIZaauv8IX4WeyZYpQUH/31hsCStw6Fjn5Zq7easIn
S2ssVDPDwSgGoEFNHoEyAaIagOdHKghKvMHvzMeI+Hkxwu1rv7hGzy8ex7lej2J1CPJvw3wCJ6jU
BFbq5TACh5HWMWUoHpUIGajzF3ywnonIzHP8+4CcJkdVM4f2y29t5X65t9x6dXfWcZDT09p59wvP
UOf5fM/2SBXr5JWo5VBBT8/RZXKw/ALs1ZQ14ZpEfzzE8OvlSxIljfu2qIu53KuF9nx01DT1Gc+c
+QvFNMkGudi/BpNf6LKacFXc8wiGWajUH4Obmn++f+NIm1uEZtn5ddmAeNJXDH4neOJmr4XA96J7
lHSnVnvYgE/p9OeZ57W5or7R9LSPoHXOTaF4oT4YVY56+wUOXkMEoVM+k85blp/OCPtcg0n1lAYr
q8dWUwkXJvhP5t7ckC39PHEzWUg7Iiel1Sea+XF4umS9BSpn9nEaMbGa4Ed+KY4fqNriuXYIN05y
D8HtQP22eaGPL4u4EZvdhLXqT0b1hH2D+eNJ6Dkh/Bgfpo0VkowlZrk5dF5V4rfO7XHd8rU4M1qx
Xqwu9dFJ7wkeFCmxRkT/mnKiGAd/S4KD0U01t+IqLK+jkJKutpkYRzhgzFZoEb5xykIDnpgJ6XAR
zqlS9a2VoLw7VvOpCjFB8W3275R4Eo+gJUJsef3nkQMc68NYnmiM8A2x5WtVFtYLlNMU2Yl8VxhY
dQ8QtesXI/4fnHjJE1v7QfyIAjRUnZ5eU/WhteAa4IDkGq1LX+exAiZ8uiezP581SVEXZAcyKtYM
qpecDh999Uc0TdQnRaLFxKotf/sh1QXTdfrAYBfeOe6vvTclgSUjTygU+WS8/CzSpZJvBTjer7rD
P/+qtxncaCFRnsqgZW8NFFtOnAW9uZNpDb939SC4JOwhpLwYhqq6c6qdZfbjhFioA7mEFD8HiptT
PoVi03aJgx58e3u6e/DY+lv1E/4hHgSFdz5FGGBET8ECgMOzrNdOsZ6zZKf1d6byqGejM5PwUZ2b
eDF8r4pAGtDTn1Hy4TQRfyTMd+pU2kiVE/OKfh9ZbsBCEGliPFVBcoOKoKL3SzIYZbBP99/97DNX
9SpUtyp4HnSVAGeMyTxg83pHciFFs3PzTct2ng1Dv4pekLkui8aRZJ6203nJQ5EUx1aWUONnNNWB
9EqQmqrRM5SpVwLZSbw/yDmUWbnHShH5uzm94ywHl+nGoAB1+5v6exwslG4JGYbOwMxlxwXzYXbD
YXa2MJU6BLqwDrmC2jv4FysMzQpsT/RwtptQBCF2D5RliznX0lAetjUg08yXBK0OpT7TuNz1NTbP
ePgkPjI6i0CG0uXr0B8PfW6lyi4IwY/5c4AkYRFgMpExGTAvrj0Bubgpv29lnfw3YlePvL/OyctS
jLv1dD7pPDmSgUEL40zPcOaUfY5ueIqWEgaFdGcZqA0j9jdVyOLa5qxofQrFSv72GWyGSzPBVXnP
4dV5Ws9Y9cwSuJ634Ub/o8pA7W92oBhFsYe1kpaOTG/7RChYTi+Ofotufs1O1UFHVgDGH4ocj3HE
7AYv8+lsP/FxJjU9EYgeD2M/Mysj9msOopBjLXIiuITPVqxMPR/3Mg3IXssNJp7cXYTbJ7qD1flY
/kevC2+COCX/Tk8dStBUHzhi5ukAyR5FEGRUrgQ1qdW3FBQoxwZkujqAAYiKlmtjCqc8SJUP8LUK
e5xfKG8TBS+e73LaJ2QxpDQJnvlpD7kg8BV8xuhHbDmxLPL9LYbcH4ll7cNsPwrIdvet56uA+b0m
16PFRed5mKgcri1D4ebdE6jZCiU1uLubpVRsUhbbgo9jFhLT9Wb6jrM/KhhWDmNw4QXZAvizbbHo
YveBWc/uWitDAGn1ocDB/4TEaCKp+l4zTMFO+r1Ex7YCNBJsIY2ovu7QxZg30uo4B9Vmu5fxIvQ5
cYqiubqoo88/Gdo2sFaHm2QY0r8IeoKA0tFt4w6PQrOVOR8StZkYoXiF/E1ghxmmcgjl0Y174fhG
0R8SX1LpOkKMJT+lhIdhzpEQxiulvyNa78gO4t/HYEJUoiVFlloAcJqxAyktpLirNcH9GnxYrqY/
RHVtwmekNX54Yt9CJ+2IkmvwIK9THBHDp81q7tYpTXk2MzTD7thE3JTucK1kSVG4pz6C6utPk5Jg
2UOoGRlvzyOVvw4DFslqtdWOmHHxu6/24GFYQbQPvKRy4vZRBygVWnjKUwsn81CbtbZEk6bQLorH
7985sLD55OdEaHlXAByfBK+zNzf6DzQFe9FCHfA5VhDho8DHXGP+TEoN+6RTQSgLKP6FNf6oqvgH
TCbb1mEITmu6aUZ61W2ftWpuyblL4WHmPEXqUpldzItXmEkxDjaECLNVZ0YKEqpuuoeRY+/dm/ND
tBt5b6ljCXuPPHKyMXccCZEdcW64nDTdzP32wuFCwEUbwBrlhqgHWtxdxBssxneIgR7PK92SSQxM
6XoHQ+g29j4Vsq59pEzYulnotT8IuI2XBJHSmFO27IT/VMk/9flyw4MCzFqBug1uP/U1f4+wDcbS
yH1GU/gnOGXE5WYvOC9tYm8hkLedwOxGRRvhREW+ayPr04xIjH19xjjf+ns8coA3fg7gEOajdDLe
PkE/4+lfsZ11K16UmNg4TyxRdJGvwe3HeYCLKDrZsLG3zGflNopU6+ZPPPV78fViJD/Vxa4ry2Kw
/vG8jgeNu/znfVpOUIn/zSvlmYh2EmcmA4JSz3YanD2epiYdau+4kmmZ51FzPj6zQb2QJywqSz8C
UHWdqdwxMR45sYIQ/cw5Vzd58a44O8XrpglSRszXExWFxrvrWD7pL45BEqW/bRceNU6FuXIygKsU
m6udppJKkGcheYMRINL6yYQ+B5fxsDQkDJcCABeOWwTFMeOM4Qh8QSlAM2CwnY/3+wh/gGot4+7R
f4RBsu+id1/T51xuncijxc9UzEl8q4eRbnuoEx/fF+FquhrBDxSVV+asTVOExmeyhtscQPzzfvzu
H2YB4lPNWOeBd9xPzq/mKCWauZrDQFxMdyzF4RQcCo8USVpJ9HlNht/eILs/GyfmiqsT9fMDowc8
ft5bYkGUUd5RPghSTe4cpPUrdgG0qHb8LhAO70DzLbmK6Cmo+JBd5GVfkSfg7ctzNQzqLaRvsCqT
5k1/aPnkeyQfUzwFYdgV994PImWyKbH2WrrA4eByKwMMTkgm6/65JNylprxWyntFNads4V27AI38
IWv1IQA1WCstOTjcLrbDSUcD2txEVXxa7mYZvSsg5ONKjnY+eIjAiv7Ie2qVRW3ahsT8DvT5JQQ4
3JiGI4djGx7llyuKuNqnNaXHo1TMetf2OM6ZPBRruHE3nJcALtYd4Ck7LF64fzs4+bgvJiNGk1ry
0UBNU6/DRroGM0jRimvu6ekOdQElvqHi5o7/OCOwZx7VD8GhxIFYYcuvv2jymOC80LYIeoKWBY6n
P+Z45wKXQBBtE3rmBYMBXUWe68zHi3QC+E0a4sw/f6PakTcPK9Cuc09GVJczYYjjNRW4oxJHKWRW
DFWEupizFz3VrkHvEA9Ba6t6ayQxWTaoMqtyyTLi4LfamTa0/2812Q6mQh9UsBxD6J7DajdUs0uL
VToJBoLl1S8zzhk8NdUbodE/WrmKeRQn51wlPMCGTgSTtzgsJ5Zy4QM9GS6bumcDTQJ32eMnIaIh
wAhqhsSlWMgNXP4iM8Ser1Ave4aCNInkjBOVKRG6ETj48bG0wAGab8z1Kh3+L28dKeM+bhxdW2yJ
aHumkAGU8k+pq6AfTTooz+iCAPmjSUi7u1SnfF3ZKDJdOTTvdaZBIp8Tm1Fua7mcJLlnP8YOPC1I
3EIi1LPrSi5h88T0u63lNvlkk/1Bm9jWAvGjM871Oukm/DbknqGiUM9UmJqToEJ8Ezjsv9U1w8L6
E8FE4evTTV5eiouOjPIfQ5CvqVR7quyewpq1Z3K2Hc8WislsUqRqaT/1mSMduBXiWqEbOXlLLYuy
byb6lvWs90pI5vA9SPVISNuQ4IRDV+G5DUmlQZgPZbEwsJp2n4JxDxpcOYqK8fvGYC79m1NQ0eNO
ID7yZeO3w1sZuICsTZlgr3SvgngtHY3bRKET4nB7a1HpDewDticncO1zAk6kfBigwBZHEOE3lRix
FEFOxZX1TzNjWjStmJ6uhMegMJcuQwk3FVpuaGLErTblHEGQSvIncXL8VdehSGNmdUhhL5/h3Lwk
oGsAVj+/T8k3vN5eX+I9zDM10mIujFLM7ECxSjlgstgFq5QvX7skjZcnHW29qXKK699EtfBeQHuj
wbiON6hA0ONQTTtWf2FSK381g29YJqoe3R9MEgXog7Ps/K7myOWfGb6vrpb2Wn2PGxgAtXdPz+/9
WeSPqdl8lj7vO28h28JIVU+qI/+dvdxpdDrLsoj4TXSIPFlJHScNlq9x22MZziOEsvnaFJQb83PQ
0lCOwrFJCVKoUWWBaSpljwwM5oktqpDyqtsS9bcv5PU4n+qa/wEoHs7FCNd2KqQWNwfR/qoTCEdh
HIpNXOgRFc5PB6XB3AV3vXJ4ZXX0ZMkt7YGTaCcvJxKhPq0HPDc+rCkLv+3YTqooSTAC40SamXKn
QAl7eLcq/QPQkgbfRbOTeDf4ZrL+qgS+6lEbTLcY8psS9AxW/cMQNiq9QLDpnERgtgYag7zN29rf
eVTUxpBR7UgiOFqaku78yDGcocdwTnsx1za9V6qYqNdsTh5ioQ2BgT84/7GYmXRcLjKQm+2Nk3NH
rzi9BDr8H8HuLZ3q+hFLDnP2EPLZ9m1SkxUhWHro1h4IDR6dSMdeAKDduqmYQIk0NN2m3S2KzjFc
FbMYjtGorwFoGwGPBBizrW1k0RrIigX4RUsLdtvG3q+Q8ZC12flVY17+I1a07B+NLhqxLgnUK0+/
CwnKrcuT+7AjHkZVSk/04vX/DwYF1qukXJIzogv8qFtpfPVMPSS8fQqqQ6EnXDCSnfZ+GJg4Nvxb
uNmLenHBFn+tIrusgE5L2kkDwCSA/ZShxs4a3XPyuIy8PDnAuqSbyJCzrvhcS2qPum833glul5jm
9kvfHstCgPLcQmCmossoB/XtPj6iHMKP+luIWeWvDD0OccushIv53A3pIwj/44fJwn6yaD8pmhHb
GPQDfE/UVADPmJ1Adj+Dw3JZG/2Lzo6OlMWtDdwaGzxCXCZ4kHpvz71GMsR9T1A1YHl5UrLDOD54
gZqIUGAsSExofTNSNS7Pm0w0Yq3nkzZZHSSMC6Tvt/aiYO5Lb0+6+fi2tMZCMNZed0BEs478Z18z
J9S3PxP7ToZ/YpikwTIMeCWOQFOAJxYM8w3wv+q+dfYLgN0+bHXE0kw41n9WZZYDjgmEQkTzDRvc
CsP8MieuubUZ2af6rSd2Nuz7vteyd6oi2urDvHcI6CSPkDstkJdliSSCeITx+jt9AekLdISXC6oW
zZnoHvNUbafHwJD/os7zEHj7jKfcOQ0dqx64pTA6Yus49WQd1ynK8YZVu+GGg9iT4jpUH1+Rh66W
BKdMb6W16wL/hNQqC6y83FPnIXSOtnmU1O0SOygSBGtdPAYHLEmTdG4dFx1bgeztt0dloKJw7w+a
HsJ34x7ttm7OdHqSDraDM1p1bzIVco+jjsfTwdAPpxxeXfXbvCzZYvxLnLHFLCut49BsTK/60TNh
ACqXP10p4vhHLskMhM2RrLLutda6EHQW2zdE1g8Bb0dP3Uht1h+0Sj7lHc2D+HwS5yKEPo5EIsMr
yaChvD+riMY2kJfK6sFNumK7Mj4TBXdF9kvEXU65nypqqb5LpfrEz92SPxrB/NGuXiQQcJoDDRNd
NNy19Cl5EfDmLOjk/jRH7Dmk/Q/DADlNPdY3TuAEDrxRPg5HOX3/yfNdhncWU2KU8HbO2eyb+cwo
itWCSxZeY9jA74xn5Ow15KZm4aVvKUPo1owywxYeCIRsLFMQjGCJuOhvz6k1QHtVryjpYwco+UeC
rVMonWmFuCUVa7HRTALKzWzaeez68NIepxQbiYDmTGOMkrEjoHoWgNpfU7MNf9mrrlR4q8ICGKaI
YirEgCeeT/lzqdoDb5QVmVe49rRtI71I7fVchAyXFLRRIPlhrBDdwNKVOmV5OpJdvkc8ZEDdZEmt
MsTRshIK80XRowU7SO4StgEkIKSfJyypMpbkPSqdAFEAo+p9tby6R6vG8uCfiA15S/340hAhJtNB
GkvAmW/z4RSpq/VIVFjW8/Bzr+lYjbub8Wew7ZeY0fH3mvmEg1egNZJZO7K7nHQgr/2JFVSt1EfP
AwdsZmOd4SagMZ/04kkbC8qOQ2k5YtebvWcGp1v82o7QpxpEaF7zD600Y8Uc0V4tLYQy28vdplW8
YNrWjxRGdEYqS/nMU6xtOFI7yGIfDGvcE+tc3Q+IJRCelwb4HRK1sHW5AB3vB40XeEQNwagfMeTB
ti4dDMTTALhPv/M3wUH1aEp7QmNAHKHDRuGvQfMZBdyLbDu0h0vutCGY4V3MOOQDS02hmpBUZ4MZ
sLWkVduRbQ9Wje3cJ4jC2Lxiw6LK90KhDTUsiTtQ8JQSc8otcQAbOjZiwRjP9dGGtNDavohRmzKy
/50enXGCTjGAOzjn55u7sV09DZu7cm+e82z8uOXw2c/Ieo3QRATPD6HERnB31XFhh/zWgcvW1oio
wi5qrUJHrs/eLmvaOmt3/5PioUHoqLnEnrkrDPgqgtfYjTs7LJDtuYoMtrTMBsK8kPYBkPKISGwN
req+egcqeg2FCWxVY+Kf2pQCirxlpTJ2M2o4mPuZ42YGed9HEBOnB19f/aRZ3CTUPp1gGkhB7RGc
VoGGmgs2NKbWezWwPo9o1uhA54GoK9VbRrZLB2fhvhXcOemyoHT7XQ1nZIRukbw8nm8iNA75SY2S
/23r6XNcpZs3HNeivXj7j7lAi3gb6BYIx6mcvl+TDeFqTQSfLUphdy1xUQPnE/SiiAvbWv/CZVBn
YBWC8eY03h7mroo6fYrUNb0yb18cIO/MhSRnYy3zSOfHBBTKQb4FPLyTvevLaPqLUnGrhQpcPDbK
h5bkPqbUnlNB/PTJNTsGmQDRsF0+G1ZPWXpzdclBorFRjCvmMQwfvtdtEZecDC7Bs3TQAeVqI/i/
BounqQ//7MxP9Pz73wjgHHWVROClRLnx8lo3yEzr11Eh0qzNKLaMPDN6+8cUKv9WU4sW+tR7z0Ey
0HWzRe16cj9cjVMxYYTna7mTQ0Hn95PsMcZ5bwA4PIbNgY6TPsMANLSQs4TCqAXRlhnze3fvnUiA
uajKdjsJM20Cwph/yglb4Qz3SvcRx5TpF8EutmGDB91EEiOCbkzxzEuwIAzPZiSEM2rSZM9jA18y
FykoavST+5pkAEUgWgKH2+R+e9rdWpYdKpmpKk9RpwGKwzCRu0m4VhwlB8aI6197hTsmNqnBnASe
hkoKtifd2XjMRaAwhBjURFvPGvmYJZjI1Rj8b4wqBdbM/zgjuLKZMG5B4jZ04lUbAIR9JvuSvMMK
9L9nffZMIVoFJXnOrzkLyQVrfLqxoBe2QfdrywpynyGGZigIZ7ubveSO+tdjvwrHAYN50Ndczos6
YxofDltNz7T0Or893Pig5ZsBTNZqgiswvEBpaewp81UKiRVJWDINmay7iJ/G196DAGqflfZNzJNa
VX0nifLGeLIqUeq+Ig+Bh8ixV7qRxUrrK+XMHvwJG6E34RNcGeQXiP4PstM/tC8Q8nk1sA0z8/1/
FGFk6J4SmetTVkjISI8IdwPJw0ucyvOss3ljq1Mej3V1fy0KVR8lrRhR70F/RdtdfjtGq0j8n6xZ
iXVFwiU6rdC1/OzYMnJreJU9fasC5SVur23IKrRUd0fqBaWulbybM8/3pklOXUoOa6gXvJZ+mWTa
JNNMmtha2k/n1dxzr3IwFq4AIBnu5IZLgG3Vw8Ca8t28wKFgWa3A5sFVeqjO4wdslRA4CsxP9N6O
YQJ1GQQDHY6Di/gy8C1X8qr4jRFP0tv0ApQ7bZ6YwONiVjXdaOCbITvJYIRJ3OOC53zJi154RlQN
3yS9+MB7JxTO637qN85gigm95yUQlT1gwJxm0v4ao5eyb2vS2QXEKWTFz8KOm5pflu0AJbctY2/Q
ZhCTAdE1u/Mi7916vx0W4v6eLg/io5BPJu1TQop2hsxTlvMMynwaaZJZgZ3mAV6uYVkeLbug2XnB
aFQ+WO72bVPzw+a8j199rhPaxhztsPwfyvz2VsELcFobFqBEbLzPTZOaNmztBoU+7EfmgN+j37jA
Nt80/aEJchuk8T42pSsQYQNyeT2Pkj1459xIiT3SOSGUyR6khsUWBNxKunfn5p2afRNw1VtArW4y
n8KBwQ1QxY00aJY4k63CXOeA1fYlTYr6cnc6Fd4E57L86Qr0IjO57e1EYYR4FSCWIQCWANtMzjWv
0ToDc1Rujyxy579VHMfFOWwSHdlwWu0Tc8PK7ot8Yk1Gj4kHFIylLlZkkLpHtf+TVeqmHPB1X8Vj
lCUwP2Do0NdgouMMqTICXBom1vpyLLdhixOLVeCFrUwDWbfycsc6XksigSQrW+SxTrId6TSR9bew
F8fnO/eq55pHhR8678FMYvh2QEquuXgFnGWKzj2Z1wyO1q6vf39cjw8SdBTPVZFd1exCMl8cgJ+Z
7ovdwh91smGSiRE3egulYTRZOGUPDwxr6sEZM7bF/h2lwLPCBhFdDN71LBIEHZm/db/8rz4AjjCW
qhLJHMNQMJNkNJ+6MxeykTM93CTkpmsXKpe4NQOTTxEu/v1450zV3SwoMEpbRp4+FXbsJzgXinDc
Kqby0GLp2+v0xfetzedxP0i/sSnvT3dqmevypAcXliFSegwhgNVU+iqY7oR5yclnKqwHDI+TRvkG
FNu2Ly0or7Suz0I/f7WveS0U77v/ai9wSG5ZMhcqKS4N70l9AsCxb8LnvIJqDeYgSc1PWmqWstDe
8MTSvaJc1zH8L1iKhyF5F/0q9j1EDPFBHSEaZHsNBqOxahMuK7mhpmctveRRIZr5SPJkcySpygCv
wObZfk6zI4RCKm6DKuYsDGsPxV5VpYHxtdsJkQm3gJPgnQemDtJW42piFLYHfdeZU1+xDWSRrpga
EtBYmvwzQrw9o5iFnzqgOfLcrc45wcZK6d1onyER5Ei1D06dYEcyrDiKfUM0So0Dy8rJFjRqpvHE
lRxWk8kcfqIVcB+VqSX286P4LkWwWFyIgCCBhN1+sub5HHFQe3H7ufBSFe/SkvG467KQ9qbrfASf
iQH3Q7BVqznHZoapoCHcjR6Q8GoVZ5oFrGO6gW7dU0l5SLtDG/d1W4xenI9jTytiTxvUTgjn7zv9
kRgR+st5uH8yl0hPdenmnwBO8TbfUeNH0Nczh/S1UdVlvRiU94untk4MpzqHWOYHPGpcqJP/y/kl
9BZmLNVBoGvrW20HvonbEUqJYrwavaVsNEHry8ayE7cCvVoUQpxtiGBdn8Lz55lqtSIu0Ji7F3D5
5DZ+NDUG9uHIhsKUznHyqi0/ZIUVVoqVobXJilaZgDdMXpF6gBEPM8y6LL6PRV902DHB0+VxWWd+
SM6PZhmw9vyeB/ywOI1Eep3JgI+6UuRK510fQL1F7waID2VrlP3CC1gCtiGQbwZWaL5kXhsS6KNJ
aRB5y9w2ZvCpHFwLhg9bpPfhv/M880QdTrwrV+FOCghNHdU/2dTuhYrWUzcYBhkENXQF+imOdECa
dBW9o10AnCy1LabPKKd0kIS6fmJFY6oTkBypV8LJvSAo60xJipAMHkO5tPbt1DwoEbFpL87wC7K4
rBaqg8qbcLJnp8ACdlm+ixNdGXrzTq/qff33r/4uWqEO7Z39UAVdgQ6xFeGYKdO+JpKvPgoPYxb2
W3iHZxCD4fwkZ3nUAMCkl+HqC+vmCoi3ExaePb4+kPD5wWYGJVzUwg+MdetHg7T7qQ162lN/4fp3
7LuZ/YuCLHyJowgfbOMgsxvK70qy8VmuKEf1hmRVxCssgB3QLKq1tweAXVyW9UaXPB87d/Hk2FYX
tJJft5GlQ/BjZ/wAPsL0tiUChBLc/V7GwfV1VSHW/MNM1MF3akSP0Y15KcQWbVDpSSMskyZAWJLU
U4i/EVgrCaqsqQu+PaoXFjY3VM6KyCdX29QwwvQ9VzliAI2dZac+Dea8M+QM8+DIPEk/Ws0NmHVM
UTRcdJa7arzpxLWnEGV9v0nVkwHfeys1J7baeqmJJxIo8cvt4Xk7RatjoNxEEacsh+EMbJi3LlJ4
4CL90wKhFAMS6KFOF2A+CK9cvKvh1Kc1N5NV/B7CClH9LEwuMA83hAc0qKJtSCMH372gUusDntZu
C/9c+r1HhKzIGsLrAxJQGLGSZ9Haqsrv74aoD8V2uHZpldm1MNFqr1+/VJnUg2avttFsc/kMvcgd
/KdsCh24KJqqHCYkUuW9NL+IySgfjHS/nzIZR5OP4tMVTYQZiTjMos7jljfZId3qby4nvUW3w+Wv
JT52H2PvlWgtWS8TcVLtcsZ+P+vOAw8sacvc2TBp70+3EJaDsUdpIbEJatncfHvruUQx9IiJgh9K
7lQb6cBkYsSOKrJqRQ9vtm5f2SryNXpFHhPH0AKmT4g/cmXpfCRUpzqqfm2ZDH8sJV7Fpfkt00ex
NdfiI+H+YQjG/lgN6AiA4SGFwuWeYRd1b8JIXpeKXSHWF9ABPkpuLHY51/uTRrumcHazNXfcu9vP
nOd+mRnTw1IzJcGW8tjkmb0H/g97o24iwURwZaMZPnePFJeuNpgWb7sJQlr7B5XKCogb2nJIEyrY
9ISsyA0zg6RfjZpNlaB3f2M3DFui8KVgukSEdBWkEqBDfV5O+xQ0VjysnWHVvoPqTkUE3npTO1wQ
L/hiXbMadr2GXOIdXHFMI8IHWa5Nw2NjPIAXIh45IvStqCC3CmkRj6CRhkwToteoQQ7yFqmLOaHb
QAqdOwCyz5Wz9/aY6kvrpXV9wxCXgA8q4xrQf90IAXXMUhyDAWk/3V4lYiX1SUGOUQ1t9VkQBKHW
A9FbouZ3fAq1znaCcTb9nopgLrXxYYt+Z92vrMHo2xmH5Wqm6ZsPyIt+5IuvsNS/4YQUN7GJhaZ0
d+j+jY9YEFO93RNf9AMQX/2sYqc8n2Ycr97ofvgSsh0ZSWTy0fIY/iE6g/YfPPnczmAavTSi3h+i
suNN7NFMW/tvWMBBs4hlPw7wnlDfM6XSkLKsstxLvacX4oi8/IfepH2BsYlmwgfq5C2C+alITTrr
UtFnFvExq4/IsQKKr3k7i/8SmtJmsSVy8dSSDWJOFktJwvMz4mmiFibd4p0Byzuex5BA9wxPZQ7u
hQF569ZE61HbKZ5mTIhaVYrONJO1wP3TwgMEhAdMukMaSLSFySeTHQSzseBltJrQ4wQDE3tZKmtj
BRdEe/3Mcr0GvCcCfGvWZ7/zTP8DO9wKm7YdvTUJ/3YBtlE7sSLW7oU3qIT6PwuHORXIccOYq8bQ
Iqfdl3lESZjJMl4ekHXVPn9FRGIB4duFIpkiSKylX5yzAeN8HGPC4y8jHPRK7wrJBkcY+NU+w7vz
50blHjzpcNqRgbMo8aJ3CkLJDS3uoDll1JuM5un0G8wjT1cqBhT9wntjFa/63lAf9rdICb9qlH0k
WHOwAPuigkM748uNFuExJIJqKihJ3hqIoRHOXPxs/ujpuw0ePs8fnYSq2cDSzZGi9CV2vI53nhrm
pHn5h0jrBLKGrHstCHIrSlAcCFASp7udxW6zh52oWwcAcOrTcEoY0geNy3DkzNQ6JoXi7FEjnF4y
nAvTmAWIu6AV0AC17gmADRcPQOP7Weayy4kG6Z9TmuqTdyfe2JC2vVWsNt3/m0iHLBoC4uN+VSv2
JiwAIGm1k0iwV04JemlcPcsXgsMoRdyHOl1RjZL/OTT2F8dU70cKdfDdgDYni7B8AQNTPAjj70kl
J4xmS4WKsktehm2qmvAmSzfmLGRCYl79JCFm7n8Fb8RcjceMXi/owDa7K03H5kLqEZ6S10lw4WAF
iwNJeB6Seqmr06bq3dcFaF+t6YPgJSKx6NsUsi22SqAU799Hwn8yJhWgRexNMf9qhyva6Ue84Lf+
NaRZo0MyOdky3bYKQJ+JN+UZ+7+jaJu4yrRXrm8GF8WiT6K6WxDuglKpTvPtt2eR28JSDGYoMkZm
fFZMjuWgAh5JBpbw1JYuo7tP3Ejx9CcQ/hu0sloGIhMdwFWCH9Ro4awSPWpxyw2p9SdnTAeHYtFS
lk9wBCbfd+eTm5SxKi0gKYd9QXnxZtiOzmF4fLagSzWM/+d7mKItHyUySAtqdOi7V/djHN0gfVxQ
XuK/Jd/sMQebVleVuDaBlWDGV3PPnrY0mpCVK8rTHbQ51crDQi7LL7IUhkfXYyWCRy34k8buuwJW
cB/GbKaFkTtOtQhhuhijn5J2hS6/QvUbrYmUGZ1nZsFiBySgev/VQ/Q8AUIUfLZ5dDCiPHlqmM9G
AYIGPMKpoUdunIDDDVUVRhMd2kBzO13XbQRufwQJhU4crzZp0vwlIPtwRAD2eiBqk9KT1/JqJFOC
lvBbX+Ky5SaS5cHnW6aHB6vVd3V8gzMGF+SPICi/v5pCLUQ98BKWZcxFj8WNr1h/ZqueCr6cLNh4
U1JEcC5iC3LaET5bYcnCqdoB7IWQT3c6ALrHKC/fN+u7IT8iOFNEQYGHts+85RwX5IqEKclmLC+K
bg3OVH+YzJ39+Jamh7fJxmVA8XkkpL3Fr+LlvloOYEHoUoq0K+dpUb64D67DAyolOm51/YdDXuv3
oiMo5GitBVw7wFROoeaMl4WVWmT9BehoVyz802TznRYPjgYW71lf+2+v9KOCt/HOY206jnN4Ak0r
NhNtJqQl+oRJlolxsK8ETnXZMRXsXcktGPLqerZVoMAR5ht26hU4TXY7ucr22P9fg89DPZDg3gMw
SS1gSPluj5bcVs66yiTgBSxIBRfOv5N/UqS45a1wOAJnerlRfH/50FTdOH/oN1g1qEqdctuYfkmo
fNOlP9VyDAWjoJHXW8TyGZhvLZB5jNgbuQrYuXQ4+zBBavoiMKHPsI11X/R4SDHnTWcJIQMnLr6i
2ZId/Az9Dbio3XQuiY3uOgHJzie97Zxfq5itIj0QJh1G3tE+NU35LonoSXsLcmL+QVNvmVaxYpzw
L70r7siS3XaPJku3dI/QOEpEceB9TZmGUCHJSXpNBPuE2aoyWdG4n3FvKsbDvGElXQAc7jB2yq7v
8netbPQuWasjRzHk1589xICCHJTejRHfyo8QyPvpCUDFmOViI1Q0GHWa9lQvWknp86K3b5pQmGTD
yTfZHOgog5+c8c3DPT5bC/oDDHxhBQ9d3AilP2SDqXfSlBJp5wRSe9msadjc8pt0TdMY4R1F1/dR
AcC9sxAj6p+58jlfuk4paDSqtEEKcXddOZ4/RBP9B86MupGdMnHOSCxgD/hVwbi25lgIdCa0SrOt
RXyf68KwRZC6mRAtJOuFmjY5J9vCPz3ybqsvf2UrbvqlKHj5PkA1p5UqodMe5JqFbpfWG+hR9jl4
fE17n+ZzQRyNDpEBrLowXof+3TeK9wKBRcaX3JAUiEh9zvGkFzMqWZVAeHDBCMO4BGeIh41IhMJf
Gf5lA73FOXw0WmukOctyyt3WzmwKs6wPcJ6mAGnSExojG24ngFLUfDnneNz6WZPqKHnncujZnXeO
7NW4HzJHsbeKchqrQ2Es+HhsW4inc7ceCdum3VGgI+eGPZXZ5nW91L2dCF1S+V+Jx5LfyLMp6YtA
l4mcuhmg1CyvVVDAgW5tIaupSbCCtgUQc5ayavQWQ7W0qZdu4VdFlCUnBmtNjiK3OBuko0oeh+le
uGZ4pCS8yNH6l1gBayRquVXmvN0i+GzOc9nCYZ4Pd68O+za7+24clQo0faglkPwVJLBpUPNmSNce
ZYEDVPzBpEhDlI9so4Odu6+FQIagQQzEwFRgHT5Gb8jpZeAFYjz7Ob+CZsGeTz74JkplN1AAOb9z
5oF4dwjvl9B9fnlan795waAQ6S7IUEvFNjFZn4uQBufY7z2mVtXhTqV3OF3QocGUPeJnBJQj722J
IHZTKgW2d6KVkUXUL+roKa+VoIkWWOsGOxOTenXyEs3XpRTTNpVq1AnHSgySyoPNY6NS/NMJt6ZH
t1HY+dUgcZior1B3clgpOUYzcoHAK5K+3CqMnb0Zodo7VC4T7aRmrCEdFs+HPkH5yGSu+BSwv1Qu
nAx7wmyLKW0bWuba/n1QXGqGBkoEcqw3c4y8ZlUfiOCBX5F/D4L4JmuuBZ5hDRpCjxqnrC6Ye/Vj
m3nHCJZLZcGGqmav8ncBgqeBCqscpKZOWQ+yXjphOJeDfbExJT6uVmFQqVwpAc+Uz5vQ3iLicNjC
UsNrhYtm44KexsN/n7+2443UjMvQdWBHYzFowBlZ3hf2J/fQdKKTwIo1XHZ13BCY0GXroa581zW0
ZAZpyjVoVisSpaqGBRbblLxraoJ1lQRuzpMm28KmSafOBHmqmMh3D+dDzebGjZvZy6HRnTf5NcPJ
1LSmS3xwB6rB1scrVTrFNe65nxtiOGr8jRFlwuOH2kWynqq1mjGtRnyPRrYGYKvbzEpWavquw2Pq
Q2kDKA5NOyI7iqTfxWySIMGwy3xqMGXT3nEJrZGF3f7TEAVHzLgDCb6DTb6dflye/zS15wMzg0uH
v7byn+sj2DZdijVJV0innwOV3tq3/slc56ioxuBBZYLE/0MlwW8M0QND49xj9xLHl8OBvjFlFeQX
2rjgk6XcMwVlLLNK7saFGH0lI6ezw05icNWLsdAcq3bpv2uhPJwbcnmFPeFA11RrvskRZiYsl6yD
dzQXYV0Vdmm6gevaFskX6GUeGIu/Ir3PsBk1NxDwDek5iM9/CI4wgYjLn+AzWNZTP1tv0itrjOHG
oewu1ob+Pgj/QfN6tNmAPkOUG6IE5bAoySQ2PJz2edAAKJQl6dzLHXNarMYW/ip3zRo3asQN/wFG
FdwIsSkiVfnH+NaUuvxlMtXfA9eFgzimtAjczYNkZOkjxTh/ptuFwj6450tLy1KVJbLb5NJVeWeE
CzjzDomd6x2IBUFNAibhscd3AeR6KDJETi6s0s3oEdt/OFVP9K/rRTMTasB9h5jGhoQYgUV+RYP2
cdnbRR4qtIAsgtBU3ZhOdHrqHPr4hUkjG2UEHjmiSbHQe1oWOHAfJG9cV5hqDiyaiazafMw8nTtG
iJ5fipWTmQRa9N1Wl8JEX0pd8J58Ua9T4kVfimzuVX0f4BqxTROEf1byRRo0WVOfQJlNcEeSiXfp
8cm2n9Mj/rgedKEakPtocv/0tOmSi4k2FIYqKeigi7JvC0P9uFFeIm5eunsGVwsIEoU7Fr0aQ5dx
zJa8iWBoAYdhJbpaddJ6Tm3UI/f6siiY4mFtkqO+niWK1yP7sYUQfUWvIVuP4cgBtucsGSkD76/K
W0d/Yfkr7Bs2zQhx9FgbHNmzVVGyibWn1+A2GIpp+f97g8VgdfFdcJ9M4cRrHxyzQuPQ9bxPMlMu
M/WNPVTp7MNr2DK5fRS8F6TBw0kMTlrM8xmbMIRxg+NZyy9vcLwnTanQvjlqr2sszCfr8dcOBeyh
Bxq+p7TpPP2YC0BlVHiMf1MvTuijiuZ9lQYtY/MDa8KVkI3uELhdsyAPHBPi1OlCgsdCdwm3UI1g
BIQLr6YEgDbp8EWbaSXhgdlX7cyyQErtfx1HKbsimYdOMva1W/UVTFugKa0775VoQ8vCVSYhzM4f
NPiiqhnvSkCe/H0pf85l5xwvp2mjZMSv8XTEJSYZ3/1aSg/JN3qm1Z8qsKKE3h2vT5YADGmpSOFN
g5DfSghMuEBDlSdMWqshr+B6Ijxb+GfrbNJQp+pInnrIxkuL7Dlg9eOXtn06xTLgPRNNdcMH1pEj
AvERHzvnuoVD1uw4PwXX8OKzxMF4Fj0F03yKD2FaU4MkuS3ieBkdRH1DDpsVqKdqtoplrNdjfctM
KXr4pXxDzGyX0I4Sk0LOMil7XRgkenef2akCBPdOdkrmz0QNooY2wxANtVZBpZd1I3KTbOOnDHj8
Dy64cUazGokksdUezQD0YhkOn/9N7ahUWeZNckSL3hV91nm7/aSQniPj9OTuA0vUFz6BwwhPmKu9
0K8u0wQpfnJ11DN/Vc8el9p7To0pdU9/ablQ5LhUND/QgMOkJHreNwUdX3ZC0Gco5aHtQL+h/IgB
FxoQ8R9DZ48aXi3gumRWFE2EYtN59AWZj7hWDwheJxwbJLGcB+WWuXP+jLnel0Y0/w3R+XReS9Uh
jxgilq6jbbv85YoMV/tRjOapZethXedDLgxMsaCh0LopXNC9j1PAkFoBU3BZusufp86XZIiO1ADv
/1CEOOmda+gKeBARBPk1Q9cFyTUefDliavZB8I9wHiAtVDJpPm5zZlTaOTh53XT47rovglzpVC6+
6Fma2w4chWyl86bDnMNJpaRGIRDRjTHku4JCkorv80aR4dxZBt794X3l0QzarqkHblyuSp4b+bmc
J5JiMM3VSNHv8CClAIPRaQDamxE76Mqt/KzSg96h7cQzWjI5f+1YgDicQjr11OA6YLd1GZUEc1xQ
hywsGCV9AYYbiXxCLEBSJJF6vEw18LFv23uxTlJPyY4iReBxMWnkUr4jy/jIZXhSv/vsZo9lAT8D
QAaHzP0vpdrmlszbmqr0RpWkE9Dlf4B90hR3dqBR+QeP3mHiW7PNYq3rVctip6SflRLHv4HxtoVc
Qc98K0eQZJCbxB5WLvTqxzgnTr7mrpAg99kUZErAxtdEfwM7xub0rHLghTBlFsqDdFMdAnDjxrpz
okT6tWys5+6IyT31AM4FCTyv8/ILnuZuOMD59z90hQyGA1astz2pIiN8E2EvjH8BUhUkpOggI1FG
yI4+zEI7IvVI4i9ie4+s2KD4QX3AURfBAMxU0n7SaSopX1+XzMWbVJJy8sCCe12vMykoizlWXMyB
glP8EpX4/iPlPUQT04UGBmIkwvxiUvkGWyuIPI7w9yZrIqSR7lEC5iLwFyU0xSeS4qha9l0KNipi
Z4XxtlrabjC36g3s5GhfpIHvtKSdJ7T5MvkLjNaYtjwMV1yFEX+TjClTpRjQd4tgUs8J5vK/AqBE
ycwBfOk9kXbOrJe7aHZnOAwQsEhpFTqlh3kk+rgKdvJYrWZfGbftotHmFjz979nfzes6+o3/RO91
cbfh/JDaHNL4+Tr3IBT/Htlidc+mcEsiM8uNaAV7JPhAmhkhoC8/qjOPY2HFyJPebjxwud71kt5q
CpVMCZ/QWBtC/2El0/WLhl2aTmEQpGWAZbx2NnhBFce03puFX5E8m/HlyPXer90QY5PyYh39CwNr
ogwUgFp8fyNZEpwk/KCcitisGpUkbz+iaWrCcEHiPOBrX8S/lUzxieHvghKA7k/NWIVtbl2pqqpN
bUgN5wjjdsfn2SLSEsck/VER06P9zOPLfNsjg0hj75GDC7Vd+1E+6PWBXbMR5yNC6l5SGTRVLcLX
2cg8Kz9J6ultSfoRHU6/o+P41/3xGKzWJ8bILtcfWAXgo7Rh2ugKr9xAfOVZNE/FkndTnNay0pAw
hxUzn8ESZ8KS+MMywmydrUIdHAK86coU53h4FopWEo2u2W0WojUy5a10++Y203pI+i4DULkUYKIs
Mekdv/0HZ5PFe179aQjIRBNSYFmXX2yiZudaDhfl6v4C0TzugxKM1qcWneV++05Itizk1mEp8bNh
pPqWmj13+CdIzTZ+XDfHBE0NiYn6x6Ipr5RLQMLoIw27/IKTNy4Q8EETGvOTmOjrEhAGCgeSVewJ
9QLan8BC10ZnG9A9EnXTrntK6zstSudIDgajUGP/C1qZc7WGbpQw+Wtrx11EJ3fivAP/rfvhZJ4E
5fgWnXKbeZpNnKM+CdywrQrOsoYLUnSuxl4g4Y18YagckJWppopnrSBldXi0isS8ZC9ZXVxWs0/L
o0H2e7wfI3CUF49XRvSKkT1e9RSZ4kwIZa/030P8Cri8M8uhNrO8MbaIvxc4qOXxTdALfZbQoYNx
SYppGaL6Y9TOAnQHQtKr/16tTZS8RvT77kAA0KEGDoyEb4k42zpfOpEYqtZTaiZY2ddU5bUYHgfh
YRZHFMjBosdlBDKtlI03CiTb5bTaK6iW/OVhwpIl8lHhTzV/GhiotB4CO5W4Aikc/yShvOqgJN+f
W0KM1vahqK1hUy1akaufuL5d5+ZktJwOMBAnLYKQKeUFLkKdVCLg7e4aRijeLLNHRjQWDTR4sbcx
IrA5Lifj+34hjOF9djEjirE9/j7xoPvZ/a1nNO2Wf4EwALSKo8SPF3kI61G/72earEmW4TRb0xEs
T4ozDvgyErP1ji5g7oplEjVINo0uWqIFzXIQWdjzxLpefFKCBZYTMRm8jKMm7SK9SHZuu9CkAIrZ
Ahwm8UMXASti/kZXZvjGSlkXtOr7MQfJyjUZ+L8vwjZ4U+8pVhgNr+z0yhXD2FpMKMwrT69mhHV7
E3S+kCCx0N/khcUeWtd3IElydbFU/S3kZnxKTTPK84wHmFMFlS+go5YXP1/Ssrj1rnxulcp3MtVV
WKrESCQXsqr6ZKO7ay5YF/I0ZPd/zLqyqNkHQUTd3wvTUUhh8wsz+2hGbZv7n/p+vRODDy1N+YwX
EtdVVw+Vw4u8TnajMkpTnUzjqWpcT46zSqgHpi9POmO2cZc2Sa2aX+zIpNOP/qvjL0yf4sG+1syg
G5f58FVBq1zTNohZ2kZP9Es93JTYsm2YraM7iSyu65mhB/hJ+Vu2fCfRJcEG1/HD4GZ38W3a8kpv
n1XQHFTMqvu9kc9Lv2myQTeBVL+riy/iCg34q3yDfxCuIAYjUz3JPEMQPjZDbouD4Z+w1cCsnIjH
OpVbID5rUszg4wcomUxdz4lSut0dN99/XIjUJjoVNiTKz6ZZ0l7TOTs0IC8Ex+a3WflNNDKs6tv6
+AoIBXg5bqeP+jsCfW5GciQWLAIM5YJX16lcOV+vdAs+hOSEN16vL5UBcRQXr+yANxw4e78s9TtS
D/mQMl6eZWj2vZ/RDzKp8ejkvZ8iryW2QqVPM/wRf/Jf6K2xtdqt1QVFzNwPoLlkk1iGxwJbbPoj
qnU5ltI9cu4B+sZ7uE/lNjv4l8FHj5y0qArXZfxF7dDJgRbNx/pyLHvafyKp2kibTAwcy6OZ9xbq
dXhtE9k1Z3QNehLgICoC/EKtZQqzTi8oJ0sqHg4riZe7mBx+dB4wzKSKuG6kEB262Hkmy1q04EEo
r2nNfTGauwWCRZ2hYokjdfx2ucLfpCropGOJTn+j8GYH4RLSz1GwAvassh/uoypIKPBK2wQQ9eWi
j7ELmRg+kVuyetnUkmPc9rdTPnYRdsrdgJnLlUTlQunk2hlRwW0iBr2B8fqQI7Jb5u7xYswsSYX+
BxKYBY1YgoPB+gFTmE9Cmh93S8wrsXD6hjarGdqPA+MPO1YA5pX/chvKlFi8tRMcr6R7Njpy0XVN
vYx0cJRKYw1ICnPxPiCw7hQL7F9Hop+J3NpprHUp7ixNXMdTGJ4tg8lx7K+ul3NHb1BlfmovUWO4
KPk35ctcPdyGbYpJHQxZ8lcKYJ+TZALEXkruxHYTYKX710HPcsgvXk4oDSLIlDy1TjHKRIncDRsS
0hbTVa1ioNhHM3VlaoPwHoxSksKrjj6WXaoOdpR4M4cKKDkSqFhIo/eOpo7AacJZclDdKqMa2MTe
bXBFyYFBlmo+m27R+206gkxjD56mA2dM+XmrJrArQzWNMxShInzYfP60r2Po+fZjCe7zjPW7cQX6
fAL+vRdnx3TZ2kz9LVQyE7BBJr1xzmijTOt/xgaPmRnQkGhM8iNBkOSLCdE/bq/YG5YO7DbSHH1p
HHCsAGUuadrbJ19nXlsrR+3jAChREdr+yM2WXL7bDf8cHjnKjqTkpTg5SSykXxXFVGolqHQuPEG1
DcA9VsFyTMAhdouXeGLIeeFMiVQlg1ejM50bNCxp5nn8XpSQtC9Zr8r92TCCxKGm9/LT5dl4yZzp
ZJgYV3ZYryUhH/V7KEBwLj+TT45pcnGDBG+i5YlZ5e7Fn4nQ3oaar2WxwLHjCMw8mRVRqc0k794L
QQEZSJYp+tt4viVk0N1PN94PzBAnz960aOrc/34Kj5iNa1APm/L73ijYuIA9gSH8vlshBHhjWqDc
87R3ymtmEpLOLUveYJBpJMs3o4X5BtGwWB/Lt/Z/PrBD4kW/FpKT4W5xwM6do0+jGtXWPn+Kllst
7laweau+FGtBjAzTFhofFndVLWjf2to/s4zcmWGx4LZaPzB0RS7ViODKjmt1sbEJk82LZ2NGhk+/
oDhz1t95sBmDxYXDkIsj6UectCL+R9cOkABjUOXB1sEGXqx/c70rLESvvvHvY9xKtB7FMn1eM09F
huZ23zb+txaU3F6vKt+yxEt7O2a3vv2xIxT6Bx+/c/AJA70fJZ42yMR72+u+h49gvpg20ilfAtws
x8HXoCPbbbOIyzCQg1zkvk/ALXgTCcgcsuOGW2RfmVPnCS439lXYIv3viQOwKmnOdhxVrEx5O+n0
Fo+BBPBpAOHt61p+B89xk+uHGHTg/Ke/e8cwAPbeQcdCHZsKzE+HltB27OXprEUb0dDKiUN/VRdW
6+6dYN7cRXb+gC/TX08Z8p30kI9hNDlKYbMkqz18k8IxzerwSFDks5aD2SYOAHYJBzKMz3kcUUDO
oxEqZMBQvkwTObcCUHM/g6i6DPCvayGvMzSRFZfamoIujAbyiUvxBEQLT1tKT/qpWgIA17BWgiss
MBJeWEvFxQHWSLve1WY9Gz+EvXl8Q1J/i2a5jcmZGT3aAs4L7q2Yv7K2P4eRYAmzbSqV1FLPNob5
SpAwhwqKGk9hPuD9ziyAYUZEV3uAhtqReXsOoZuiUN5+Kr5VO9jMI6e5yHee9H9paUgp5iZfCo3o
9ZHJd+WPuID++W/1nsQ3RBK1pBxTZeYpO7X7WpU4SwhFoyOnM6s9q0OPGrkEuGzFyy5PuX9BhOTa
Wxq7+QjWE0m4sNpC12oOyB9JLPCCVw9gi1WmgS5tCbcDuWs9PjtmtuXnc3RySgczO6PsPdz0vqkl
BdILcghR9XKyk2dDoDte89RC26E5HLX3YIpoc2B70OaCS25loJ+LagMSOIocmOKpK9L5PJScz8od
RsssGwOkcUSw2w5hD3DSvfcMSxjfzrmsAuriL4bbgjCiVRTCEwQPEUcDybyFiSKpXMj4Z8KLPhQm
pHVUfP89kd1vDvO22GQt7KWKk17/SjA6HB0C1DvqXhMUANXX6tv2LkkFN4PVW/u6mVdaV6lGofkA
kwJJT6WbksPblJRmj7KQwcy/lwx31CHKqTGohKOhAHDcQACfONqJuMu+ky0VHHIUlJ8V+p6dr23V
H3Of2N0aUOkqFZyyFDFbZSZ8XBEvcZZQRq8r4MvmFjGDOZROT29OTC2Sq0x+omNQvYm0dDIQXI2T
AEQV3CA7f4xLF/HFHxAIkqXRZK9hxLrvOC/lGeEYCX6qZnn0xR3URPr2RLmLpWFFwvYry3RfGam5
y0Tt1TPCI8yea2m25WwDnWJLO756KULi0BiNmHigdbxxAih7s+JOBDxNkB8oqy1+pEW676h1127h
0d798RJla1PvyqskINx/dYdP+CDYepARHh1dRwx9BAx8Z0jYxVTYHv8vNE/wIgIXo6ZCVsHWSR8g
YPfS9aEEr8LhggqioOgWehCH6g6gfd1Uzhj86szTw7kCegRhQAv1AdW9+N6lAw0a77N7vM3nVYzL
E76TXmU8D++38NIZL1sYIieV0i44jhQ5RKc0jXL3f3p+m1WCX3f2rFg1E5+pl5syJXnJuXHWened
KgQbKZPgcyI+mSWL89ETz8uKoAXDBT5qnl+1P6+458rnusAXcHDtDkI9P8AP9rALsKbZJDql4voE
tAltR3fss9kwEBQOSl00nzttp4jMDQ2zItDdGT6Hoc2sX7Hl2IsWYf6iis0PboBNWrEVXhqF3f4y
Vt9Yt/YW7tzfCTCKOBBmPLMFdVwWZiqtz5En3mshrR2NI8LdXn59352SsSHrUW3Ddu8LVeNMoj1p
Vr4fU3dlHI4OMVFw7ID3LSPyFrIYWtIYXa+hJyUmSJg9lVktwTzKQ0bkM7HKF1LjP0NlfKN2ZBq9
KWBEtyfx8bnC2YnTnuO+7BYQtAdhxVybKAanBVr5nplRc5DpeYJJwocl6tRe0+ewE84f4FN1oPD/
Jp9pgVpSIBppp4VAD/WP0MYSu2h8TG0UltQD79Od2jxJrOah6v8ORMUXQthOFifiD6jv2vgmKqt0
GTiOFp4JGf0L5n3PGFriqYeNu4ux6E8lwyHtj1kXZh4EaV4BJAhSzKHp5JMRYsPUpIY8KUcNqu5I
uSNrXxIV0pVojsAWgRMl6Xnnta9+2+4LaN5ni5iiBBKEHgZh6y1v56jTUw0XLwO6EJnkzjwSnkc4
eZKhMaW0bmjJDDZ0qMWln9wDSyTRdllbsc3y3s5Bx2SGXOJikFCPxQ4U5jk9H0N6EO/lnbKj5dmv
2GRZNYnWHa6y7Eujnmj1hDpwvK32bhHgXRQ2dXvUAKZUC3sQ14y9B7y67zdC2Rf3acSp6mmVzTax
N7caRM9XlqP0dDHAMYVAxoZjh5t1ohNRitJhcnCAcaeBakfVqor4aGKjG8QGUiApbfFH2mpAnpva
YQWyHrIjTGwsHGroAOrVizkBaqdGvqROP4DHIvD+GCbXvuoxLO8Bl07uYUJP2dCARXAKPepfKnY4
amkwq4sUju4kbOXpl1Q/pqa6ZybUiaUOPMzBkj68EfNjq4x7FzNuwruMM5XgSy4r7zexZIpdJYon
XnRhFqBP4FrYfC+pnI6PkqUiUbL9p3LnPC8rYmixwF9sQgVTYmntvMBrhAuaa9CO65SP0vCqdiMx
HKYp2xhJrF129/cJQvVkdX5jIONl/u1decNsghCvh5fnB7NZDg6cIzH/7QvVrXXD0Xiz9rELqKtH
6GIM+RSLVXIBDPHZVqYg5hzL2J6MZ2jPaR8ttWOAxOv9sNfrEfgrfqunCHigcGch4imOkCQG4tc9
BY0DNoK3cbaI2EhSNzFtrYNe5t5gqtgMz8pe4XFCSUumBQDm2FXxAGCPN3Zc9zaIqvBdeMuF5H77
ooQb9Mc3JPg2yIhysWwDS0KXgXFrrJIaZGOkDsDqVZo5Q8h2Vrtqxqwsn29I1UO6D3lOamg895lQ
Soj8lMMTDWliaE7w91N3ELNDxxstGVDf09DZjduQF1CzVbFpwp6Y8rIin1SIG+RbnNXgKwaxX5TM
6HDm1DeubmZxyGjLcVStD7bmoPCAmhX1KLxVx/dAkDd60NyC/U4yV0Hjttc0bnfV7IyeM3eMrYgL
MVflzMM/JTlSOIYtVVR1P2ZF5PQrN4GS9Nb1MueeNWyM1C2ZGLEnDeEvF4mj1O1wKjmIiAnbUXZo
pddoVGJdcQQNu/r6GSXLZK9WU5S26QeDMd/+gHAtLYzba1i3Flqr8uj9rfu5TB3F985YSihsC+r4
Fb4RGEq+Ha/S417JfF9cVi46VCOtIFeLsatDiJ3XW3tQUdIxDd8Y9vV1QR/8ZMaOeaUp8qNSkVxL
WniRPmemXI47l2Lz+psl5OZp0VqmfQ91vzFakKDpZ5khv4qyz3zOzSn2Rd5f8f1UaQBNK0JKAR9V
N/ZyYUX76Ih5aGrR/9jYxdieTsSrmqHXtgDAF9cI8R/khKt4M8QtBdpfAcQlR2zMPd9gSFt3kpaD
Pja6TbPNOQXJ2tjNNM9LiMJZuK/Ojkpk5hf8TqVVovHFncAcWIXYluZyheDR6Rw08zPQYBk9psuM
PuKk1LF/JEctOxnzOqmLig2+HgUPDDeQ+hyBVUxRogH4jjoUBhd4k6OthKMUj/hCJm8N6E6PsIFZ
aEmdDiXzWylD4hJimD4iiIY0flbtwS1yyWcWSVeuJY8TSTSlgWPU2i2frXYhclOMytKOQ4NxZ2ei
3DZMTUuwz3BehEG61hpiaD1MrwwgdMsUD8MTvoheIsLxBmJoGqBI6j6uh3dChePiwqdvKwyXOOnr
B4vgwPzXVz70mEbL4OI/k1n5UOme5hb4lFVorcx1uB2ZyWKaYjXdR7nxU43QnRonNIDLf6tsMDUI
RnGj2yr43YgEAU/VjHxLuNzqvwCLJhuwtp0Dff9MVwU1Pkni7GdHdDziJnZ5Qx/E57G1xGlshSZG
dl+hsCwd75/u0qkBLYiR7zOO32mC7DeL3u9uimLkeCC3Sg4ulL3nCzUtapczHW/Uk1BJUbrUHBEZ
G+UV1BVCyYBFDozqTO5vvQ1vkGFEGThWNQPRQ6JeziBmlL15obRV5+Gdgc1SQUyr+UAOLk/plbmn
5gVDNeG+/0WbpGeHqqjTVimWB8usk/PvH1K5eBPRXJB6MoOrZazximowS4HfIAA1F3OnT8snIUJK
np+XYcppuNbvPilGR2CdztTDokb/5gpU6cNc+nswpc5iDvZ4NqnwSCuIPZhb9R14ab2UKGT0x3os
MXb8UW4fL8AhxvYmhPkXuDTr2y33ureQULekXebsF50dfwCkvRcXfulFSzizvjrw1CQzr7yt8QPz
0WWu4xMepab2vWGBt6lxWvSRMTjYz0xAwSD9IqoBxxE5isU6DwsGiPAmh396odXq5avIb0cglKb4
FcYGw2h/bnyCt5b7112nK5MM1oToMvLUzY+5vaRpWIrZX8Wgz6hzziu0oyfOKTDSWDXy0bMfxEuc
AtQEUGPtIoQADE5XZCwWfUbFjVr9eNdCLoR8F1P6/kKn35xj9RKsq9UUgQBo/q4RFokaEnxcQO4P
dDiF0RUCtWU36+tMJkgvNeAQBhN6i15QK14sP8OSeRdIzELQlZvlrDXFGuY3/9UuMH9RrGWRhO2N
5ZHZ1kp0/WhqCzflM7fDIIArmTol5YyQhjB5a98o2wYFfLpEmpoelx3dmNBgXWs0yIdW4Efx4+8T
aOq/ijOwiUcPtYS7q/W6lR+lMUqC4QEu1epsVP3kIZxlJV2lDCZz0ZJylx9EFXRpV9BtWiy1FcNM
s5/nP4ObJJ72SADvcW4zY0rXfuPMZA2iiwx4rcluFDEpPfKZEIRxNUZeqo316Ekd71OZHydvJJd9
77nDhN+s5+xd+XsyV2SOOY3QJMJ7E2qNHZjQ1T3e/W2/puKPGAl7xTdU9ac4aAggcU+dEuP+Rejh
oIlb+pp9ZK4wMBMaGZpAvpI/qm7keQbEUwmPPu86iuqunAmDfgzzG5cjUw9Z+iseJDfi+g4StT5z
AjNz/0pI1QQ9qDYmnC4eNTl1hBAgnYFvrfUZPU8gUDZPClbZmcahb2pHynP76t8fvLaxW0B+2QDc
6v12DKsYBYh3K2cudWxZrFccpqdjLZoDmV45CQgn6dCFtfY2vo1HVjJt5iTLrS41rL0BrQrimIh5
eqNIxkYeLMSi35ZCJyVfiHgmGKpW1CoVpZc0Yikbyr5BKhTabMObQHQA7HzXl5r94BWO5E4Xlgv1
nDSWD+kkgw5oWBkCZfYZHErt3KsyXi1cj1JOEtVtaw6gtcPz73d5wOBmbsYEbE+SBSbrygHs7X5E
J7KTKxNSLX6hg069XpPaNF12qQylW7IxHQb1xa+h3S3s2rpQttmaC/JixcadspHqY9Y/xaO3aVtH
7+xnog3Xujg4jEKsV/JEo3Ep/iQV9mTDUcOzt2sJ3+bv8HCDUdQkmlWF+rgmz89H54Zebg+xMfGp
GU4IjIXg/t61RO41Qprjh6RGh7wv2hPmfioHIGsDoD07AqJeLysb8GpEHIOnAxilTdSU//+OyQ1T
N7LsuESSNKBKFSK1spjgi8rAVcH6G0PoyX2qe9ixM0PoqkMuCq+PsaUcJ+DJ5WMs5zDhnb4nWThB
5TE6kRtCclhPPuI5cRQ9rOY/y+a+N7ZDrj+Izr1nGZBMNPiodBDoGm8TgN3slGgR0txEFJwaboYd
FoIk13q6lQ0DhTn7wqjtP+MWqC/R8nK5U/EiZeJltEaPxY7rqDqshoa6lVRqAbaZnPoAofmlnd8g
5wKtOk5lO33rP6BbXePZmoZBUUk454q/ew8mIuHRImL4cuBgki4bdpukqxIo5NCw+MO0iaSkS96V
ElL7UphmWPSROlOfzHYoVvhOj8N8cXd+gnBXju8H7kfskBgBwpTJAKZ9irLndLBA4eYnFxVPlN5X
CjdKb5kaCuEVIoLqxTN6EGML7wip4+yof8lVVe4d+D8qPmiZUQJPAslLbIuhDcfuCDfshg6eyUC1
jBQOflaeDwjVrWRqvwPXh7lHQlNyt/PWGv0gmhn3YNMc0/RMNwS1HXQqfMR5Cks8DbwDIeoy5fIZ
BOQW5TEH+GCaP8QBxYMWBByM0mpI/j8ejT9tVnMQv3NoR+spI5EpmGL2iyAlw+tWk+QNsqoiLytu
DxITe8NJ0UhNBSAtX9HBtxXc5pswhCMztpFnU8MZU5EzoIsD4y8mqY9NOQq3naquBcIe9vg6wNjh
fWuEVQrKy8RBbSOkPNH9/DqJDev1XrL3GqQkR6ApVw+mK31wcuAKHeOO3DNmGjUm24UYnAC/QEAc
0P6TeuFwxzkv8mfrjVnbYvdW3pAcF3C259AUKSk5VHOFVAliEtwt7e7ujtXC0n2IijvULPwwS1s1
DC0POh2Vnl2cazVTNkWk9GZkT16K1H7H7gJFfFu8a9U0A38O2VGm9vd3ngqUu0AG2GJogt3qs8I8
yJGD0zYWlYweJyEIneIYbJpOc/GaJ+Eho9FUueHnc4qNd8N2MUNT+L3o90APiAHA/lLsDCI2ImNG
/NIwgzjn7EFl12E0zU/JvKPijoTTsiUVVwzeinzAsd+aw932Lxsk2s7vagp3IfSJB7sta1gwiPA2
o7EEqyOJ/xONC1IwbrwsMxzta5IQCzqC6W/1kuq+RX+OunN8ySHCFiqAMCUMHEJEjhVOMxyujoyK
+Zx9midhuPfluumtOZAq51lnXzdJzB9Yw96M8jltAwjrvQcSz5fWaao1w4+Zvv/ukc/2/fRoG6oi
U7Cw0CIs3tryzJ9Hv6Ud8cAL11OjiHV0GkQ+aHMH5FlHZCiHzyx7ZvFSQs23O5Z4q9/JhlMDH5B+
ay7aTow0Y1zTScGz8x1H9tgdJyJ0WEBvaj7HewGuEX5FdJHzSXRcxIqukpIr8UEq5KemCHP4SF0l
InxcS5FtCpSGvzMnFvp8FFbHkllar4+hiPN3jI9/41hZMycaGYjUGaxyf26S+WqQKSI8R+2unegB
7g5VUgSu9c6xRyPbsWthEespTf2F0DxRALcYwF9fKjNCbxlMEVrxo0h0BZ4FWo4Mb0xRmY9nWg0g
4Ybt8Mx85AEoVyvoXexUlvzycxZcIe/9h8ExFNi4f9h9SVdZ2CvD8AIEqNwGTp6cx26MdBJAafib
oj57CIotymljtxs2nAdxAGgkAggVTNzEmeJ7gGKnpmfux1hPXspmzRn1gUbAZdVK2nH8EaJI+LFh
/nqR7akYGsaeswY4A7Huqr9VgP4Tu4fvRCOUy9F9DTjWgNL9L9wYiUq31AQjfQAZPwujj9FCHxT3
KThc4/3YRmhOXgZhlcxLFboTEWPaPpump1eC+WEPQ18Pwk5QRTR9ctYCSl4sPS9uYD9i10km/bix
rrw5e5iqcP0e8mv9CusD0YedmYWXSBBWEGKyMSyDxt/JidZHZuw1tNYs+T02rtKGUo3kb0ASD/SE
yZjTvbkQSo9pUTYL0hrNVDG3b7O6dxvbpHIbebDAkCuNCbrJwjNFSLT1X1+IKQPSLFoDMUHfMQO8
/fjofAt9mQGIooT6FvcwiPaqaTyTTPDGD3ygKu3FJEVKZlTNT1w/VUW1NGX9/8SrgIz+YbP4lszr
P25K3jD7/AlTraOwyY5lDZYA5NvxI/l+AFl+t5IzbjLFtwb2AU1wyuU5UqfTvEYIA74GtNSzR8os
NqDvztT3MDcHhRwqKLL1nyEIo9x8AueMSBGLUIafKi4AqeabF6KjH8WBzqmE3/JnWeRQ1vCXClcZ
mXbLNqjAAhceNRNgr7/zvlc1cC/GAfN5NPADI6O0kSuZbBp08LEYDtI7bipqrBi47G2b+T1aTyjB
h1mkmNszcv0faFJ2FUHyoO3fgghklmnWKfpUMiWl5DwZMfY7FTMszTD8zrED8Q+g/4T1LrY6IxIP
OdVF7L7BhScmHvDrdEDBNdD8jchB4t7Gjp4kOJNNVbhYF0oobZGfDVXnyG7oR665WOmLr0UlbFL6
P/F17uawlmMlG0y84OrSNLXvhY+QIY+PLX1DrqyIW5e+YL3SVETgY7VcQLVARwqKRWUBnq2jMVsz
e517MBoqtAfinmbjfl6gW/0iFxvNji0qK9c6kJnKxg9DxdQi2EqqIBEIV9oVHMoib7mrfIoFVLav
fG0BLzJcnkxG9UasJpiAF5oRTmC59ZBF/UlX94l7iAf1Nv93U3x2aBZtfQzjCeNJpYt10TqCn7iL
/i3D79wLBTvwGh3xnWSeR2q7mDr7+NVZ2Yuvqnk+IYMskIOn1sKk8mfBfmbhY0uvDMzqtHwQH5vi
iCx+Gcg0LYIUtdmlQnGj1/MkZ9k3z14FRX6F5ho/HWJLxCe0oN+w+SmaT1Sd1umVBxvaxS3ZVfHf
0NXzC3ByGAamLcR3WZw2SsvmuFeg3SK5Z6Jlb8gHA+j9tw9+7w+fFIicDW1aHgIjn3ByGIGAjRmI
diqKz6L61+wuDJx1roogZU3kb+pty6tNdeHTKVfJcPtlyvDSx5os6krliBybsePTeO1MugJixydI
MFbzVgJbY536DvuXFkQdr+XuILD7AsyahPmTjcL2dBCq8K27g4aFiEqzgqnzwh7fpR/AXJtGjpqh
7kutEQKCEOw+KIXYvDUMKPXrhanj5PB2kxmbp0aQfNCg47hxa2Q/o63/s8V6/n9mMOxBVyI7Bkz3
37Nl0Gg4XqZJODc6Ghh6XL/8jjHjn8MvcS56pBNP3o/0rDkhP0QrmwHO5KpBkvzy/xkEoG5vLL+D
XDDnpKg+XpUvRjinY3n7z8FzRFpotpQGdxnecsEHZQ49qtMEilSMT6rHbzHE8+iX6mi2CYcUgDV8
gvIA9JWdfFVqyXUGE0zpjh12FeQN+P5dhICtwVLkhHspk9r8hUzTIo7xE8jQg+C52FPMta0JCluB
uXmLUI/ZMP0jr20BfdSXjHeOXwW6C3yNxSAhYX9RpSj7zyfoYBlsqvfz8bEk5MBw1eXKwPHRh0QD
+k/qCpzSB+DS4BXk8Tzn4Zbub6AMmmLpKpDKoEbVTM7MvJhBFQK+s2aaI6HNJR5yMkXKKy/KzjCi
vJRnNNraE018CJwxYZUnCfKDIBKGDQDnLBcqmhZcR5DGv5OaN7H0TyavA9uDmTjLlxu3n8AIXZaw
JY9AZ884+Xl2Q/8YA3Tk6+IwBBxW5WBl0BibTbx8DzMlmrs4jfZ3DpVhwrPUkGjxua488FA59FHR
RyBv/dvo5DX7KnmxIpK8dOgoQVwzGze5HNV9mCCDcsxq+iS59IWQBCNm6rt6msYeOoAaMucee5ut
IAq/ZmXVMsejL7Dt5jSNM4lGQymxgmk1OCVvRjFmz5mxCjle9Y8J7coDd6gTkcQu5UhMp/5+1XSh
oDgBBjs589VnvEd0A+BmAi0IXHTC8FsH5feXa0LDTCiUM88m1+Q6TgN5V7b1Ip1CJ7bld6wCr8zC
emyzgZrNgn0xGK7+itpwlQrgSySmzHMc2bYSftz2P+4qFXaNOwnyd7+KJJwLOcW3uOAeTwdc1baN
l8v4condLrVVjAMBWfUXlLu5Yc/U+abFuD0DEiViW3MU+rTf1620w/NY9ieiQlP1VPQFm3v5SsUF
3f+NIL+r961hrfvLPqGVJp6ijQHOeqPwJGIbfW+H+qqvBimAUchH6CunLfv6IAhzKxjgMJWgjVT0
A3OgDEyUimbIFwv7HlUT5Vu1RXtoRMTxcef8iMDUjpVHyRJx2GrAS0qui9BGcK5t0M0BgQfcNQ0k
bFnAmxPS3ftVa6kWOpePjgT5xVjcUlLuVRxcDKDstMI7URQmiNEH8OzKBecaRqpHt600TTZXzeOr
87fXNjWWGC8t7JECp/EsVoXWaPcj89K+hFlmVW6lUibFxewXmMVoQnwLjjQfYr0EhDi61fHYVI/+
Mw2dLQt/gGV4Jfqbx+ac7pWmNKA6iWrPceA8WR6T7Iuk2SDrEt0W29X15tNAT69uMhFp/L7Hk9uJ
mtKmnNawGRdIdDeaVuo9OxF3fF0MoJtQRicbHBkQ3KKB4S3qLpo5k/pwfpWJ9+Atfrv9O+Y4QPdl
RA5pgZcTlDBhaqxpOipUw5WcIlsBT9gIRdBU6mYVUNBiGmrJ6MWa59HoAL4ke4fBTKflPItu0hVg
0m0X9qWf1yFdilmf8+D1nChY8wsDlRnlHa2UsAn9SgDT12X3fPpEtEqiV9TQyEgBI00uuFvZI5W+
HTKtIhkOMGXqk7qzxbo/pYMtJFfpIgJis/OFd3KWSLf7NavkNMZPFvB6DrZlRUFo9KXg17DchTRn
EOmu2Ml4AlHEOoWdp2CsizX/GZ/OK+9vUCRse+zl+ZYfpe/EGvGI894rOnZJGS1247ku0O0nVsBo
aEh+H0dKR20BuBXbhamDQGghl/5UKeoCZimy6G5VvUbRfQSS1YeKrKTpipXgPL5XDC0YC/+9ps+1
A6ptFxDKCNmdsWU2ODKbz2L1Io052drY3JWKEQmmus2a51XdBg2EKTvMOi/0/EQK7PyMQPenfnYC
t0Q2et0E9GeDYMY4hx7ABTgUmWhnlU44m966muaWe6YfkPU0ZGHb+NY+9d1HFWCIaBtkB7u23SA5
Hp6n6vKU66q8wsNYuDefcyAyWkWT5eUxcbKJMNSUWfxmrnwYkyILdN9IOLQqbawDBhLK3KREbumA
IawtfNbK9QkhpBmAjPi6KmZ1JljiOlvaezGDDJHTiWsA+vE/uC3L+ay8Ook5Q4gNDjbzwEFjBOwc
TlZzkVEgivlEhwbT351h+mNJgJubGPDOfY1loAKIE2ANmjf706/7HidTUvJlkYhaHfawWAV6BYo9
8aJmqZu7vjlH8D3zzouCn4hfsqgKBPKm6V1JFUf9o3EBGGtCGElfudn8KY3Pqbp5ub4tF1wLvrcP
gkvhklPfIddYlm0nN9DfDmU+nD36l+Eo2FGtEgM0a3UGAlb4PMYOMBsTW5SwJ61JiaSgsn6kC8Ka
RpwRkW7oEA0+cOZY/3E76Vb0qPoKv8ggd/U9+OU6JVCaYiubwpX3cBXh3894wn9SAeUXCOwpKxjo
gFFFS9TGZOg3BTh6rpqY9KSDlfqfYJLhNn4QpBifS7kiv4ngxviCf8x3KKRKmB4Y9TTWTdK1ofDU
Dk6UZ3oxnLB+CLM5phhVDlZzsUQC12uIsuy9Da2N+jO9acjthfimPrNdEip0u7to2SsLCpatVfnA
Yh4ul7Eb5m+oXG37Nc/tGLgXcXBSGBgySJkGijbAT0TBMxJQJaOI4yxCHv4U50R+Kh+sADZWYX2Q
lK1kSfbJz0osMdCduuUXzcTsnhOOr5aQp06G9vKpfppw6IT1M9X3ij8t8+v4wTicFXEItgQrv0vh
gW53um6NStXyZH8G5GVcrzQvonrqFAKWNG/GbVN0d29PmR46vreKsM2KgDVwRk6zyS28TXltSHJg
T59n53H15M7AootGq8D0dQU2aAIazWyhIA875l9Poldh0tpsbjjx4Gjn6km2jksXwyOCrKyTI+P4
SGJ+poV1CZcdiBYdUG7h5wRLA8ROM4BYqr/bDdFm5ZlguWMTIWn0AUrvTZaw2P5iunCHJR6Lg4v3
WBo/FiDskH6MIYhv0koCHIe+5Me+gA3MXh1TLtXDPdAszgNgn+tUvHoRMITQhc6cRrZnnOhdTFEs
0KfW3+UejoiX6znX8A6D+54GFM2rPrLr3VyIQWu/j6xiacXxkmoJ/AEvSNp05mu7mEfj3cvaztg3
Lr3sNn3HTsHb1uz2MRo5n2A8esArStGsCB6HQCTp7TSPkVLAGoThza4JJJMO1BYD+5LCf2S0nQsF
ADlI85kKkEkKgmvhjOBvYK5iEdctMkOJIaQe/whETA/sPxjO5YaYexRxQJ8+aICmpXarr6BsPxOM
O0LrNd63FBGwaHyXDLd5MiheLvw7a6uFkqOWXQnvYllKAQZjrsxMYyOcDQVbecX1x9fQ3FdHQPUb
IfzonuFZm2sGVgbiv+Cr8y3vqv9SyK2ND0huqBhY6ULe6metqJE+BLhgEHn7quFleSvmlBbq3LEK
vSSM0oNCGWQhn463CIYCO5CvF8Jolju7yn3F4m6clWW4Q+YWgOpbB+2qZRjjx9fq+ksHCz2r5H7K
jULZ6vqDwyv3fzk1v7RrvlBC35MwMuyeUyGItC5xnywhAnohyulkKknx2K8w3qtauq3lQDk6mZfM
y8ToGRT8ZYyLQEaMGXFBYB0qwc0GIscVC5HQcRjxHegJsYhXNLR8QFkX8Afz1NFA/2Bw7clykNe4
WE42KimtHYA8pORAjnwe8QhoeMZPVuupXs31XfeZVdCr9AFiY7Qv+Mw/OCQadHOVIpWlhDikenY1
gKEDeJbIez8eq9xXYtBPIT1eQXb9VKK7tsiMKqttB6kjRIjUFQ3t9e4c7XoFy0PwxavSPuNj+7wG
a/GUsGldawkUB3epgHtzHR7Jc66zgnrez2bYMcOitW1A49+uBoT+AYV8O2bnoeAqaGoznzTHVHAH
afza/NHix8sIVQlxbGYrCWv8B50XGMmDr7tUezLMjyoufc5lHvt5ZzoqqxLME0FiPjE6Gww7gLqn
EQlKI85grdThwDZs2wq1SIiQFB2GscgyLEJrFtp6JZVcnTxuG9dwL/THmn78tiPh63nRT0cPn5h5
cFQtWGjg6I3508z8BeyAuHDQOYgKfWXidslRKHfhQVQBzbx73CriNCNZafDmDUMiVGrkdZ98mZFE
oVZyJKLQBzrF2sjjBU8xHNmTrPW9lxO6EydH36Z0ATHVILN5Qydl2hZtZrcaAbhghXq2DJUvlHl/
CntwP1XUOEExgGlSzUECesxWBKNh48A0v1OL5myWK6SGSJ/oX0ohHUJ2h1C+pYtiJYJvtyuV/1Tn
98mYdJc7p70h7+ILn1yi4UqxUVBdo/hSSFHUgYiUiY+5BDKOi0GA32F0B9fmMV/7hTmH4nQrU9HR
r4u/4D32eGhRJUNLWXsxQ+IRZZE46THSUAs2PpwSXG2XnXT1TreoUfKRunll7HQuHeMlVGIJdMhP
aBG7+kLQHBafYAi9rEo1Rd+E2+nmU3HIfB7xNnQEOCIVVdGvtek/JZaEs6eB+D0SAf9Q0zPBfr2H
YjcpsgYUUMKiIbWdy1nqNv0Sdxfy2Ksbb+KhqVmRjgXxzIXHTLrv2swIzXr/uNxdcdpjA/wKm2Zl
n4dqKbz5lApe7oUxVpKLW3RUzjTbM5rqRBoDxeNzpMuLHnlDF9FrvS+6xEvS/S4okS8yfRwpwbvB
BfMPbNwkFNr4oxSLWHyB6F4HEgimX9dzioCyizV7FSeH+XDh3ZEPfiYHzX6qOvl7pwoVF3oU0nYf
Ytkfix4nNO+7AAhiksQrJp7vtA2Y5dnp+/hLfwU4s2Ltuj1kDEoJoHoVGQFm1tKMNLFQrJtBUwwt
Ta6bqdULhLQaCPnmcSgHwK9YLv+Uc9U1u8rtDBqlAFz60NRuFWO8owJhJ4j8uAhbdWE1C3oVtl7q
xTNFrgEH99gWBWqmc8ZStatH+xpCSgRoS4AuNC7m79SfToFNtBJNXzE5g8OzQZiPDHHrYSQjDnSe
fpcbWInzrAhSZtsRLvyprr3iFg3L7xf2A9dTW5+60BwTz1Aqvb4sQLMkgHJ7o36ST0vaWzjhC5hG
9k1wKKcsGTHVmSQ0T9V2kdy6TN/EolUByzhyV0MsB9Z3agk34WjGGhvh64IRR5iPiLpHKeu0x/XQ
XuDWSA18VV/q3VbsMiTTSeRw+c6TTITHzVEjx2iUgEPiyWd41RJsScH/jd+kVSxGkr0/3PmrInc1
yHljJE6jPOFCfA+UdtcNuf+UZireJ52TqqzGLjAxyrLezvuQ9w+dWEF3BJhunR/iqjs9iuOTn4If
zCINZYCVFMcKIDfU5RMv2m6pAUqWNth/tcLKAJ35aRJglBxwBKOToZPAj9O+bSwa0HA8qYBwJUEp
ngPMVKjblxfT3g7ypeEqeYeUACKJjjKNJmNY5mWVP62+7Uziorz0k4ZpdbeokKmkb+N09iroL2J0
pRAfuQ+H0v0PauqMdshPzOoPBt+6H9ZZIZhiVcX/bDCxvmlJPHxuJDMsLJ/o2tAejMSfKw3a82t4
RqOU4YYmj6Cj5xbDN8Ljaahu+9qAUyJX2PW7tgL/smvyHflUZNoPqFotkFoqS3NZRQKHHwC9/THt
VOOUYBBPv4eTEBUnK3+KCFzKwcAZTYRKO4zMavkWScqahdi05OnjJPqlCczaZ5Bn6FT/AHmBjU3V
dO0k9xPgxdoaPPVAeAMl43Xjsi79+e2827TBHDrPJ47NdwSjs2pDsjpQWk3BQuL0yMkU4x6VzKBF
5LNwXV5TUjZPtYmYTYOiWQvBuwQ/Zc5zSbMBMugFMECTFa/DdBr60L5zY1wEnxkPw/KHRykiZsGI
hw0jWsLEimuqoun/i7LYBp1p7lOK14OK2pDu+gNBj4YJ5P4fddBNTegbEqgzRCvCt5zAJfolAMD1
f8yW8IlYh/UeINJL6xXw48gjJYO+H1LGGp8yzbMGRYyLzfdHeqZn6rkHtYopLyUj098hNRvDt64w
4SggxkiAVO1ZlGBq1yRm04x0iMB9Z6/TW1qOWsf3YLzo70GQ6oYJS4UWwLSR2Bv3OzrD7DA0mrVM
PZNUo8ZyjIWKZLOV49mqQzYZGtm7eRx72WeBI56fzS5BdTTeVcY0xmYWJpDYQ8tBiqgXPVNxSNpk
njPrSPLy4f94dGHPUrM0W1dsNZcvdZ5NkPZU4p2sX2pcpfyqiu9YCrMktdZgdJ1THmhXjlpF7gVz
yCDeq1F/XfcxDtQ84v/8BeH8j7OJ1SQJ3jpa9JRNgg5WUOEcxBTfjv/6e/XBmHyC/EI7YPbcm+Fv
XpUNfCHlwZNFJ64j6NSGug0jCfiDkNhA7d+j48ovHHvvMbgXPgOihtxuQZNDU/Jx2hw08BcjQHEb
H0pMdam8IqeeKqMlI7r4oRZSRMUxgD01rdWAE/RtQT3IO9TXNuErqZOwCOrIlE+/GpqvmQES1Fmo
YiS55cnDwKzc2nNwnl5UyiNrNd83vNngwP2lhuHmNKkWgNnhafaGTVBlJhOuykawSpPIWPpXfstn
kjUNKAUjqYIJJTXY1hRjItQLF118MPl9dhmDTiRUIRmNEWBqt3kPEOD/kC5BlJWusK5PrcEuECX8
hNo0e/5hLSXlAZMer6YYkYwIMjih0Ji+LrpRic/z996hhTyXEu4sFvKqMkvpOCqczqvqBL2aI+LD
k5/W6wKDldVr5g0kEOrr/vzJiTvDQtkrN0PmkAWSYWrWt+oSEZP0Uo5hQHC12lQiY6h9xXsKfiM9
RRjyx/KryHZZ8QJ62Jl25RKlWExxcMy+rz9Iu0kBUlv/23lnHNP3xnpin/KfTZkfsNqw0ghB8bWR
yt1zoOqotPx6u+bkZK7yTeBs07BWZEXtbhowb+NrEOpultsWAyX6TXhSlIoLqkGedFDd38q9D3+Z
B6F6/93I3kKC4e65NXxZANd4JrpBuvHbA8klqIZ9W/7vT8WvtnelZP3c+3kYcBSyejwB3OyjQKXf
KejV8lIilq4npCdfnMiQUK9lDGN+9mZC/TuXpPT5UKJ6Y380ZlzJz62Y4zIHF2gS/9kYNNfR8z/D
akdBNWu3hJzPUzMWJIdzD2SeA5ArOzbO8D3qxBon+WlmswzGTV4prujSjTpQIyioZgFqEyCYvGLh
9FS+gfAvDEcby1Vn65PBUt7JjW3coYWYMbo6zs5SKhMLMhTGUK/doXDw2cqoQhvkDb4OZ/eisJbB
PUfh5eFSdeQIJaxxiHJ3c7z1pIiu1mYugmMD7fGKYPRNnFZRj9ZKRLAZk7yR/TMtmlYDXpm1W/7T
XtQ94Hit5gTUmqdgPzUstnMXGHvDGG3FbZovRzCCB9Vm1T8gx2YIKPyfudyR007OtptagBqAx5X4
+e9rF4eTu2aaRFtTDSZaW60aXU1ukmSvHKuwdHZxPZsNBVVAQ1YjUnPhTfgqdUt3tHcpuHROd5Nf
tL0343QMeHprO1z9xnogKavU5HWbgvxEsBBHmNSCaDvNimY0eJyuRODxFB7UidEKAYRBNFNy+7uz
/k/x9Sa2aDhutn+l9NYIrkD7IH8acRGS0WFMOu6oplekAajvVfb/+qdHpuU3h/WkJlNvuFWqGHDa
6UooR+I7H8HLlnwLAn9RZ/7OpKQjwcizBFAbUueB52XRlWt2MxoZVqH7hyv39xA7TcpHDhfolN8z
Yft+OWFu92EgpIqpE/G9iq6qMQCv59lYmEEFKg2/OdFennYeFRoiFxxX1QDvq3zfE0Hw0xRaG8mZ
E1iMgRFklBKtgtjBlO4AwCxaYfmNtTucKMf1Wou4j7Q3OBMmdzzH0TSdDmDaGQDSbFnS1gmxhb0V
ILylhMoDlkPWSsdO0fsY5ngbtlKQp9BeNWhsb5BxXEJ276aEW9sFmz/75oktSkYSnrV1s2CSdXa7
87RetXMlV4+/HMnnWVG8IyMNspE83sOGFRDuStYOYH2xpGFwSSUFhhbOp4X6gY1HNTJnvHZ7k0Fy
lRJfgbHAsBHI8Z1Nc6WsD8oCFj/yNvOTKmkRrfHvEtHxvLOECF0Eg8dXEUevDxuN9fC45WzMU0AT
uoN7HjquzH4w0LNMEtzy7U/Zo4p/ovhc4fItlULChMQD60TWXDWDHv56jMOEUqyOl0U+OUZ8n0XN
vDbV4NYxxuX3I1kmD4ocnqzVX+/s2iZ4d4SOHb7s4y2OwtNNsNRArGCC+hFje3hA2Jq7/VktN6BE
wsXZAYC+tdb2fPsGklnHaF67ChgS3ES/TW0tw5wv6XjHF9alg/6KdFmOaTTLU8cVc/7U4r2ei5Jn
eYVyBGEmBfFBVNXLlhgREqgzoCL0kmHvxUu/4zhEEmgKQOimwClvxbQ4H7FcwYE0QJ93sjPg5ZxJ
Fvth8jUInOkseIN4YOg9CdKADKWyHhb2O8nZKhCuKm4pCKjvhxBBWjorvH9Ef2ebjlCvFcqaVaxu
O07BiRF8mNx5PNNMBDFYkHzn3NOk3xaGXktbD1hKvX/co7Bj1cE6Q9L9h5lT074Z/nmM7Zqou9H3
+B556l0br8B/ae1R7SzMUUCfBg8JCAW4vKm5IbpqOB4Tg3msDFgWIg7vcIDo0l9MRrugtyqudysY
OJZ3oR6qnhegd2nx0+fKcKsxxvZ5GMLFp5HKTBNZokZMK0LxI3ldW2TwygHRPQR7NLeP1M8vzczz
SuPaP2W9PAsSYKpNocDjMZ+UWBVJ//3EHhTPAEYYw1d1lr1ll3lj1Y5lfCsnHTDvCF4E2amgDEFT
QTglDTo3yXvuhJR8gr1Kw9sWPvjpMXQH4dg7f25vVCqBaku085trhLZG+jfZpxFFnvq2zodBo1T0
f5MryxXHKYpltCrRdsgvZy06ZFar+S3s9XHHVbsTRCEtsrwpLls69aVSlZzEkJqPspI92vUDCMsu
Qds9K7cm2txwGW4p5b+yxcfExpdBeNQhdYoCTtL5zf8sAUMCRANdlbv+tLf9JoBf1Hj5m5BNJJCM
RwQiHkESurv/PcoDbdrdGNfabcS7IpsYbX0oaqHgwvzl+6KJWXf0ghWbkBuISHaGwjGCAPJvFi8d
K8CWtihOi+CHate0gjbvHTOC4GtMnpZI+rCtQeG8wjUpfuo7HiI4JgO302YytrSWs/wDKT6EiYS2
tbUex/xOi30Aqa1r32bIcVnFKTxgYz/wKimnZSiIwJCnGEcbqyMUehyxU49W2ClpvIerMhZYTk04
ROdPRJwCNSMt+6ks+7SLo+YEQKzuHTn3js1516efa3CWI1mN/vTrY6AeDmuVABjH7hUwYTmMQjhM
Ll1DbhM+7BfcW6ddAGBhjGb3WH/mnvMwQ9Gd15A9MqZ7tLlcXPBumyCVodvGbYiqC+N6f6gvcxyK
vXXs6IPivzCXpnPLbVX5MWj59jk7dR2vQBxDWmiP+b4Bqdl2ZxH8KrB65ZXKfAXjAm6Oq/6LrwCe
0Dku37FjHht70sRDEBG1K9lBil3oIzacanHC+Wp26dsp/NTgYQ/wL2QexIPFIEUdrhGzCFLcTiMy
zG7TXixpETVT7GT75n4riJdM69HuRwj0FklBod9vDJvmZ2AiIFtDuhlxtFE9knJ/AB8A+Iqgpoq8
d/yNT5O/Z/ZPSJYpZfKimUkt7GEQ3Df5wAlU4i48fvG2YPCmd6Zc27dfqPoPH/NxSEC4o50kNDKs
8idC33mhl6wPPOkwu+XYCObegQF4C/F6moWjoSHVxB0UTiuKcl4bkxgInh0xq98ZWDjwz0IaZzX0
3Cc1XCsZRx/9y+lM6ziwwFIJ36U4wZvJkFgzQOx+Hj+m9XVwED/8XPgJqT2eylTBVS6eZ+XSfP5r
RGtCRLobUWWDOe3tgreLN2wx4vgV5AQ7EFW7KwoP2qPffx0bdmetR1XPYQo4o1yv7yNGKLxsGEi/
uZNzt0iki1jZPk8P2xJI6TTMvl+H7EGkEDFOZpbZxyQjx9Ki7dSUMHijQZJar0vQ+OvBUYm/wkKU
6K6/gLdz05M4p6AZybWB8+bnEXIwaJtiUiiRUWyarqlVLP1FyRMIRPdQ0ezKjls7uEiAGSotkWLQ
++v7RgfTbcRpWQ0AO7q3H5FpnYup427rqY/i2NYtrXhBzY+EKBmYJPswKnyJEWkpN9JwuM2fUs6u
Wn/xaGkoaoBRzohip/BJOJkpG7vCpbWV/cc1vdr8bV7WNgIlItDlcpoKwsSz4KA1ixyjTo5YSGfx
tkly97XVoTIO2248oCtX6LWPz96KsYvd+01NUIkzT83TlYXXZfZA46Rgb7/BepUv4+GQlvsw5Qam
29O2ZQJbEgIdhNOJ5GzfOat+skAhUt4PQCwgaxmnVLFRUlTHZYWHcvxNJKaDzoTUz+QGQK65sBrw
JxoH7+e+3PJ72JgGO8V2kQbC3RrXGCRyg2TNVcCY/k/oWBFM4rSZWhA7XjCfOEvnAnEBJDWQXMOn
hGGP4BPP0JIzwY4nEa9KnSkKNw1y/f8hBlbm375ubjsAIFD76+toTQywAvR9npV93Y5d5rtzLQF8
JmPWT7Ddkj9+jHtK9XFNbE1T+gqHs86DD6mEJfIevMvk0C/WBz8PBQKPmKYRYX05LGn7it6b7cUa
xdO9jLJi1oJT6ggGD8U4ZTvk23YLveZw9rUfN+PJZ/Izd792lv2Q1oKFmKtzGGiNDCBGOvawirE3
NeiZ1S81wo0mgRRzxw==
`protect end_protected

