

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
p7OtZBpltt/h9CD5IsJBmAQ+bQJxazkQVbRBjNJ7LWO+cgudo/XA7alKhPL+qAE8nYmt8n/nhFV7
1FHJnU9EmQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o0V8lbvMs2u7Pr48iEK+soyjigqgrrzx5HsGK4k7Ph8gI81XWNRtIljFPpaeGwucYu/H+gPVGgh4
LxNZUBJhgeC8kZr5P0UJ497gR4WHGLQSo0hvtVYHYDlrxnVk2S/+il/2gMAwvI5YF/lKiRUCJMb0
2mL6cpx+2git922rE9I=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hIqrLT0Q92Qul/GeORaSvJHHAIqLk6EmPwtSD3Sw8K7TFMN/pzvjFhA6g78oxGwtYju17YRUOAPP
BxWjMZac0YPGSx1A1AySaj/jWf8/sND51mJS4hxixMPKgd+iJln4gROFDpToYNAZ0eBhqGsKoRPf
Exo4YtwLGOksTW6jkb5XyScrMy9eg1uc2W3HXgQfQg9hr9gpWWe4xqhKUCFXFb9eiIDe3eaUQ22t
Qgz9S0YooH+uhgkKhXgOsKoG8s8RO9q+oyyLd0ANkoAdDySOy1H2+qKDhuJHoo8oHgkWp+t8x1nO
sbVK5ZibMfLbKeRbGwFkFsj+EKfWfOy4ck2AmA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O+omGGx7WVLIBeJijOGvFCJZ1IO2vxCm1x3fAW3H6+gw883MkRTmRZO0ddVzk3pvzQaBPeJUDRsY
1XbF7OM1C/khYSkVv9TjyhihrgNNT2rgkTkWtfQNoOMnsmtYkK2fHBBMyNXzHPZRBh+2VgTZHxjv
olfJ+wvlLAdf8BqZKWo1gutmRCut9sBqwVpKtMbEKFGRBnt2pETIJcWkewW45hEmUxoPlXpgWrRg
sESpeoKuutTTWJor2paEV2RoktNIWs/+x82raY47L1AIZ3uy3vEVemolA7/fyBhQXHdXuWEXntN5
bzesBXIrWmoZpCMSf+IISz8dywoKgC/dpdCKGQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pc9IPtPXrLLm2VmqSrmdhsB2/sqloTepqxhS9rXzXINDRuCWOADiBYd/5aw6fJ/PtHP6hvfQmgPM
pe5Rbb9vXhfZlTdZe6IYAV6ajOneMnpE0SRKlyLpgkbpQbwWF8Ta9x699vjybNfWF62AYBS3D7DQ
b0t7dD7uNK3C2oBkpBFbB3y/rTrUlQxN4AZtlp8BUDmTdKIOwvLfH64R9omltAgRoa9eT5fKR+NB
hJulrR0XnMdnz4MTDv9F/TNStcRrNIf5MM0b3o9Lm2heOPvkpoBOr22fj5c2jTQHuYFT3gyiU8GP
rFykj34Hi9/EcnhfJs9E3mtp1Tszf4e89AyXHw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Rp2qWT1ngiwszVInFfAgNDsqirvFBRH0fhGMVLdTcJjuZF6cagj0r5deSp/lHSGQXbQ6hn2NE/pT
sVS4xwCY2B03TkdpZqI4G+dZXB8686b5iwRUQ7S4WwcHb3WXRb4Df1OHJ6dgH8h0dIOxvwXXNlqh
PKzd3cQ77q4ZzFc8bvI=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JmHrUUSZT8PLNYfmwBtqUH6qJ1p97BdaA2q40RVMw79ZG2/5JMAd6P3xNNzdIISzZU+jzu0NYPxL
Z/zfPbolJrCwAck6UGljZ/OOpPHLUDGkBAu8BIP536kFNfmsl2/w8PHTByudSnwDI/YKiNqfsxGP
M6Sq3+TkXml3dJEoLhHWDNi1mL1f4wADZ5vEh09j4ryxXNWZ0T1vCwLDq6JQfC0fF5S+fWguWeoy
y4GDwuB3WNo6v4nkxnIBm5jk34GhklMVorbQQ90znGRfAejdTRlBiH1jH/CASbqnXiNzj4+1wJ6K
83Kv1+Hi6TU2vQtu3O5wYTXjTMpJrASuG6iNvA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
FYLl00vjC767GBkxsWuhl/zAntvtir2FQU6hmYSR0iWYPnMs1Pf6ckCP/mbqUfxyxZsF6cXX6sSz
moaiM/TRUGNpjPy2C5nxxWE7pMoi8xKU5GSgsyOCdFurQ632FGHu80Y0I/B1Xkhxo1kc5FMwVa+a
uaSc6ISNUOxA8oGoIcOg71HYO/0SwgqlW+mkgtKOln7rJUR39fjJfBdfQ3ZoY3bXepLUlCbRuJLJ
1l5MBg8B1fyTW+GsxDJq0fDsinB10YjwlPjdmDcO4Z3HrX87KfB3oQwUIodu07bSuHD0XJRPfc3u
XmYvHMMfb//0I8sIHrV/kT7z6AAmzNV1FCz039bwLVmzqt42RACfqXCfNo65rJPW5Vh7rcLLE1tK
y/PoKBUPJoVhV1xwo+9qMoFHeBl6I7z/zOKBStoIm0rpUZ4lpbwvIGhjgfKM0fnvyeXE5ygHfXo3
xMmNIIPyt3sY1jm1ulTy/phtWm29D+yOXWpIqKcPEkfpxOvVZYRi5o5sLmVc8cCF2SDI2RfxNC+9
igMHYf64nlfCgVw1Sg9xucZiIx9d1EtS45f7dUVfhv8aufoWSotzYOczxlnIoMuzR49R22s1dBhp
+lRuCdbPgmZsciwA/l7U+fKLqK+7hdXDdLkAUVnGChz8FW9r048gQPTtAvLrNhH0ddVLwgGfMSO1
RS9XddCaIcZeQAaOeSdbi5jii3/jq1DitUnraH7Q0RqJzOp6xvmQiQTDCHCihrqIC0s3pI87SLsD
Qu8ze78OJNM+Fgf9grq0qgSSncjuOubvYD9HzvFrZnIF4eVGA7i6HXltcG3GdUt+n6md/OoPi3Bo
F7CEoTHpUmOLdxADvfLH7KUeCDuPVbMzYoUw+2s9zck4zeC9D67JPzUcQsEVH+Iy5+J2WtUE0uoK
oCCzMtJn9tOv56VpMEcLi5RXnWRFFVJhSogyl9XWJT4B3ZRpgj8mRAp6bo7votU6iuZkIJWJGLFW
NYPad1P2EC7MvDKRZYdO0M7RuVjKacIKKVCWCaTj/9FdHfJwTVHNxmeUyQOEBSAhhRfMVuqMhay/
q+sCR1GpVxzVLtQ5e/ZGhsvB6A/DJnFAJmtXv7IfEEM9PJh+RtKU9msSgX5cWEE0KJotwd//Q1HD
6eeOyoMVIevfuYea8GqYb7NKMHfStrPM1CHKhAujR5ed34lb+yjUgEtpNUvKibk4UdBXMT9E6IOY
Yl3euI3Pa9eBcBQw6r9KAoRrWB6VAfU/Qkw7ax3BFBi6cUJOuEIwBiPYt4jW52xcmqHJEsjPMIcm
FrdrahJxxvWl7PHH78ggd8l4qDNhmOBr2wAddW9mhCuSuMsL8zUASa06fF4jIXiMM3BCTRza7+lY
vPnkwEtF+UwDQTRIaZYnyL8JWW+r5lucIhWf86jCgbRfWJsWQkkMUcu6hneo292PQ1DFkU+KsZ0Z
GdlE0848xQ9eBbIkUiNVxV3H3tx0f98EiNf9d6nmOwrVo5kf1pex0iqrTMsLG7t7BTp34JIlSbV/
+qTAjCOok6xzXKS5B9JJfyIOlisesDI6JUJszk/0R1zyxJ19lEQWCgr5B2WF4cSo0294fSgx0YyB
PYh2BWQTWqRgE+pRfhFNUXL+ddHteM70M4WIRvRvYrgOGxVOMqij6nbIhujeRWH0DKlyN1LBDjAz
045DEU5B/CVI8exhbZkXLIT6XcxW+JyJuj1Zt0gGdnSBdWoqDCO+Y870wBwbNRWwjVU3xbkQyfbT
mf35qaWOm6uY09FBUTRG7gxtrzrFFucRl2F2lVuWCm6dAtoUEC71BwDx81qZ+o4Zovugu+xTO1He
9Y1R6rFhMVn2LOJqY00lgKOaKA7aWqNOaNWKPNxVvAsEhsCzXAVNzTpgaQZYujobxh6986LyCtTP
5xkjXjUdZZXcuuiYLytMZMw8e4Mm8opTHN/22zSGWgIwuMgDZIg1LBhhOyR9hg0RoD7rr2SWIhc8
uZ3SvWypU0qKW29LGTNECobF1xwdVeAdecfTDMw9sosBBrukHDo5ZCJ/Q95O2doLDnVOp9MYgRq1
mruXgDIajD+1BYXvB3HvB6X52d0/Vs2umCoJR0pk3ZNhNUFeuPekX+QE8+Tt0ta6LWSABv8y6yPd
eGx8WWOy5lt7Ummx9V5OG/3vNwRdm863fW0whuBRILMEp27iteLR4ux6IkVVpoFAFFvGYxPW+Ebj
plBegLsYfkGnoVY4/DAaMuU8MmgrAnXwV2BdxzHqTQYJN0NtVpUKQc27YObg1lC1ue4orQVEV7xc
KJqUkr38j5YvKe6mbAtgcguqYxRodV+tf44v8lZVtPf/IIkki3aCQJuP2l6NJiWHL94G8v3nQKxg
Me7aNqWccLHA/9rUmq8s88bcERrMpD+ycLym9YkuLVrvhMCcWiLNwwHFmoVuDZNjwkQKCeBGZ4C1
5zEIy2N5RrKju50wpKsAQFcayksrtbftNufA05qx00cJQPcdsx3+1XOc1KrEzeQTo/qyZop24uyp
2V5G87uALNVxxTlbWokIBscIEqLUuH5kpG/iGTMJ7ttoYkd06V7SHrxfvVTEkav3MR3Sq9o5LmID
W/J5BWJd/KXQ3rD7QWRb1+z0iRGy5x2q3ne28oT0+dGxQ+vLjid03Em19Uylwk3jXkK31KqatVBc
xcHmfNJLrIS34tZXSThlcWhD8ZRrYeXySfIuDSdXWpSsnL1XeRTAEaLj9l5m7fUY+YbnVMV5IKfY
NL+TNVUouQhV71a/jACB1xx20qfnaIBN2ZEZSTXrbgiN5g6SjGoBlsxgTw3GTpTi9dB41mLbxMmu
CFtui+vdsPrDRV8iay1hBcZK7vLQRHDsnAELLc+BXgPMGvRgDGhqjQiFNlvwMI29nd2Cj29cpDXy
zpzbOl5YR9KXKYWh+22+ffx7OsmeQS8l1BOJmAxBfbTKSAc10nWTUOuCy1BsI8L1AEnm+lpYxLUy
HcGg6Md218E2TV1F+MOPWNlL6h305tTnqX7S9c4r0TyKUaMBGbEopT5g6lTepU9FU0uJjgRCKE4D
sXmhvh6NWEYMUba4vxmOZN3zccyfQUKH2j60NIF6KM/hcG0dSxABpPIhowpj48hVizro6SH/g3Ke
1n4VCXlrY4npbVMgmxbt9J5oVkyyL45A1XjY0Hk1xNEWz7ObHGDkrBs1t9XEyQt2kTi/ZQNrObT7
/xmk4IFGjC7qIxBkLpkWaDN38cU5lMlCusPD6kE1mSUDaDjpx7U3j2skNKyUIFYifJODoHXEyKRs
wAnOfGRskU+M2cniZ6VXWKwFWNrWBqpGU8IGXvKUKKLpACTCuie5MJbmdEWvCEQ2yUCYcAb7lFuY
PDaXTDjZ86IyzOZZR/qxmLRC9jp4+dTJ8yo3L1TidRC4V4SC6v4uMkwLuDJFSaubiopfsIwJWt6K
d8TMPdFwIiXEaj4mro9inJSrWCiSe5nrj5QzdjgGJv3CC+7DtzPcrSmvHQM5ukh1bwykvJXlTc9f
JJo6lWS3O+syPEvWtifWAU++HKK3s5L8bRWbp+2yNCHnxzVn+cBEXeIL3B+6Xk1NI0WqZl3432M9
qfLQYvE0dNz+vJVLVBCKo2cS+crb8qhzPeRv6kldzVW0OtqPLpsnXHVUUva27IYCOeIsxeflA1kz
b38It4E7z2IWgrq0sruqz3dh5icYerx4xigQvL9y252P2u0U4aoJvO479dYFOa2/rUiXQ4bYNJTK
cL2KqzZ7k1b2rGwk+oIole77GhVYmBwkg+3vf8ceMidWO4u0JkGSFKDLJZUuznVzcOEOwd7yrmzJ
K614rlJ8e3Ngl0iR61ftSaCPHtdSo0U4PuPbIN3DJhb2OxO7ROln61zqdoY3wHTzNnXak73RiqEP
joO5exs+FwsHp0X7qDbe7b6lyHBWfNosrdpwfkBZj9IpAJl4vmDd6rKYcTerEOAowcfwQwGhyHv+
9PejyNmtzmHPGKg+WNRvVGiHVdX9XSvslZ6z38Jv8IxMAkIvSz3KNGo6BWIPjIB3RDQRrfe+xtGE
7Mkzk17jZXxP19gvHdjCdOBTKgb3zy+EDUXeTOXz2MAYoslEVDXjeDRs4IIK4Qvfnrr/WR3KnbK+
A/PhJbwUGvDnfCgntvLPOaJMsqZe6XWmzm2dOP2TPPJfE8NrZxzqPEGPyFhih+WNAGnwqOEumOk6
ehy249VcFwH44xEw9yVXYiw4sreS6eQEeVKC0EabY2DTVqIV1y/aSKWWjgZgmXtRryplcDQV91k0
WrW/aBBoqAOtbk/x/OYXDRiWm63xpS2bYVdVN+W9ojV2yGvI4wBPfJYRfImDxwKlZCflJzoB2PRt
uqpGHg2zIfegJDZ1zd6gREYMKpZo90wWnRjDAup/BNVuKC9nQezGoLn/dmWr97NNgIQzYhHepeyJ
2pAY/XAFJy9kgjMLWnqmeeM8YelTXZrKTi6UKZTIWPrf7DAXBjaGSPxFuLat6VvHeBPAFekUwC1l
25Xaex68o7h2YqbSbH539sLoMCSj/6pwZgKIVJZZk84ZraC2AOatp/+eb5FM5vAJTq8cgjgwr+ND
7usuda5SJvjdc5w5zpGPB5wbw0MZr9ohUhAS2bKVwN7t0WxGibICtVbme+ONYM7DNKlLKReD2Bdp
KbyVfHB0XADPirJm+74Sr1msZ+taFzvHUHvyXJXGgjxUgVe9Nw6ul2H9/u07VO+WIHIXqVyOm2LT
9SdTWSKih6bNb/+R/26oPP1Brx2UvVLe01eDQGTO8+i+qi2IoK8Wx7TGKzGFTjzGhRer38QPeLAe
0vQ72W07dLYxq8fe7Cct0miTZQvIrDjrec7BCouSCBTnxXT3VVSrqwBShdFpKJMIybT/bZ3Xikoh
2tC2YN8DjeXNX+9eFAHelAHl0CkkEZH/oMOFOWMeuz4I05cmFVzoT6EA7ShGMf6C4hGSUkby7Vxt
+Th3tZw0Tl3bB3bLN/mdYYUdeAqKG0yjdz5443I/h6ln5BGHeYLFD1NwGjji5wL9nVg0SftHB/O3
M3UUq6XNUszaciRG1qslSvTZqGVWn1dpXrhTO9wvy6x34Hb80v/sbJYBEBr9FzIFMWFcDYVUhm4A
+BM8NDBvjkZqIgZEG0pi7N203S0k/5jckeGHCbl330+IkygU8k3GJwxsk4kPoTsmsi//JYMGy336
5TeDOUfmD7llWOKkt1iko1V3MDiQEeQRKK92vSXkgqHoLFmA0QF0IWcs9Jkpwy4yp8nk9z/eun/h
T9wJw1pUCC0zpwYpezGY/jIDRxBCntehleKC8QmKuQ8yeGAodkoyspJz7JjIY19GdMr/POn9Vss7
ZRIwyR4D7OC+iGX/M+4oruRVpG4M15JF1uoxb5baDWsu0G0l1hplnC+X3eONxzdW57bRSb21QT4U
VH/YeL2VuOc1/xjZjxZdD7fUg64Rs383L/2QfqTL5x3M62kGd2jEOrKUDe95FNTdtnCaXxZe4+pd
lFfYFoM6C8VYVPfapiOrxm33ZKiFMipvtodim6RJF3RaMSGiDXiKaSxG1W2laZqzney+EtIGu/dF
cPwkMfFZ+4sKkEYa2aRdo9axvF8O5iCrDQ2iiF8G0nSSqtByA+hzDr6gL8Tsfmn4Sb4+57m78eeh
6Hyw1qMkwjSwfG/ZJ+4oSet2oL9wX0wknlwzbfwKeSufX0RN+nYwpZYusKFOF1rKCFqRaUCrkRrR
VwFhbwKfxVGKYpzZPgVr6KjnerdLrF0QlNNpA/m/us8Vy1EdJUO51hzdw0FqhpPCWxWMofX9mJKI
odVDqbGNLuNllNtIzF4J1MLCIQ5VAc1vO0Wimm4TkTS2iSnvmEXCSHNagYOdTv8ZVKXx6IuVAlTh
cxrskaxfZp2M1wtp2NAc2PasOSoYK1wrrL8ZkVjmxYswXiNOUOQRadIojnP3GYBRs1OT52od2LSF
bHEd5MvsEU4w0cfgWWz9aPeLrg7dQoBcPp0GZVyUI5hZDRtm+KAEbbNlM3qJufeW5WQEjq3x4xYH
k5oNjftDdwhQIY/dfNRoclqEiSgM6YtF7OQaqflhmBtD9gYsXmzOr/haN5/KXZJJgaQV6w3Muhrp
MrW6CZsqcu6A90h8qU4J4Jna/MuWyDV0B+cI/ye46Dry88tTQaYMgMxIpMQvf/0xatF8dfXFQutE
8HapTduhlinQAGVKKNqP89t0xpmxxgn25NVmcjuO8GzATA7K7RAeEBuI6UeJVf1hVM3L55jlYzgX
IMeya1Kj3lFp67YBP4/mvPaN2Sy/5bbVuH8C8UD246J37ZjsvjAd213z6g3keM/SuUbaBZ2nbQOj
g++gInrR6bOFDR6EjbiGdurEIjkG7emXJeA1TWDsosTi3yR+YbiZtZKI7w5PXwZmba2he9XlYoo7
fJsFRUozs5G4Buj3slC6QvFl7rq1YuM+xepfnEf6fI/e60HnLfOEhaHQEW03ohovboClXOrzfqaD
HKUjEmtWqPN4aP1TGB0ETMXXAf5tbG5esVcT/fD9ET0XNH2tpPR4S1k6ApDKE4q8obWc6IZ0nwKJ
tdqq8cbcq3/OY6UNzGYHkLI/45GZs9AaqazRMcQxqwBS29afvdNuxVUOuTa4F4zKQBhzB153AwoV
8TfRmLMLa2POz8SbwJLXQdLNdXWB0szA1YcYxLcsFVG2njLGyNE5nijt19evtklFb5noywAdZVCN
KpU1p3DDcEqdGhZ5TbbH20dn+yxw/J3jphP88oQJSouKEk7vvmozZSAZM2WjWxpiYA2jePRL++QO
FKZHaoZM9ab5uRBIsn7saFZt+GOnXpu+UDVv0Dm38sESMnKPm4OxeR0Fd65XfzteTjKyXQ4/63VY
3Oc2Hvih/euk/PiB43BvMTsDuU73qabZnIlwAx9PC9jLTqP5vrZYDh3y9B/n3RawZffxl8ASuc+m
raRiA/rwzh/bKL7Cp6wgY9kw1ZVFx15HTHMpfiUU2vIEQZLs8tRj1x2G8zUFiUkRrUR70molbt2h
RWLLagHMQAGappr1REXxgcmtUMCA4H+VLCRy+8pW6X/jGOqASCai46r9lCNdu2ukwI/+jMiuEt+X
4FA+/OmvyxQzOKfI/54cUtbXduQj1HaNmKBtPmBznDHqd063FLUIjUYNdzpWgzp8MvL5XlO9ydmW
z+oxmqe3Ln/VieN3Fitijcb7yihIDR9qrRzrXYk8E4LqcxTj7tBLmrDY8jL01E/mX9+wSbwoF49X
J/fWSpAiBNCVDemQtlIK7glN8AVO6Wr1zIU01DlWM35fp+z0Kbv4X2AAUX8nyBl9t7rm+PfDKvkE
2lcBKMb6JtRY3omGRAo+UZxRiecIMl1YimGyBDTyM4g0Lp19syJQO4S0z+n2mb2jNWTvg69X5FvP
7n9Wn6Z/60Brl0xTVsSfvUE6MUWz8epAFHitUO+RdTKKOTLhLcDXmLehjgvcYTV9lhmThr5M9WZT
zopK8by9hQlBI8Ey3U+Vg+8YFjHs+IJ0hBvxCd/sUgkdcKgJybDmjK0lCu+QzuhEb6MZFJNjlrez
q4wS8OoNkOfjJtM2GOvjArA4eho9XXvc1uLliO4jQVv7xL471TDGzArbqgqBI5ZmOONVtGKvqCac
8LS89nL5P849MR9t/uDHUHpNbxNYq/PI6LbPXNSE1QRZ8PxSlaMGrJFd5qdpUt5O6RSpSw/DklNq
wfOENqUUYKLyR/2+zqWH6ejQUj+tkK1FggDjHJ1vjsu8Pfi4dpymQaqx0r5G8GgW0SC+4pq+VwL7
Yfr+nGZg526jWhNTpZduvfmGM7h1BCYQ0MYRykkUYX7Wa3u/XqR/K1KepyMhJzlubZI2WTg6dO0x
lD66iKKpuFJYe0bIi2YB2yRaypX69ZGTVSwPtSWnVZ4HhwTdf/AVmhzbvqqwfWfVUO0npfaskGq3
m09NdMbUeEob/11g1cizeU/MVdNdpB5lIrxXTMbgBiKjGFWnIl9HNFIipRhGNn8t0AUT9AlUa15R
ADX3g+oYQVogtwHwx4xuzR687ExpbYHgGYAgcrk9iKP+N0B3h8hgd+xsPJMN8TDF/DEnX5pUwTyg
NyIKML7GvmWD6JrZudtE+1iu7MQCL5icdLhinETs4DvGpz2ZPQlxER4M6N4sYYBXPSqAWpp9XDZn
tVPaNJKhJGg7bpoQqnPQS+Qw4/L0AeAHLvbrxl9tVgrqLidDApe4pq2MWSJo8sIXhQkD60pNJsej
WPFeg0Dg6K0rOy6D2pgtAZ7CSFCLd0iCaeFqdIx0NFSYxjFm0oyMerCbwUThQ+kffd+s/8M70UZ5
gn+hU724K4Tq9tRCvDXwAqkzAr7EgyrDCzx1Lvn2jPpI9VLK9q84Ksw8k2FVFXcFuEou1uQFkKsJ
iTGmM69RYmj4BHrTfis5u3tH6T1qcLBWjGXLqbY0jhFMlFH2d66T2bgvZfAvmn/hQ1aw3MULh5/V
O9MgdnDf9wmkwfdI6s+p5bl/yBKeCSuXC4JzJ5ZRXy/hcgumsh1YIDqo8HFIJbMQCdGj3NWEeu5a
AOycuVyoYRkXpvvUog0+HNcr3i7T1PMEqYILkasnorYucvaqw92S+MX57dkb6IoslZA/6PwokYlz
iW88i6OuWpg8KkrJG4VHXNb1ziQ/htYeHc4FNB0FjU7KMDVtkwrzz3vuQ/eCcymkk2LxXIUW0J03
VLAVs8SYED+S3p5XKGQsPyvW+kSV7uh4ItFkrBzzA+yOyWUMVnHbYfVacvwKgPxxdGxeKSyj7gZV
nqUAC+1fCacCIanNE6zgPCVaXQ6893QDbuNQH0vfHqTsP+uhhsse12FMpSw7xllTIYfI3vUgvfii
G+C1bc5EI325z9naQQ0Wzi+E0QeYpoN+/cTenHyZtAqv88L+8f0WJuycZXMkBHo3b883aSyvAIyn
iULtMgiprM8F2OjASgSvjDqh05gqPk/FKn+S9+hn4AHpMXgIO0FGT7dj3cFVyaUWej5GWQwBuTz3
+qi39riAGN3thf4E42uxuPM7sRh61INNKfhAGWElUYfxUfXV60bpQiRTJA7BJBbf0vFvIcmT2VhV
7pqAbyM5DejyekfdLgX+PdLdltaJ7KNpMIuzAiXg9Ne03tSwHsK1DQkj7nM9QHGWM5vMuYbV8AqR
sHaGA6nleKb2SniWRdbkgha5ZfWapG6DCZf6kiOOVo5iyJhynJzzuAT9l6n2FRT97obvYtTkQUpi
YRj+vKn//5cWc31kwOn81VRLZRRfs2+pIwLV/eKIO9hIxSwZz8a4iIZj8h2G+Zb+2TnvAYdGjusg
UfrCEGccuO/uCWcrGmP8OyKZ6D4PPf5IC4w3Lq3tCI5lVrO/OrpYumiJBrvIpLHZhlE/GP0DV706
LK8frfEAog6a3wrHw5UWc70mcTKVHIYA+IHt6yQs7CDBF6sgJrfYfSWe4kEZar1C6+v5fJftNUzB
3dJHzD/8xy6t3+28k7gY3HF96S3XIZyenk1za7p/vHPE1E4x/8kf4oIEGDtXG+B6AKd+cGeJauXO
Dlj32JF4guFSUdfhUhb5bSYCzcReAHNpW8ZIQF9mhhNLI41+1U1Hhpo/xk3B/kD/uzCp7/Qj7xH+
/DDj9TcaL9CVoFCIo3bLyUZGGF9r1c4nQvKuY9GN+Z0vPvLBN1BCRsKOfrWTGeFtZLzEvr9d7Eiu
fCg0dTcb/XwS9a6ajBD1QNlpcgth4McQF3vev0brgrYTTP7JQ5E5nmDX3yauUQvN37IoQ6y/d706
ts36RIgexfWtGWxSopgYNKxdq70PNl1eFej+u+TiHES5N4RipYruD1KH6OvSmwB/ywWg2scaFotd
p3b8Km0LQPdCE6rfUVSZOQ+52LXAZbONISCgkmmPQqe8zZ2wVzyQqrQID2D5Zm3vuFjYU7Q+NEMd
8lbKpXNRqjO390qU/0etntYMvTKztbJvUm+n0tP3QzgaZiUqU4Pb4vO71g/DHkW0+oNxkFTlmzOw
iKNppeccEqAexbjz4uWe+cxYDKTRe6ZRvqSF7fnOKlRloA+c5TkpmtnE4U6DYzK4Gf1Nx0QEOQtN
2rlV3zxoWsx9tEPrCSe4Ut7J5LfHFzQtxeqmwfgd9MxEtpKwmtf6+Z4JaJEobgMqHeXDq0XV0QgN
MK9LHGvsfZdUKlKKb/h1Hqv/S/ercVWNIO+FiGYJQSsneZcc8yj3q/VtBT8DK6Mvmtgi6ciYwV8H
QdjrUUcf0tcIvAkQTQz0WeRDQjcJITf4x6/VRN3aGwFuks9JWD56u0vHyTB9YSgFDpaSRr+fHEsT
Is7jKIGqGN/zdefdkCOWqzv/Bk+O5BMjQ2DlXtklvGR2HINc/ZFQ7DIk9oKXGM7+rjYO1P/giWKd
8+32QFeDFz705rKCrvZpYdBdyrsEDWp98e3OKOE+jEYRGT5M9igS08s4F1JTVm5NDSmFFU2Uq7lQ
FGePDEP2L5mIDAyWEKnGd61qqQWJ4ymgx2+2c13S3dCmUSaH9G60Cn6gZnPl+JQ35PY9LJkQhKzh
NUxyfP7EdSrGx4VTomOYuI8uRaOqSv1hM1XMjWoilM5jTh8UNnWmUOtZU6QCewzb7R8KJagRHh+6
rh3QzyIBsKr5KAR1mQ56ZANrvGAlSEoyMlL7+nbZFPntWRD5XFUrOq7TqbOPhRq/4DYWG5MBD/XK
20hWp8/r0U+CYUizV85B9hTwTGtyR6nOuWACXBmFS/ZXV8u9Yuxf6471H0xTqCcfTuVnUHVkSwp1
YLt9elL60I/BM8qNAuve7WDdiUvTvQt2j0ZAqCfdXzQirRo6kiBrEyRgPuyYAwQ4fYz2lNTLMlNg
VuvQq+E6rO8N67EXjEUmp2oA0Co+Cqd0lTGyNih9YTQiY20W36tH8p74+mF8I4pmVOOdnq2qGZwF
b1RxG0cytnXqYOmbgEPQ52xb2N2Nwlte9AI0Iefss0reeyQsdxNOJdrpouYdVyJ/zaRSXwSqWk2Z
pU2pqcTB0C7SjkmYjXmF7isQ/OTsqfjq4e0O5x5CgRorOoKOpyOzysIt9wcIkntIOhkx0DaFbUEk
Nz4JJugMp+D25YSdGX5i5JnSmr9zwebmY/yVIG6tBZxzNmtC/YTzvf8wSIpsTcN7TtMfnPxwzBt3
7JnBPVzccjX6trZwVvhNHt6NotwpBvXVxv6ozFACQwVj7PWez6fmdgCvTArQ92NE0QRLWq8r8ti4
bcxj6MNRWU2AbyLwZ8FX0gvIZoLs8PYSnZ50z8B0oa0MmvE6Mt817nLR0fc++siziZsyl4KyuPrj
asKalFFvGV0XW0JZJvThZ0BLlXwdcPK86YIQTt442Or388sQAjK1UBncNznNMYmaU/AKCOnAvUwY
12Frt5am3fS6cUAJCC4P+BvBqW0VxKund1eLEPU4fDW8TheDTUMthcXjdbBjJCbAXL7m+SkFupkp
WWUeZjl3hodbWuTH3NqWdM9mGerYQT44fc1jakvgCzJmxct5WJWoC2Cj7CO1WPFT90EUIXSjgHmx
xcgXHEgXqWw9inabQ8DyuK/FX2GLvUFLaWCxNdlvDm96OoTcNuHDsdomk/NBkAilXU/4JAU1GK8o
Qg9MPxb/8VOfBYMVzzbiU6j52qiStavPT2mlw1/sWuO5/qEEo3FIsWjvguIrhq5KFxp4jOek7hXw
82UV6AH+qNN9LZfLMy9tgjkmH0jzZWavbJK8gApNGAoO2Ma34V1arYWF8ff+fsXMpfBAvBBWA/Dd
jzEckFmXIYCeVYuGWwtWChQFO2gOL3SvsoRisA7mPI+7RZyv0Om8achaLy4hoikBZIpEgLGC9Xla
hy53rgXqtC/Dz0TAmiOT9/Vi3M3F1mJYje0upIPj78AIgaUKt4trmegYu7SN1nuEVQ9yuID7Xavk
ZEeDBX0k9ZeSnfjYt3rKjHsQokfYFsx0IaQqxg+bxTg7phu9BRUoEwc8Xn6cX8PKcBMivSadsyMY
7j/wF9tOFnSdNCsXi1liWZITYjp8Y/3cRnfzmw9nn9pyOw/sqwBMfvw05E0skqcGBGHaImHDjXtS
ScBTLbq9BcKFY1ZTmM7EfN3C1i8aAZXVBqD1cC2/rDiTxFiULqrc+nwRUVQi115JRsw53S0O1GQv
y7DiJvQ6MPGqeyi0Z3ZPzEUCxcdTmELTOLLiF69nsw6mJu8XG+H2qyDAeB1pwKUTEHYNM5lZqeLE
AsBheMsqjfIKDk8O2r8cGB7LrHEBnecjDcxXa+lMU3+WOgIFObVgsqN6NYIzTzK6fu7lAeqOPvEp
odX0GrwkzFljXh3O/LIGjG4jofKfJSRxovhjnw6CnfbgEWh5Xz5n3QV7T7YO6FsQxvmBhxjvqgpl
hPGg2E1p+XuzHJN/ZBKxVQfdEZVaD8rNij2tU6XbU68zbQ4N+FgXgmHQ3X8rMVD6ZacfnYOKQZx3
bpug4ik+Oe0JGdqbCxnxLkc7lbaqjdNm1DdemT6QLSRZS3vRv0xQRsCna8fFxV8W1mv30GCLILXX
+S8pSUWUNSkV7nu8D9krukwAvl0Usx7gZUK1rp3qIUUvgXmJuXt/2Lo5bjbrtpnyzFVID/PeRKcT
FlxqBzlAiGV2ZvaW4Tp3fFq4X+vAc36FxfNdKwLcFnorxkPRw0lOsoD8XCGb4KjsXhA10WszKTot
vm6rROf3pOlxoBSzDD/cBBebc1E11+ugIhy0ZdM6e8+ItJjUwXGt82RcbI/Su54nThHGjC1qxIuM
GdSMdxZMnC21qBfQDW55QJ6Pel5Uy1z51IWsjf6Syen/PQVDaNWzG833O9UhbE4Wl/FegTZ4Aicx
q9DCgNyWWWBOCbgHcR++3d4wBo9v14prPiXKj3Agu0IaPqRtAaV0MFTz1f2Ccz7s6dWFGa8U6y4B
pPjLogvOqWLhixvhGvjQqHOpAWofJnGAH76AM1HEyDhs7Mg66C1KcMIUssjNU6B8nXcmwql/XNS0
c3i6AUL6oFnqPNfOfUkPCft9w+tU+jgKWFvtM9KmpNoRZQ3SOkVJvT4SMN7WePE0wzr2QYXdyHth
A7PA1t5sb5hzHICTB3f1QcSLfb57l1lRWhQyroManaoWntueiLrXe5vs+o3adAw6tI0TWBHbHXVu
77CGl8LJXbd+Oil1C1nr9aVKdvfB4wlDly1Axvsdmfc2787YIUPxQNqerXi/4477dvahZeHxhHG4
TrLR3u9EV3aoTgvMHOsxahaogV8TzKoOgFDPAPIfZsSb/yit1hTiy2fg5EihBeO1LKVWIJxk36m3
57BxN1xGl45LxbbticNsy3HKIk6CCP40ziZx3PVb/uzMsM0YkHbnfGwXCWXyv7wq6nlmAS4m1kR7
OACRER5ZAorW5Cz03J+abKt7Fur6I+V5ECxS94cvF7ZyrEY95eOAwT9/jNOnQkL3ZaBfl9LTb/qd
31Sd+PnVZSxfMxsxJXEjBQ3yCvzts1LNPgtaP2ltwoPffPJqSV3Y7htjBLFsRoO4rDGduwIF0vvZ
p1S/m2vdSuc0XApYCn2aIPmyzC8uRCb59ZnDsRS8BcBNRM1L0fYUSnQuMX1i64rUyg240T/vPy8C
SMoIvRTSJlpl9UJG0OXsb6c/CDmxLi5QJk2G8pIJi5H698OSK/d5v3AazxKISuISTrF0CU5dXwgX
UvCY6fwrcYPTaHiC4Sms/9+FYgqQXROzMp2CLfVlMaqKNHo99mQ10vEMoTtoZnVqfPSMtj/76h2c
5vtkNzmBBZBn63drA9KndeYvWWKDtDQybsY/xobRnIId3jxUxczh79Rm33P63cOC7pudOWzjyveM
J3sa5mDeMieZvTdCJXqWcuUWqU/sSn/NdOwaUQLSasYbIk0PctiWnkKUrdd0AsCbtnjRlRrhj3zF
I/Ij2d1iZQar+8wlEce1ZZAfM7AS5vTtenKh5jd7+gOebVbQxOdJgAeUiAY5mzwZrMLaf5ijVRnv
amt3NqpGVEsmJkXh2aoZ2Jj1aCuUiZ7mc2R0U0/oNqCqj8E8YxpqMEmEHCMzrGQjMa/hbDDOLrXl
GOnqMPGxoBIJzObiWgYdSnWki8eFG0nGZ1bDGUi+ssIon66L9nAL5vSdqdv5oHN5oGuUby5d7Ist
ISWr4EtKP25YdZax8Dekbj+r4KYiBvtVZ4m1IEd0wjFtTNPnj6PpFMX6LpnBPnsScHZserrcXklF
vl8725R4azePUOqb1sW2s1geylUK+Py6SGsmC1+fw7IvdjUnRJS+8lhXG6SNC6+58WUSRaEKqbK2
qZh1uiGpTyBdGj5uUzNCjPR3oRA6CD/094RPS/DaJPEfekHeYPvC1/TntCVRlwnrVgpuiXJgcpP3
AfHGIoIUXCpsoTIjpjqUKfoakMWp+zM5g0Ltkhdn/pzi+W6jE+DWSI3syPRIGk2sZ/cU3BxXVLvy
pJcvsrEi7yZ5z4TpRQmrnonJASVSicBOB4lLqnBrENMT2dh2qUKvfnHRKOM6xzMf/p/3cpVDvJD7
vwdfHpRxL+VOF0ckUJ2qIe7Yo/g1A1ZpwvUMubnvVPagDWpPveQX5cGlcgg0k9nseIQs1PuvGpqP
Y7Wf0rqG/Iikr/vrp1aXDUdjYMyQy9bRywP6pKiuy1VdpThJsziqRrxsjwP637Qh2TKD/TMyYXDu
mYHTJjgd8T3VVR01SvcLkpU7IdOf3Jks3s746UUIFDbVYP/IZc6SIo9QLhhkYHnCRWqeMicb16LY
ro8i8yHk8C3wdGbCo66JF4GRSzL2XOPeVxo1C47VEvW3HD9S85z4rTwDyXthBXSnAnGY16Yde+sa
EWQqLjY7Jj32MfwRlqcWK7Z5EFWfK7MOMYU1BlMlwwI9k9IfCG/0613c/XXUKCJ+YN/OYbjwPgzz
q60vJ/GEdP0ui79bdYRnHGk6IBh3aDzuw5FuQmgOOlj5Rp8E847go7OqIjrnvWRS/IdJSCMEGcwO
969bvOobzvZgL6mDQRZ4Of61MTUN5AVv2Xe2T//SWbAXAYLkmAB1Y7K96hX50HjLPWhVDXlxogg3
nddA+TllgiVl1Xgza02YAFppbaCCixmQIDYgKbTVaFVkikKYPgro7fByz2dp0mEwrzO4HyMt2CrB
pjkBAGjSIrWNUtHc625Z/ijgGRmCbhu17HB6UeyrxlM6ckuZ0m08ht5sCjWxvP/5BWQ1LiPFoUMZ
TlYAInsgCNeuorlD2aJMovYZvCRMGwAD559rP3Sdh7ZyFVftjzbTriRbqgW19MOxVEjxPGDFUmKF
bfDIr+zBeXjPuf0cAmvl1aR2thyQ0tBL/ELKpMiaOhb9VWVDjp94jI8xnArRTvhxhDeCC+E2UFYC
+CM6H19EJbZv5JqeTzwyQpjC+E+3iP6Ul9ySfrOOv2OqVy/KziHVXHht3wbkCksB/WMqD88ikhrA
MWP1MTu1w7sNWuHiWf4mYaN2iIIThcKGoH6BWiAKB8Q742z9QFma5JD5qAYob19rNZXgCbyYrwVG
orMRZoCUZ2sxjTcQ40SOIWcc6Bp+cLNs7W1iEv9teW37+siWjnfYkhksCPN7FpIH315WCAPkBEy1
cWaEJBpxnj7C0GjllenIx6O3xVbe8CMucRPa7DGc5TkIFblel3ffso+DC9dAffsjmym9pEaqB5Cl
1Md1/qZMyYEmPMRXfrrS+1EBmrJ+9dd3QdnC/9nKWkKtptfAGJ477WN/LT+1VpHmEpwJUoxCLJEl
RLo7AU4i9on7z6EofmTAmfsEh5XEIOB83GUvsyEK27wKEwW/BWQl4lqSgfm8XMzZjncJPjHbPr73
hSEInIdr8VrqY/NojCP98gAsgHOgbPhAEzS3TJieCh2iHglj2L30KM9vG7lFDf6D+mwJZp/j6HLG
bVdToUUl8/AhgEWIRmlIPlFsOTSWm9Ki+Ulz/jOg3O9FOxiMvDGBIVhBRiTk5EptGeavl+QAUrCo
hRGvjxVhoPrKVlF9N0Kc+zBDNvekyeIO2VNsShDI/jA8+M7Pt95Kwi3c+TMO2OVjKH0sb9Ozwepd
NYsSVLhhybIo0HxKG6rrrq3taWDQ4d+5sEAzp5NRddvLFJ/2Sm3wUBrxEXkAtKTryo09ZphMME0t
meHHwO9+pNdTi1ZJkS4NDnTA5i8o4BlhFW2t9y/8NqfoswCah4fT//8ihT/fAzlDQ+BC+axVSbnG
WvMRuKkrLXqEB7ubbiNaAvEGXPvLesUEiDb08borY1R3flW2Qwy/qeIzEJth099ruJ36s8hJFTia
nGLbgxuCUHZwgFcF6ol3BixFRK3Ea/B+9VDxFloODA7/FM4wsrga4i9B4vN4T94hw88rhs0wNL6Q
KgdQyieeTjsqEgO0uAeIJxQg40ptEpeFRBgPhqvmfiMe/KOKHWtCv5fQkq6kFSVBak2PuPqE0cj3
Nmzv6WWiPtwMRElV38I2SEgGA2CHC9PbzILLNOLhKEZzbgrGAhNvL+XZanbKxLObQwzgkXW/RzGK
uTCxRRm4J8k5VCNfQ8SIhDV1Ybqp1YXiaMNQLKSW9iNdREybD9lCHj37jkSjJPR7muWibqklhGHr
V4nUEjBNTj8anTP6fpStdMg6NXYS/5KF0xaziE17i0KwigBYzcANyLMWhJT7S0haqkIluYss6dsL
sqtqTWSmaekfWDeAfDuzg8cfWMBU/LtyiuX8ygP5K+LGyxu+EAc86BrkbydHx7yQOJ7ZIMoEEfKp
pK+cguqCVsdgd8jU5wy+igtfTI8iqyNcypu50N28NdpY4NHO8WOWKvetRdf6oZsmIqlgx+6r/GGZ
NCz79yj4jMNAVsSVVMEPn/u3tA2TIdzA47618bDbCzlo3uaxof/F4TYPEe0qTFA8f7aqEfgfBOqU
wrs0J4/gdYPf5+qT6bkBxRHV/iLFrhOQ8c+0QO7ND0+Kztckz8fs4HySsF7gWb83z+NA+wG0kHu1
S3HAhMQ1MJguRdlkmmx842iOz0UIDW6yQaY+CGFx0j7/hECnNxMLBXZeDQvLEATJiQ759zs2ujIr
/0alfffqDdBjHCImZ/LXf4DouD3Kd4o9gJ4UAzqKE9Mm/8CyJO893LkeL0/5VGgTy5BgYrWIcaL1
Q5BtNNe5i5eKxpXUwrX2gynfY3vzr/mzT3DpORnqYct8um0xge1n4C6HulmphZLXE9P0QycJ7SS6
g+bTXvRVnvXF8DjIrT3p2b+ly1QHB3IlrsXjT0zT+JC3+YTEF8AgyUXPH7w5puVO6I6+aDqX6xFV
OOPCFl1h62rCMghfLjpjtlWpzhou9wIQuUZHh/0MY6OtHT3JBTdghqNt6jA75t3MK2UGFg2ZnzHT
DL+hVh03nxiYi3LNe9yqjlJUSZzDWcGgsLmxKhuK6pHshCjsrBlAtI5UwxmI5oSdeZ33j2iqeTa4
yeSlHdJAKSQC92pcsM2k6J06RcNMCqVwxIrz7BK+I1GuXBqbcNILD+Duztuv4o0dodEFeVIyzGqj
L7gDlZ1drXWDy3ndnKrcgw/zkLUPM+ilyTResE9ebCcR+Bk/opG8QNBhdB5wsXMpPZDllV5LgBH+
DWL5mCefN3lJ1QEozjfcTSCaE2nmMf1Bpfv0ZM70DXRRlDwrZ2bi/rFY7pRiiOLIt9muf1L3Trp9
JaRT18Mg8nFDa6DhXHGGGtJ/8TCXLlldAkoXHHphtTpt9/gsu7qTdIyOotx9Lf1ZPZ76dZFhG9sZ
desYpQlxiEE4lxqopPH8T4D7//zvoreDGUh9ayUqgmB9YaMVcvqcl++Udh5fcku4fvr1fhypoYh7
wpFtMIBDKkomdYTmt2VFD4kYGNdeSUtEtZHmcJzHaEC7UJ1UO7EonJywgIEHzPoYIzWijBCA7jEl
y7NjmQ/18KUe09F7wLwAzCn38eu2YuF0NrQm3Ao/PgGdkdzLCbMJkFDCVfNFc/8fNGdLqzAlHO8X
6aTf7n1V4z+slz+iNls6VCusrdtbI9D9q1IIttLQMArYS+V+/CgR8DrE3NaFKx+7ytzqRsPIwK+S
Jz8BQOya7wnP5SXYaY/zNA9Hv4ZApI4ir5Kbk2MF13+4621Co1VwGBYi0eH0k0ti/GQ0C2A9RpIX
vPkW/UVP7UgNu2tpCNv3jB8Eh51ZtVhQGGzt4DWzoLyFvE4q27UI3wk4A3MJQZwIth3RRvFIVWDQ
DsmNvwyadzR4fE/xAfdbBErMNOd0zFxkI18QEs6acHF6ROt3fD6wOB5q2jMU5ZiXU4RChD4UbKWb
EV2EcHSjj0ogRH3ukaPPQ/LIhVUQVOQI5JGZIpaZQzGZu/33M99erHy4g3bUq5eqNOjfB1lm6vBD
Cov0SwsypStc7tkV+yFJmVdTTOM46TKDUDbG+qK2d8arBKpDLVOCgN1ah/aiKWJvZdjoHICqPFZU
7z8NB9phKjdzpWNDo5d7N81kOAJvmJkXHgHy4X7d6FgOu/HNuxRc1G5G3zS2BaLFV0vA3GyHpFpv
eg8bHKgK3px39e27QEzEA4bT5ShUM6psC970FQu0wmIVv+pwkHt/eRBCLmGWXBTS4dir6CdeMQpq
jMOGGBf2RQai7EfCDk0RoQ/yKU14l6kXqPcHO7R82BkwftHMzWks9cc7ZShuziJ4O2bKDLtEN0+B
zNS8zFwRblNzC2y0WmkkJRwvuiEYFkaEQ7v/ragI9vJLguMA6y9VuHsjeyDBMDNyLiP3uVSof36O
fSm8xMKbiRGHt8oRYltl/ZHWWKU27ppkHsK0KXgxnDx1q1egZHJy0tEB/MV5NtYvzspaFiCY7qPl
5IgtW8UfBOd1DraTPTbXTgQbi1KBPM89cThzBShl+KDJLOD3E4aRlB6lfUjuf2/qddLeaNfJS13q
/IKfNsX/zicig6fGapJbZgbdfCwo3E4g6/wg41+CCQSKa0VacrCC3e0gCJGEC9Zd/jh2i95HxEkQ
Y5rjYlGZ8FAnzpPwlNd+uXi/CM7XxrKiffdDvn/M0CfX8OuCfwPnlg7mDEu6rPK+HHMOUyD5IfsZ
0z016q6v3BS0AfFdUX/iBcXinXfgyrgwHIcehiHIS3PM9rWapf6Vc0LCVGjb2bnWQux6GOD8zJka
L7UgReIlOCjrStFkkHpzpp3sCaS0IFGbXOSl/Ff7DGy+8BA/ABprMvPzb17ctbcf9+fBe0n7Rfu+
oJKFQFr2beVFTfvT8JNcikY+5gHHBR/giqFISQvaP4rGKyMXN290IE7LJNR9r0ZhMkb0Gyoz+mWm
6rF5Gg8BYGabWFru/YNKn3QeVwZNDFGS60HMu1gXau2X3qJKWp7Otnxxuv5zgKBBp89Q4KKRu/Pq
Akwwzr+gno/yPdG7uhlTdkLC6+iGKpnB31QrgLEdSaXqONXUPXeCTrOzL6DJWYaGhfH/sg+0dbMG
RpGzxpHtjLFD/YTMWYIuwqhn/A5QFFeu84TlPU2DVc+wJMA+Jze2hLk8rzeOceXSFJCm7Gu301fO
bZMLH296zWAe+cNxXjlo8cpf3yJtPN7kCDx65ZTYZNeW4l8ocO4fOAjgG/5UXoBzjuCiP+8/3Kx3
t9YgRHzLBs0KJeZo7qdFrM+YFXej6hDH1qOz1QhWOSTqBvdGD3YXTclpY+opWDEu6C1ciIBWF8sd
BqNRNzGn7akX8+pTClmzW1/yruRajOv98I0R3xw8hEJ/2AhWiMklv8N6scAkejWP6+OEt/lP+y6N
vye0Ecz9AbtkYAoJyVIHqkVPBfphEwBzUobVlCKXF4yB3uPJRba9YBS6etVbSn6taJo4eE0m/Y4G
jVJS0jgwUlp/mlEFoo5VlC+E53MmgMngb4RigaHbNg2+TOzm0UHPdkKB4e/uYVLa3Hf2iR26Fidg
opITvPCjsLsJs4NfEkKYA1jm4QKfxzB1yA+ppvXybY4VuUVnng5uJlTcyvZj/ODstfTXVpsbVGeS
SgzSU1R0rYDJ5PYCXfRmxaWQuV1S8tHqfxXVKhxKV5dp3fH8iOV9kDOPivhXSF7NR9lBsCwGDk+i
EjzCIkx6pa47/lKRTFsJZLOcxTUcebTO3hB2IS6+8h2Kj34U1sbsQBlUCzH9Wx7Xn4BUnJLW4s5T
3tbIyj8NNfspCNAeC8rtub47EUYNsBxMq9dEO0zTbMTW5HDhyD/oY+HVEBZ0SrVr1H+w14YCpJ6R
TdbbEVqC8JV/ljIGkHJL2MifQQu0jFYb0uiF3J/hdw7bTJtBa+4vefxLL6lzCaWR4ZPzUYjnm5n1
+9yyLBWXnMJDEyN4ovMWQwSdAJLs+qTfQ7BuN6B0EYJwMtYWT2voNqwgGd/uesEZX0C7Ll6h/piL
jwETEhsNyBwN4SqA5Lfm/daq0tXOAfgXn1RXXQZpNVq1aalNVK/Ci5YNmGnqYNN3IIMLHXR7m4Ew
q/g8EiaWVSdlOGi6AHcQQgnVqEdAh1rHDdz6asGyus2AJW835zTUOUBx6ymo3UhztIvahX1SYTHK
YgwkgYSmQg19bbA+JL3r0k/QK6T+CMFBR+Bq3tmcfRL4PjwVyQED/Ch2QlE1I5Asm7/YzWQiawG2
npHR3GPkxqL4Pp4PhWCjDNVtda6mZz4CoOWHEpY/4w472zMzY+i9YItXLt73Pl6SgSMGUzidf7WN
ycnGmTlCFK7KqNCZ5HI4uZ0ZH3TFIAsxs5iXO4vqjZSmptoicR0BwHCW1q2H/bGNj+xMl211CyAB
HChxhIbN51d5oD6IIXOHSEqBj9ebODqMJ2mVykKUZqbxPKg1Mdqld7hej9JbY5ss1exy9A56o/XT
KQQOlvJ2FCvuyKKB9DVxHmCcGBG25qfZ2cSZGkiozl9HLYUcvOIfd4sFXz/qgV+DlFsEMjeGwtFF
KbH256k87iSyNhJF76zcam9/Ack8LKwkeFXS6SYxEj16hGW8NZqC2kTO/MDdtSk0Xp3JLON3ry3v
b1qa4RXj6vbVg/aAuI8Sl+RyBiE06fh8w/fjJjb5Cpz24HrTZJftPzKAzqzR+v8SMnCuJqKp5lWE
MA/im1lbH70KwOrEW9szUZgaCdacW+MEA+x3RStZkXlUTzGIieQelKhUoDo24s44+nyXL8pw9KPD
dg2Mgg8hEk+lYcy71NnQgZOe4oYkKbLnOx/qU/aH4Iqu+SIH6NNNpIFFdsZ9CHeZT6xoqXQIgTh/
r35rgQiYW59kigLACPQP1jV+L2jvRaOvTxu2uxWPGUHvb2T0H5gKoTAuTbPOMWydkZeR7eTpxKDo
kJ6dAd+vTB/Ib/H6JbAQIhtiYGg5fRmSe6uUmYW5ql9d5Zn1GZ6VOwk/anshsZIocqFSZmc9qkQE
Q8gND6HJzNrJA3HeQeDoQSNwjWsycSP6o/8TvswGIzPwklsSZ8Pgy4BPgjGY9wfF55umll4hD8//
Omvr90l0q3sun7lsrj6bEzWc4ovS2Vcw+cF7estRJb00I82d9Ukj/LEgKSgIZkL6C5MvPECn1JQa
xY82XtnuZyFPjqwp05d0Duf/Gel6FCMFmxezEG+RtqDc0ul/psjFh9/qi2mHvqZvEti5zKmq8/AG
6Y1WISdIuhS6r37dxzHfa1SD+aqXaKtF7zgjmjYerFqkhSKopg3tt3RK1U2MNzHNIO4d2dWXKMpx
NbcetUqudCgwy7UfQcyuCcmZ+V83UrbFfqEY+syBehVb3hPV1jB/xnU2KqOUMsX5AIO6EEYE4qAu
lJ0ipwYfLXPhf0yH6UDj5nG4VIumNuNtIUyYi4gJWrX94mREG+0lbY3OY+7+QkORUlKkeDsQ+u8I
pT/JLaqkYzTeHQ5+on3vhtTfmI3ueuhXNfDSSxQgiYon06fw18QUuVc/9eZetsIA3EF/NyUb1OeA
x5UOqPEmnxdyPpqvvOaji+ZOk++cczx71GS8SLu25MsfUH9BnsafHmXWdzxtR1P1N5ooP/2+4o5M
vhqJSATjGnqzglUYeJWwVWraY1lVvxw+R66ZUM2Gx5xUHhPgg+N0A6mFU68jXc2WVU74qGUsR5Qs
5E7ZNB/N6EnqUT6HA1APP0ASfgeN4K9RYznd7Kdhb6AWySZO2aW+BjYcxwr13fOZTQuK6+iAWkTB
+GGaFw0zhAsOqkFEm00H6xAzH3JkoEjsinKqklgfyi9QW+HIEqE6IfxDmqDcZdLafeGkZsICbPwm
MQlJL/r8+4MKHQJpFnkrkVKuvG6PKEeBDutf4No7YqS6o3iq6O09j4yijQbEP96MGdLmpVzd5r/i
mcZDAlb/V9rBwySKbyw3HV1RzYo6095aJLwn6ka6NU7eG4LxOTQTAVIcG2DuUQ4eFJ9UDE5B/gsA
Sb9sG8UkfQtMqYou5xze2/lemPEW8WASIuyZb8ZRAvjHmtNN6+NQbdHBLcTq1AJq02xMDW5P9dlc
DpWyh9HVNQG+D0yakmhhPE986FuSOMzp2yGROzS/2GVvap9kgbv9LXrPHhSk0um3gL5iEC9PVst4
W9WFLoZR5tKcH0NfmFjkKp41TOisFAikqg5Pamsg9vllrgg3uP6d8jRVsVzF9howLLmBJ+E5qbyL
cwfaQ2eegoO8NsHsEc/KaFj3t622zEM00L7jFtqT3UC3pF655jkGRZbTOZxwOC8XsD48sQF2G6IE
qPZdzgH/TA2QzKyUm6sUCEk6+n+cNVwinqwO/MHTHv9+jZPSlGrjNeORM3Xsr+hdbPiKCAEO8WBF
XQk3qYBGviOT41Hu0APb1/ungw8ucaWbW+39cfM4Erfmi45ALYGCySq/lY3AKivO9dzJHng024cv
BuIFd3rF4BdcHb3gDb1/aSPCjM++pYwkL+AQPRjQzqAcYzfcYG/jRtS0DWKS8oSuCaZoAHvVY+V+
7t1qAsQTy5KIBanEcxgs/TCHcgOsvy5FFVwvmRBEyR3Ckw2FSiJ8PpeW5nlKYz+mtD2e8sTFpxCL
HREcucKSI+VO74Cl0EXZd3TQHU12y9IvR+D6YlvK/u2vWFvtl5k3pZfsFnMakmKLUK4CQw6v6/I+
W+rkVVf0Ngy84+WazO28KyRN9/ckqQmnd3+h2OamunxFTzHbHRGaUPt/BOTOmW9DJ6aIh+obIU/m
PysND9Ff9cLY9aICj2HT4sECHUj6Cn/EpwfhM33Z4YlYRYo/fvWsWBpx94L3V6NwJerwh39Rl5It
lAA4wO75rohlU2hTf3Mxqvh8DKj/4oFPYMwJ0K6DEHELl21/W0mWubzJec4Xg86XRyV7V0KqaHKf
1X+jX9vHlENFi5h5h0e7Z0L6flu2NP5x6zPUiShvCNyW8HZb+Rx4oeFajG/90GNFtycbw/Djf3Ft
ihtmHE+LsLccSjwXvbVn7wkYmZd0Mo8L3M8Oy+nqoscu5aDfgcsUT2dJFP5xEELcoWVjixFEob8H
hxk7YIYO7wejXEU3V98Qg7PQtx2Owyp+uF+egNUAyGgzZh48AMHzC4lVnfuMNhgQrT/B//omYPwJ
quVW1+GoYWqNZQ5BOSdbB0fd4RMYEUH0J1uOdB+f6khhjASsYF8LGyuziLD5fKJGJxtGtYLPqP4Z
qcg2hiGn75QutH09N8KLBkawGDI+hcq0AlnYPqcYvzyxBSdr17QZcGAiW3ksVPUsi24LVllOWtok
JDA5hTHYEMddomRI+HFoI8oXHpQEcH4ssadmm0sF6QkstgRBynY8fIcsgrycYfv8gb7WQCI+v4wA
6UJ01S4hu9LjD/iKVKNUCUyFzCbrkPg1scBw7+mky7YFIbCSFERyCNcqZvQonFPseKjhg8dMQTvg
W3sfox2rDTBMZ1obEd2/dtwJ8fyfRdwxBzXFyZbIls0KKDkX60hNrWAAayMH6JjZjDKBpoVVyvQh
4w6Jo3jmKTzJMMoy1I5O2Qs4endVY307W6aS5oAO9MY4/IxZrG5mgy7CnGIzxcoln0MAsDBFXTRV
GpYy31/MNc4InKEO2eVtXh6/RAd63SRxZJfAdU8NIbEihFy4NE2d81bmkr4kcvh73hSJuljI2MEu
OMUEOQhj8y1QNmBADdYtZn2unfwU6miVSCaXcQbV/AQ/8SPqSA6C6WPXXI8dXRQ8reOnB7NP1ksR
gb0kjI/LoHvBsyLccYSPAepRzlmsU+jLuw3a7QGdbokA8/kZzHJAnAGlPEPB/wR+EQecQNLstwHd
37H2BihAGSY60IvRqFBtRQIPOpuMbarqFyBPvvao3p/aIV1rb2l2Xdv1/yA42eg5sbMAXCJklspQ
TOk2XbEmH9TeLFpgHYvC+bGThRYUInPCXwoA/nyMlJ3K1yWvkW8U3dg6bKb4eLmvARCQ2YtzygoB
a0Vx/S2oE5JqbcO3zW1eWiUmBnxKbggk4SFFq6dVF0kiS00kA/eqD97XOXJfS3NVxY2BXwpZBuy8
tzPG1VeOqjSkiNn1+cri/U4UeZCDqiJ6/hQjfsJqwkimTsdtrAq+Cr6tUvDIpKDgttnsw/P+3pES
pClIxUf/uPehs6dBjlZBfC37NQ7eyHd9MSVGqEYqeWx4pjws9mGxEKKRlAg9WaofYgB2b0AP0mY6
FxYHmb/kyIGZyaY//d5VqzumjAtUNk+W4/5AenhOjQdpwoK/7pVtbK3YHT9ANj0zTUxDq2uEjmcN
stIAl02HuQjAlxbVo5o24zyD83H7ZEZUY8MrovI5eUJj8qgsn7YF9sfx3TtGWcXnNGsQOCmH60C0
vyj4lVKBaGdRGkB3BsMUyEZB1/dK49cW0Y8klJ4kW+V7KpA+Uz0/5F9ptn/GuhNcrX3ePWnXhXB8
MYVB1EjhJXGHH4C++twy/z/0ymaH+IKqcu/80ohAb3sUdqkbvWIzqtI7/qO9RtXFxmbOShZy895X
x1I4EaAld/mzyweNqakKuClrjrmoXiEt8DhO3Pyt8SDm3t1TDf5uihQsEve/Kx/iZN037kKcCVYd
q4HInpiokg/31+RvpsT0+dFC9Ja6Ton7cYMLZ/jZic46Tgp+IlDAmCbvD4Y+lQc16uSQgQVXWCKP
AcASz0I/7zGxfaLPtdmcnGn3z1zV/1lSNj7Q/ckoxwsZOB6+g3FInsnTf8BrcH9cMGo1CxRY8Rgs
zVrnpvdyqmpnZQ63xH5CWoKE3exDGbYmI38d3HRY6AaSSikJaSen+8VSOEzVMLGsGpVwmgoq3d5X
fyL4/7Q0IZPHkcARCDTAFFQKWoXebs4PQRuHieSYmIzhCpiH7qQCJefsKLqxtJUtZ7Gw7xRxOiUU
chTNJhEeg8nYIUfobZt3T1/ll+ufhqu6z1GUM2SL6H5pwgsjFBR1M/xSYDtDmIaCv+K9oaa2m5w4
k6+WL0bj/VG8vuUG8eugxiyinEfvtfFWtjMpOA+FFVpCoSelQ71ggx+dipkJH1s5lwp2cOtRyAfY
c/9r3DE0JP5r6Tly8pG81iQXXaoFBz2D4NIZJsaKlKcnCCptH4gYZe1Dp/XAgjLctZYfKWnuq5mv
37P3HO0+bWstktyRU/ZgZk9gFBJDIjdc1M/GnU3rZ+kF8bif/C6lZFZilGub6YJEVZnoyYF7BgKD
qnFOaFPZeozgbkD+dDPWUcIN/2kKg9NO2FylBkNi+gUItOZXFyOSVKGnICuMJxNz99avZJl7SyRe
ixyV0s3DIofMOpWQ6/D5emeTtLPr0W1QQJfPyIsuBtU6RC94y7VyYWdlDETOzhpGZEFU/X+5LCQy
mBXpfGRFqQMj5MNp61MPAUZrWaQnuJOXhmeNYRE6oBYqXs6EVBlN7E1+NXtttFTdLp8GVJgOf8FJ
uU5HQ/ZfoQUO/s4A+SJfs/ERIb4WZSZWDBCCNd3tjkwuaeQ2daIa9isjEf3dH7Uh2W47Bbo80Glu
zlTFu2qt1+My5Gh+jCPJaGolxE1KOnndn3YtspBrQ6UGBMibnRbkb5yjOrGqvtdXpKPgd3uN/bxZ
eTOiuq4Sd2JDV9o8fizl76OGktMFdVeg7dEaaz0hGNXAzmplYCuOZ0AVSGYx/YrCs5j40pTxywWx
ta6p6BnX5yuPmvgkhOoMDf1lXZoVPV3xpZg1ORWmHfbMJL22CUBmvhvEmzfE5OCCYscrw1UyqzU5
bNTvCkAxmiSi+D8YPPtnFbP5D3eFidtSbojnyi1f78Qq02dvL3aLBuqkSJZ8A5qcz/PB2ISaT3UW
Y9oy4uHKtS9qNk6IFvwaq/s5mgHFIpOPfhWVgW8N89x4x+3fP1g0xEd8eMnyu9wNoC5Y9YljQPla
UQtEgyT4SlAn7sOZlaSwQkHeo41f9Nwzvnar6Dtwl4nmBRSEOYklATP2nQogza22oruy97slSG8h
IVD1N0w58YX9dM8gNUeD05pOCzo49Azu1AZqAPTHzqaCzRXnLjuwaQPJN5kECEIt0hF3SX+1CV+s
oqObilB1xvdsFKNyByTcXEsM0oQ772HyzHVpNSa4UiU48lP0bxFuvTKXb9e6XZhVKkFjq1PtaLhE
gaEI6zp4BQzV4OgcCu1JAe8ZykVpb2Nlzbcwu9MavK4GAiTnguZ/LwYI71EetMrzxGlAWKNj9cPM
GpkyvCmutqaFDOb9NUt/Fn3vR7aqfgewl3Q2fljGiLTuooZoqu2wdfFwtQ/CVoroVjNX2ygxcGdP
SCxPLGnido954849YNou/vZSgc9SIloc1VDmE8iz0/JZJK1b6OjAcXu2cu/0hOprrwKC/mI504vC
rSgHqpl6tjpNbE5EsjBR4Yh4x9rbBNLHGM44jDrPlHfBmI887OsgiyVt76jkq9rGmmooKcFKyGdx
VrXZAi/qu3QkI/CEH8Rp+V9RZSu/BUIdD/QOO4pD+/MefRMywYzEBDa4mdN4eS/ybFhvtvU3x8wh
JWxfpKh2H8vvtSWUqGxdxX1Mv5FqH2T7e+vn5PVtFE+UxmOtML7uQo74CvvoIrPTdE7j23zHip2U
Lm6679hgedxbRQGS6L6t8+SUumhi5YSrTszTARnRvJ8OdWQ6mfon2ULwTDKGrrRCAVvzTdrJt/16
WYnIVho/Mw==
`protect end_protected

